magic
tech EFS8A
magscale 1 2
timestamp 1602042344
<< locali >>
rect 9631 20961 9758 20995
rect 6595 18785 6630 18819
rect 1719 17697 1754 17731
rect 6975 17289 7113 17323
rect 9631 14433 9758 14467
rect 10103 13685 10241 13719
rect 15703 13345 15738 13379
rect 19659 12257 19694 12291
rect 12587 11305 12633 11339
rect 8159 10081 8194 10115
rect 4663 7905 4790 7939
rect 17819 7905 17854 7939
rect 2455 6817 2490 6851
rect 2881 4641 3042 4675
rect 2881 4607 2915 4641
rect 4479 3553 4514 3587
rect 3111 2533 3249 2567
rect 4997 2295 5031 2397
rect 9413 2295 9447 2601
rect 12173 2295 12207 2601
<< viali >>
rect 19692 22049 19726 22083
rect 19763 21845 19797 21879
rect 17417 21641 17451 21675
rect 19717 21641 19751 21675
rect 20361 21641 20395 21675
rect 18889 21573 18923 21607
rect 15888 21437 15922 21471
rect 16313 21437 16347 21471
rect 16932 21437 16966 21471
rect 18705 21437 18739 21471
rect 19257 21437 19291 21471
rect 19876 21437 19910 21471
rect 14381 21369 14415 21403
rect 15025 21369 15059 21403
rect 14105 21301 14139 21335
rect 15991 21301 16025 21335
rect 17003 21301 17037 21335
rect 19947 21301 19981 21335
rect 8677 21097 8711 21131
rect 12357 21097 12391 21131
rect 16313 21029 16347 21063
rect 19349 21029 19383 21063
rect 1476 20961 1510 20995
rect 8493 20961 8527 20995
rect 9597 20961 9631 20995
rect 12173 20961 12207 20995
rect 13312 20961 13346 20995
rect 18312 20961 18346 20995
rect 9827 20893 9861 20927
rect 16589 20893 16623 20927
rect 19993 20893 20027 20927
rect 1547 20757 1581 20791
rect 13415 20757 13449 20791
rect 18383 20757 18417 20791
rect 1593 20553 1627 20587
rect 1961 20553 1995 20587
rect 8585 20553 8619 20587
rect 13277 20553 13311 20587
rect 13921 20553 13955 20587
rect 16681 20553 16715 20587
rect 18337 20553 18371 20587
rect 19349 20553 19383 20587
rect 14749 20485 14783 20519
rect 2237 20417 2271 20451
rect 14197 20417 14231 20451
rect 16405 20417 16439 20451
rect 18981 20417 19015 20451
rect 19625 20417 19659 20451
rect 19901 20417 19935 20451
rect 2881 20281 2915 20315
rect 9781 20281 9815 20315
rect 15761 20281 15795 20315
rect 12173 20213 12207 20247
rect 15485 20213 15519 20247
rect 14105 20009 14139 20043
rect 16037 19941 16071 19975
rect 16957 19941 16991 19975
rect 17601 19941 17635 19975
rect 19993 19941 20027 19975
rect 15393 19805 15427 19839
rect 19349 19805 19383 19839
rect 15071 19465 15105 19499
rect 15853 19465 15887 19499
rect 16957 19465 16991 19499
rect 17877 19465 17911 19499
rect 15485 19329 15519 19363
rect 18153 19329 18187 19363
rect 18429 19329 18463 19363
rect 19717 19329 19751 19363
rect 15000 19261 15034 19295
rect 20361 19193 20395 19227
rect 19349 19125 19383 19159
rect 1593 18921 1627 18955
rect 19763 18921 19797 18955
rect 20085 18853 20119 18887
rect 1409 18785 1443 18819
rect 6561 18785 6595 18819
rect 19692 18785 19726 18819
rect 6699 18581 6733 18615
rect 1593 18377 1627 18411
rect 7481 18377 7515 18411
rect 19717 18377 19751 18411
rect 6653 18241 6687 18275
rect 7297 18173 7331 18207
rect 7849 18173 7883 18207
rect 8401 18173 8435 18207
rect 8585 18037 8619 18071
rect 9045 18037 9079 18071
rect 1823 17833 1857 17867
rect 6285 17833 6319 17867
rect 1685 17697 1719 17731
rect 6101 17697 6135 17731
rect 7665 17629 7699 17663
rect 3065 17289 3099 17323
rect 6101 17289 6135 17323
rect 7113 17289 7147 17323
rect 7665 17289 7699 17323
rect 3341 17153 3375 17187
rect 7941 17153 7975 17187
rect 8401 17153 8435 17187
rect 6904 17085 6938 17119
rect 3985 17017 4019 17051
rect 1777 16949 1811 16983
rect 7389 16949 7423 16983
rect 9873 16745 9907 16779
rect 19809 16745 19843 16779
rect 9689 16609 9723 16643
rect 19625 16609 19659 16643
rect 8125 16541 8159 16575
rect 8401 16541 8435 16575
rect 19993 16065 20027 16099
rect 8033 15929 8067 15963
rect 8217 15929 8251 15963
rect 8861 15929 8895 15963
rect 19165 15929 19199 15963
rect 19717 15929 19751 15963
rect 7665 15861 7699 15895
rect 9689 15861 9723 15895
rect 19441 15861 19475 15895
rect 7895 15657 7929 15691
rect 19763 15589 19797 15623
rect 7792 15521 7826 15555
rect 19676 15521 19710 15555
rect 14565 15113 14599 15147
rect 15025 15113 15059 15147
rect 15945 15113 15979 15147
rect 19579 15113 19613 15147
rect 9137 14977 9171 15011
rect 14381 14909 14415 14943
rect 15552 14909 15586 14943
rect 19508 14909 19542 14943
rect 20269 14909 20303 14943
rect 8677 14841 8711 14875
rect 8861 14841 8895 14875
rect 19993 14841 20027 14875
rect 7757 14773 7791 14807
rect 15623 14773 15657 14807
rect 9827 14569 9861 14603
rect 13829 14569 13863 14603
rect 16129 14501 16163 14535
rect 9597 14433 9631 14467
rect 13645 14433 13679 14467
rect 16681 14297 16715 14331
rect 9781 14025 9815 14059
rect 10517 14025 10551 14059
rect 13645 14025 13679 14059
rect 15945 14025 15979 14059
rect 16681 13889 16715 13923
rect 19073 13889 19107 13923
rect 19625 13889 19659 13923
rect 10032 13821 10066 13855
rect 16221 13753 16255 13787
rect 19349 13753 19383 13787
rect 10241 13685 10275 13719
rect 15807 13481 15841 13515
rect 16221 13481 16255 13515
rect 15669 13345 15703 13379
rect 10057 13277 10091 13311
rect 10425 13277 10459 13311
rect 10793 12937 10827 12971
rect 10425 12869 10459 12903
rect 19717 12801 19751 12835
rect 9689 12665 9723 12699
rect 9873 12665 9907 12699
rect 19257 12665 19291 12699
rect 19441 12665 19475 12699
rect 15669 12597 15703 12631
rect 19763 12393 19797 12427
rect 9781 12325 9815 12359
rect 19625 12257 19659 12291
rect 8493 12189 8527 12223
rect 10057 12189 10091 12223
rect 8493 11849 8527 11883
rect 9781 11849 9815 11883
rect 10379 11849 10413 11883
rect 12633 11849 12667 11883
rect 8769 11713 8803 11747
rect 9413 11713 9447 11747
rect 16405 11713 16439 11747
rect 7732 11645 7766 11679
rect 10308 11645 10342 11679
rect 10701 11645 10735 11679
rect 12449 11645 12483 11679
rect 13001 11645 13035 11679
rect 15888 11645 15922 11679
rect 15991 11645 16025 11679
rect 16900 11645 16934 11679
rect 19108 11645 19142 11679
rect 8217 11577 8251 11611
rect 17325 11577 17359 11611
rect 7803 11509 7837 11543
rect 17003 11509 17037 11543
rect 18061 11509 18095 11543
rect 18889 11509 18923 11543
rect 19211 11509 19245 11543
rect 19717 11509 19751 11543
rect 12633 11305 12667 11339
rect 19809 11305 19843 11339
rect 16405 11237 16439 11271
rect 7941 11169 7975 11203
rect 12516 11169 12550 11203
rect 19625 11169 19659 11203
rect 1409 11101 1443 11135
rect 17969 11101 18003 11135
rect 18613 11101 18647 11135
rect 8125 11033 8159 11067
rect 16957 11033 16991 11067
rect 8401 10761 8435 10795
rect 12909 10761 12943 10795
rect 16313 10761 16347 10795
rect 18245 10761 18279 10795
rect 19625 10761 19659 10795
rect 15945 10693 15979 10727
rect 20177 10693 20211 10727
rect 7757 10625 7791 10659
rect 16497 10625 16531 10659
rect 16957 10625 16991 10659
rect 17785 10625 17819 10659
rect 18521 10625 18555 10659
rect 18797 10625 18831 10659
rect 1444 10557 1478 10591
rect 1869 10557 1903 10591
rect 2456 10557 2490 10591
rect 2881 10557 2915 10591
rect 19993 10557 20027 10591
rect 20545 10557 20579 10591
rect 1547 10489 1581 10523
rect 7297 10489 7331 10523
rect 7481 10489 7515 10523
rect 2559 10421 2593 10455
rect 12449 10421 12483 10455
rect 5641 10217 5675 10251
rect 8263 10217 8297 10251
rect 7297 10149 7331 10183
rect 12817 10149 12851 10183
rect 5457 10081 5491 10115
rect 8125 10081 8159 10115
rect 1593 10013 1627 10047
rect 6653 10013 6687 10047
rect 13093 10013 13127 10047
rect 17325 10013 17359 10047
rect 18429 10013 18463 10047
rect 18705 10013 18739 10047
rect 2145 9945 2179 9979
rect 2881 9673 2915 9707
rect 5871 9673 5905 9707
rect 6653 9673 6687 9707
rect 8125 9673 8159 9707
rect 12817 9673 12851 9707
rect 19073 9673 19107 9707
rect 19809 9673 19843 9707
rect 2145 9605 2179 9639
rect 5549 9605 5583 9639
rect 8723 9605 8757 9639
rect 18705 9605 18739 9639
rect 3157 9537 3191 9571
rect 3433 9537 3467 9571
rect 7113 9537 7147 9571
rect 13645 9537 13679 9571
rect 5800 9469 5834 9503
rect 8652 9469 8686 9503
rect 9632 9469 9666 9503
rect 10057 9469 10091 9503
rect 16440 9469 16474 9503
rect 16865 9469 16899 9503
rect 19625 9469 19659 9503
rect 20177 9469 20211 9503
rect 1593 9401 1627 9435
rect 7757 9401 7791 9435
rect 13185 9401 13219 9435
rect 13369 9401 13403 9435
rect 18153 9401 18187 9435
rect 6285 9333 6319 9367
rect 9045 9333 9079 9367
rect 9735 9333 9769 9367
rect 16543 9333 16577 9367
rect 17785 9333 17819 9367
rect 1961 9129 1995 9163
rect 7113 9129 7147 9163
rect 19763 9129 19797 9163
rect 2237 9061 2271 9095
rect 6469 9061 6503 9095
rect 7389 9061 7423 9095
rect 16589 9061 16623 9095
rect 4112 8993 4146 9027
rect 9724 8993 9758 9027
rect 12392 8993 12426 9027
rect 19660 8993 19694 9027
rect 2697 8925 2731 8959
rect 5825 8925 5859 8959
rect 7757 8925 7791 8959
rect 12495 8925 12529 8959
rect 13461 8925 13495 8959
rect 14105 8925 14139 8959
rect 18153 8925 18187 8959
rect 17141 8857 17175 8891
rect 18705 8857 18739 8891
rect 1685 8789 1719 8823
rect 4215 8789 4249 8823
rect 9827 8789 9861 8823
rect 2789 8585 2823 8619
rect 7389 8585 7423 8619
rect 9505 8585 9539 8619
rect 12633 8585 12667 8619
rect 13461 8585 13495 8619
rect 16313 8585 16347 8619
rect 19441 8585 19475 8619
rect 1685 8449 1719 8483
rect 1869 8449 1903 8483
rect 4537 8449 4571 8483
rect 7757 8449 7791 8483
rect 8677 8449 8711 8483
rect 9965 8449 9999 8483
rect 14381 8449 14415 8483
rect 17141 8449 17175 8483
rect 17509 8449 17543 8483
rect 18429 8449 18463 8483
rect 19993 8449 20027 8483
rect 2513 8313 2547 8347
rect 3709 8313 3743 8347
rect 4261 8313 4295 8347
rect 8401 8313 8435 8347
rect 9137 8313 9171 8347
rect 9689 8313 9723 8347
rect 13921 8313 13955 8347
rect 14105 8313 14139 8347
rect 16497 8313 16531 8347
rect 18153 8313 18187 8347
rect 19717 8313 19751 8347
rect 3985 8245 4019 8279
rect 5733 8245 5767 8279
rect 17785 8245 17819 8279
rect 19073 8245 19107 8279
rect 4859 8041 4893 8075
rect 11391 8041 11425 8075
rect 15439 8041 15473 8075
rect 16773 8041 16807 8075
rect 1869 7973 1903 8007
rect 2513 7973 2547 8007
rect 4629 7905 4663 7939
rect 11288 7905 11322 7939
rect 12760 7905 12794 7939
rect 15368 7905 15402 7939
rect 17785 7905 17819 7939
rect 7665 7837 7699 7871
rect 7941 7837 7975 7871
rect 9781 7837 9815 7871
rect 10057 7837 10091 7871
rect 18889 7837 18923 7871
rect 19165 7837 19199 7871
rect 12863 7701 12897 7735
rect 16405 7701 16439 7735
rect 17923 7701 17957 7735
rect 1547 7497 1581 7531
rect 4629 7497 4663 7531
rect 10333 7497 10367 7531
rect 11713 7497 11747 7531
rect 12725 7497 12759 7531
rect 16497 7497 16531 7531
rect 17877 7497 17911 7531
rect 18705 7497 18739 7531
rect 8401 7429 8435 7463
rect 9965 7429 9999 7463
rect 16129 7429 16163 7463
rect 2789 7361 2823 7395
rect 4261 7361 4295 7395
rect 4813 7361 4847 7395
rect 5457 7361 5491 7395
rect 9229 7361 9263 7395
rect 9413 7361 9447 7395
rect 12265 7361 12299 7395
rect 13001 7361 13035 7395
rect 19533 7361 19567 7395
rect 1476 7293 1510 7327
rect 1869 7293 1903 7327
rect 10920 7293 10954 7327
rect 11345 7293 11379 7327
rect 15945 7293 15979 7327
rect 18188 7293 18222 7327
rect 2513 7225 2547 7259
rect 7665 7225 7699 7259
rect 7849 7225 7883 7259
rect 13645 7225 13679 7259
rect 18291 7225 18325 7259
rect 19257 7225 19291 7259
rect 2237 7157 2271 7191
rect 7297 7157 7331 7191
rect 11023 7157 11057 7191
rect 15393 7157 15427 7191
rect 18981 7157 19015 7191
rect 1409 6953 1443 6987
rect 7573 6953 7607 6987
rect 8723 6953 8757 6987
rect 16267 6953 16301 6987
rect 18889 6953 18923 6987
rect 1961 6885 1995 6919
rect 4169 6885 4203 6919
rect 11345 6885 11379 6919
rect 19257 6885 19291 6919
rect 2421 6817 2455 6851
rect 8652 6817 8686 6851
rect 12884 6817 12918 6851
rect 13896 6817 13930 6851
rect 16196 6817 16230 6851
rect 5733 6749 5767 6783
rect 9781 6749 9815 6783
rect 11989 6749 12023 6783
rect 17693 6749 17727 6783
rect 19533 6749 19567 6783
rect 4721 6681 4755 6715
rect 6285 6681 6319 6715
rect 18245 6681 18279 6715
rect 2559 6613 2593 6647
rect 2881 6613 2915 6647
rect 12955 6613 12989 6647
rect 13967 6613 14001 6647
rect 2513 6409 2547 6443
rect 4169 6409 4203 6443
rect 11253 6409 11287 6443
rect 12909 6409 12943 6443
rect 17693 6409 17727 6443
rect 18199 6409 18233 6443
rect 20085 6409 20119 6443
rect 2237 6341 2271 6375
rect 5733 6341 5767 6375
rect 2789 6273 2823 6307
rect 4583 6273 4617 6307
rect 8585 6273 8619 6307
rect 13277 6273 13311 6307
rect 13461 6273 13495 6307
rect 13737 6273 13771 6307
rect 19441 6273 19475 6307
rect 1736 6205 1770 6239
rect 4496 6205 4530 6239
rect 18128 6205 18162 6239
rect 1823 6137 1857 6171
rect 3433 6137 3467 6171
rect 8309 6137 8343 6171
rect 10149 6137 10183 6171
rect 10793 6137 10827 6171
rect 18981 6137 19015 6171
rect 19165 6137 19199 6171
rect 4997 6069 5031 6103
rect 8033 6069 8067 6103
rect 9229 6069 9263 6103
rect 9873 6069 9907 6103
rect 14473 6069 14507 6103
rect 16221 6069 16255 6103
rect 18613 6069 18647 6103
rect 7711 5865 7745 5899
rect 8723 5865 8757 5899
rect 2789 5797 2823 5831
rect 5273 5797 5307 5831
rect 10149 5797 10183 5831
rect 11713 5797 11747 5831
rect 6596 5729 6630 5763
rect 7640 5729 7674 5763
rect 8620 5729 8654 5763
rect 13220 5729 13254 5763
rect 15828 5729 15862 5763
rect 2145 5661 2179 5695
rect 4629 5661 4663 5695
rect 10793 5661 10827 5695
rect 11989 5661 12023 5695
rect 17877 5661 17911 5695
rect 18981 5661 19015 5695
rect 19441 5661 19475 5695
rect 6699 5525 6733 5559
rect 13323 5525 13357 5559
rect 15899 5525 15933 5559
rect 1547 5321 1581 5355
rect 2237 5321 2271 5355
rect 3617 5321 3651 5355
rect 6561 5321 6595 5355
rect 9137 5321 9171 5355
rect 9873 5321 9907 5355
rect 11069 5321 11103 5355
rect 11713 5321 11747 5355
rect 13461 5321 13495 5355
rect 16681 5321 16715 5355
rect 19717 5321 19751 5355
rect 3157 5253 3191 5287
rect 19441 5253 19475 5287
rect 1869 5185 1903 5219
rect 2835 5185 2869 5219
rect 6193 5185 6227 5219
rect 6929 5185 6963 5219
rect 10149 5185 10183 5219
rect 10425 5185 10459 5219
rect 12265 5185 12299 5219
rect 12541 5185 12575 5219
rect 12817 5185 12851 5219
rect 15485 5185 15519 5219
rect 15669 5185 15703 5219
rect 19027 5185 19061 5219
rect 1476 5117 1510 5151
rect 2748 5117 2782 5151
rect 5432 5117 5466 5151
rect 8744 5117 8778 5151
rect 14080 5117 14114 5151
rect 14473 5117 14507 5151
rect 18940 5117 18974 5151
rect 3893 5049 3927 5083
rect 4537 5049 4571 5083
rect 7573 5049 7607 5083
rect 16313 5049 16347 5083
rect 4813 4981 4847 5015
rect 5503 4981 5537 5015
rect 5825 4981 5859 5015
rect 7849 4981 7883 5015
rect 8815 4981 8849 5015
rect 9505 4981 9539 5015
rect 14151 4981 14185 5015
rect 3111 4777 3145 4811
rect 6101 4709 6135 4743
rect 7665 4709 7699 4743
rect 10425 4709 10459 4743
rect 12633 4709 12667 4743
rect 12909 4709 12943 4743
rect 15393 4709 15427 4743
rect 16037 4709 16071 4743
rect 19993 4709 20027 4743
rect 16900 4641 16934 4675
rect 2881 4573 2915 4607
rect 4537 4573 4571 4607
rect 6377 4573 6411 4607
rect 7941 4573 7975 4607
rect 9781 4573 9815 4607
rect 11989 4573 12023 4607
rect 13461 4573 13495 4607
rect 19349 4573 19383 4607
rect 5089 4505 5123 4539
rect 17003 4437 17037 4471
rect 4813 4233 4847 4267
rect 6193 4233 6227 4267
rect 8033 4233 8067 4267
rect 9689 4233 9723 4267
rect 11989 4233 12023 4267
rect 15393 4233 15427 4267
rect 19441 4233 19475 4267
rect 19763 4233 19797 4267
rect 4445 4165 4479 4199
rect 10885 4165 10919 4199
rect 1869 4097 1903 4131
rect 9045 4097 9079 4131
rect 12541 4097 12575 4131
rect 14473 4097 14507 4131
rect 19165 4097 19199 4131
rect 1476 4029 1510 4063
rect 7272 4029 7306 4063
rect 10701 4029 10735 4063
rect 11253 4029 11287 4063
rect 14080 4029 14114 4063
rect 18680 4029 18714 4063
rect 19692 4029 19726 4063
rect 3893 3961 3927 3995
rect 8585 3961 8619 3995
rect 8769 3961 8803 3995
rect 13185 3961 13219 3995
rect 15025 3961 15059 3995
rect 15761 3961 15795 3995
rect 16405 3961 16439 3995
rect 16865 3961 16899 3995
rect 1547 3893 1581 3927
rect 3065 3893 3099 3927
rect 3617 3893 3651 3927
rect 5733 3893 5767 3927
rect 7343 3893 7377 3927
rect 7757 3893 7791 3927
rect 14151 3893 14185 3927
rect 18751 3893 18785 3927
rect 20177 3893 20211 3927
rect 2145 3621 2179 3655
rect 7573 3621 7607 3655
rect 10425 3621 10459 3655
rect 4445 3553 4479 3587
rect 6377 3553 6411 3587
rect 11253 3553 11287 3587
rect 12357 3553 12391 3587
rect 13496 3553 13530 3587
rect 19660 3553 19694 3587
rect 2789 3485 2823 3519
rect 7849 3485 7883 3519
rect 9781 3485 9815 3519
rect 15393 3485 15427 3519
rect 15669 3485 15703 3519
rect 16957 3485 16991 3519
rect 17233 3485 17267 3519
rect 18429 3485 18463 3519
rect 12909 3417 12943 3451
rect 4583 3349 4617 3383
rect 4905 3349 4939 3383
rect 6561 3349 6595 3383
rect 11437 3349 11471 3383
rect 12541 3349 12575 3383
rect 13599 3349 13633 3383
rect 19763 3349 19797 3383
rect 2145 3145 2179 3179
rect 3479 3145 3513 3179
rect 6561 3145 6595 3179
rect 7849 3145 7883 3179
rect 10057 3145 10091 3179
rect 11253 3145 11287 3179
rect 13461 3145 13495 3179
rect 14519 3145 14553 3179
rect 15853 3145 15887 3179
rect 17509 3145 17543 3179
rect 2467 3077 2501 3111
rect 6193 3077 6227 3111
rect 11529 3077 11563 3111
rect 14933 3077 14967 3111
rect 15301 3077 15335 3111
rect 2881 3009 2915 3043
rect 4813 3009 4847 3043
rect 6929 3009 6963 3043
rect 12541 3009 12575 3043
rect 13185 3009 13219 3043
rect 16865 3009 16899 3043
rect 17877 3009 17911 3043
rect 18153 3009 18187 3043
rect 19717 3009 19751 3043
rect 19993 3009 20027 3043
rect 2396 2941 2430 2975
rect 3408 2941 3442 2975
rect 5457 2941 5491 2975
rect 10609 2941 10643 2975
rect 14448 2941 14482 2975
rect 15460 2941 15494 2975
rect 7573 2873 7607 2907
rect 9137 2873 9171 2907
rect 9781 2873 9815 2907
rect 12173 2873 12207 2907
rect 16313 2873 16347 2907
rect 16497 2873 16531 2907
rect 18797 2873 18831 2907
rect 3893 2805 3927 2839
rect 4537 2805 4571 2839
rect 8861 2805 8895 2839
rect 10793 2805 10827 2839
rect 15531 2805 15565 2839
rect 19533 2805 19567 2839
rect 2099 2601 2133 2635
rect 9413 2601 9447 2635
rect 11989 2601 12023 2635
rect 12173 2601 12207 2635
rect 16129 2601 16163 2635
rect 19625 2601 19659 2635
rect 3249 2533 3283 2567
rect 7389 2533 7423 2567
rect 7573 2533 7607 2567
rect 2028 2465 2062 2499
rect 3040 2465 3074 2499
rect 3433 2465 3467 2499
rect 4328 2465 4362 2499
rect 6009 2465 6043 2499
rect 8217 2465 8251 2499
rect 4997 2397 5031 2431
rect 5365 2397 5399 2431
rect 4399 2329 4433 2363
rect 5089 2329 5123 2363
rect 2513 2261 2547 2295
rect 4721 2261 4755 2295
rect 4997 2261 5031 2295
rect 11437 2465 11471 2499
rect 9505 2397 9539 2431
rect 9873 2397 9907 2431
rect 10149 2397 10183 2431
rect 11621 2329 11655 2363
rect 9413 2261 9447 2295
rect 13369 2533 13403 2567
rect 18153 2533 18187 2567
rect 18429 2533 18463 2567
rect 14248 2465 14282 2499
rect 14657 2465 14691 2499
rect 15485 2465 15519 2499
rect 16589 2465 16623 2499
rect 17141 2465 17175 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 12449 2397 12483 2431
rect 12725 2397 12759 2431
rect 14335 2397 14369 2431
rect 18797 2397 18831 2431
rect 16773 2329 16807 2363
rect 12173 2261 12207 2295
rect 15669 2261 15703 2295
rect 20085 2261 20119 2295
<< metal1 >>
rect 2774 24216 2780 24268
rect 2832 24256 2838 24268
rect 4062 24256 4068 24268
rect 2832 24228 4068 24256
rect 2832 24216 2838 24228
rect 4062 24216 4068 24228
rect 4120 24216 4126 24268
rect 5258 24216 5264 24268
rect 5316 24256 5322 24268
rect 7834 24256 7840 24268
rect 5316 24228 7840 24256
rect 5316 24216 5322 24228
rect 7834 24216 7840 24228
rect 7892 24216 7898 24268
rect 1104 22330 21436 22352
rect 1104 22278 8497 22330
rect 8549 22278 8561 22330
rect 8613 22278 8625 22330
rect 8677 22278 8689 22330
rect 8741 22278 16012 22330
rect 16064 22278 16076 22330
rect 16128 22278 16140 22330
rect 16192 22278 16204 22330
rect 16256 22278 21436 22330
rect 1104 22256 21436 22278
rect 14 22040 20 22092
rect 72 22080 78 22092
rect 15562 22080 15568 22092
rect 72 22052 15568 22080
rect 72 22040 78 22052
rect 15562 22040 15568 22052
rect 15620 22040 15626 22092
rect 19680 22083 19738 22089
rect 19680 22049 19692 22083
rect 19726 22080 19738 22083
rect 20162 22080 20168 22092
rect 19726 22052 20168 22080
rect 19726 22049 19738 22052
rect 19680 22043 19738 22049
rect 20162 22040 20168 22052
rect 20220 22040 20226 22092
rect 106 21972 112 22024
rect 164 22012 170 22024
rect 12986 22012 12992 22024
rect 164 21984 12992 22012
rect 164 21972 170 21984
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 19610 21836 19616 21888
rect 19668 21876 19674 21888
rect 19751 21879 19809 21885
rect 19751 21876 19763 21879
rect 19668 21848 19763 21876
rect 19668 21836 19674 21848
rect 19751 21845 19763 21848
rect 19797 21845 19809 21879
rect 19751 21839 19809 21845
rect 1104 21786 21436 21808
rect 1104 21734 4739 21786
rect 4791 21734 4803 21786
rect 4855 21734 4867 21786
rect 4919 21734 4931 21786
rect 4983 21734 12255 21786
rect 12307 21734 12319 21786
rect 12371 21734 12383 21786
rect 12435 21734 12447 21786
rect 12499 21734 19770 21786
rect 19822 21734 19834 21786
rect 19886 21734 19898 21786
rect 19950 21734 19962 21786
rect 20014 21734 21436 21786
rect 1104 21712 21436 21734
rect 17405 21675 17463 21681
rect 17405 21641 17417 21675
rect 17451 21672 17463 21675
rect 18414 21672 18420 21684
rect 17451 21644 18420 21672
rect 17451 21641 17463 21644
rect 17405 21635 17463 21641
rect 10318 21496 10324 21548
rect 10376 21536 10382 21548
rect 10962 21536 10968 21548
rect 10376 21508 10968 21536
rect 10376 21496 10382 21508
rect 10962 21496 10968 21508
rect 11020 21536 11026 21548
rect 11020 21508 16804 21536
rect 11020 21496 11026 21508
rect 15562 21428 15568 21480
rect 15620 21468 15626 21480
rect 15876 21471 15934 21477
rect 15876 21468 15888 21471
rect 15620 21440 15888 21468
rect 15620 21428 15626 21440
rect 15876 21437 15888 21440
rect 15922 21468 15934 21471
rect 16301 21471 16359 21477
rect 16301 21468 16313 21471
rect 15922 21440 16313 21468
rect 15922 21437 15934 21440
rect 15876 21431 15934 21437
rect 16301 21437 16313 21440
rect 16347 21437 16359 21471
rect 16301 21431 16359 21437
rect 14369 21403 14427 21409
rect 14369 21369 14381 21403
rect 14415 21369 14427 21403
rect 15010 21400 15016 21412
rect 14971 21372 15016 21400
rect 14369 21363 14427 21369
rect 14090 21332 14096 21344
rect 14051 21304 14096 21332
rect 14090 21292 14096 21304
rect 14148 21332 14154 21344
rect 14384 21332 14412 21363
rect 15010 21360 15016 21372
rect 15068 21360 15074 21412
rect 16776 21400 16804 21508
rect 16920 21471 16978 21477
rect 16920 21437 16932 21471
rect 16966 21468 16978 21471
rect 17420 21468 17448 21635
rect 18414 21632 18420 21644
rect 18472 21632 18478 21684
rect 19705 21675 19763 21681
rect 19705 21641 19717 21675
rect 19751 21672 19763 21675
rect 20162 21672 20168 21684
rect 19751 21644 20168 21672
rect 19751 21641 19763 21644
rect 19705 21635 19763 21641
rect 20162 21632 20168 21644
rect 20220 21632 20226 21684
rect 20349 21675 20407 21681
rect 20349 21641 20361 21675
rect 20395 21672 20407 21675
rect 21542 21672 21548 21684
rect 20395 21644 21548 21672
rect 20395 21641 20407 21644
rect 20349 21635 20407 21641
rect 18877 21607 18935 21613
rect 18877 21573 18889 21607
rect 18923 21604 18935 21607
rect 20254 21604 20260 21616
rect 18923 21576 20260 21604
rect 18923 21573 18935 21576
rect 18877 21567 18935 21573
rect 20254 21564 20260 21576
rect 20312 21564 20318 21616
rect 16966 21440 17448 21468
rect 18693 21471 18751 21477
rect 16966 21437 16978 21440
rect 16920 21431 16978 21437
rect 18693 21437 18705 21471
rect 18739 21468 18751 21471
rect 19245 21471 19303 21477
rect 19245 21468 19257 21471
rect 18739 21440 19257 21468
rect 18739 21437 18751 21440
rect 18693 21431 18751 21437
rect 19245 21437 19257 21440
rect 19291 21437 19303 21471
rect 19245 21431 19303 21437
rect 19864 21471 19922 21477
rect 19864 21437 19876 21471
rect 19910 21468 19922 21471
rect 20364 21468 20392 21635
rect 21542 21632 21548 21644
rect 21600 21632 21606 21684
rect 19910 21440 20392 21468
rect 19910 21437 19922 21440
rect 19864 21431 19922 21437
rect 18708 21400 18736 21431
rect 16776 21372 18736 21400
rect 14148 21304 14412 21332
rect 15979 21335 16037 21341
rect 14148 21292 14154 21304
rect 15979 21301 15991 21335
rect 16025 21332 16037 21335
rect 16298 21332 16304 21344
rect 16025 21304 16304 21332
rect 16025 21301 16037 21304
rect 15979 21295 16037 21301
rect 16298 21292 16304 21304
rect 16356 21292 16362 21344
rect 16390 21292 16396 21344
rect 16448 21332 16454 21344
rect 16991 21335 17049 21341
rect 16991 21332 17003 21335
rect 16448 21304 17003 21332
rect 16448 21292 16454 21304
rect 16991 21301 17003 21304
rect 17037 21301 17049 21335
rect 16991 21295 17049 21301
rect 19702 21292 19708 21344
rect 19760 21332 19766 21344
rect 19935 21335 19993 21341
rect 19935 21332 19947 21335
rect 19760 21304 19947 21332
rect 19760 21292 19766 21304
rect 19935 21301 19947 21304
rect 19981 21301 19993 21335
rect 19935 21295 19993 21301
rect 1104 21242 21436 21264
rect 1104 21190 8497 21242
rect 8549 21190 8561 21242
rect 8613 21190 8625 21242
rect 8677 21190 8689 21242
rect 8741 21190 16012 21242
rect 16064 21190 16076 21242
rect 16128 21190 16140 21242
rect 16192 21190 16204 21242
rect 16256 21190 21436 21242
rect 1104 21168 21436 21190
rect 8665 21131 8723 21137
rect 8665 21097 8677 21131
rect 8711 21128 8723 21131
rect 8938 21128 8944 21140
rect 8711 21100 8944 21128
rect 8711 21097 8723 21100
rect 8665 21091 8723 21097
rect 8938 21088 8944 21100
rect 8996 21088 9002 21140
rect 12066 21088 12072 21140
rect 12124 21128 12130 21140
rect 12345 21131 12403 21137
rect 12345 21128 12357 21131
rect 12124 21100 12357 21128
rect 12124 21088 12130 21100
rect 12345 21097 12357 21100
rect 12391 21097 12403 21131
rect 12345 21091 12403 21097
rect 14826 21060 14832 21072
rect 12176 21032 14832 21060
rect 1464 20995 1522 21001
rect 1464 20961 1476 20995
rect 1510 20992 1522 20995
rect 1578 20992 1584 21004
rect 1510 20964 1584 20992
rect 1510 20961 1522 20964
rect 1464 20955 1522 20961
rect 1578 20952 1584 20964
rect 1636 20952 1642 21004
rect 8481 20995 8539 21001
rect 8481 20961 8493 20995
rect 8527 20961 8539 20995
rect 9582 20992 9588 21004
rect 9543 20964 9588 20992
rect 8481 20955 8539 20961
rect 8496 20924 8524 20955
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 12066 20952 12072 21004
rect 12124 20992 12130 21004
rect 12176 21001 12204 21032
rect 14826 21020 14832 21032
rect 14884 21020 14890 21072
rect 16301 21063 16359 21069
rect 16301 21029 16313 21063
rect 16347 21060 16359 21063
rect 16390 21060 16396 21072
rect 16347 21032 16396 21060
rect 16347 21029 16359 21032
rect 16301 21023 16359 21029
rect 16390 21020 16396 21032
rect 16448 21020 16454 21072
rect 19334 21060 19340 21072
rect 19247 21032 19340 21060
rect 19334 21020 19340 21032
rect 19392 21060 19398 21072
rect 19702 21060 19708 21072
rect 19392 21032 19708 21060
rect 19392 21020 19398 21032
rect 19702 21020 19708 21032
rect 19760 21020 19766 21072
rect 12161 20995 12219 21001
rect 12161 20992 12173 20995
rect 12124 20964 12173 20992
rect 12124 20952 12130 20964
rect 12161 20961 12173 20964
rect 12207 20961 12219 20995
rect 12161 20955 12219 20961
rect 12986 20952 12992 21004
rect 13044 20992 13050 21004
rect 13300 20995 13358 21001
rect 13300 20992 13312 20995
rect 13044 20964 13312 20992
rect 13044 20952 13050 20964
rect 13300 20961 13312 20964
rect 13346 20961 13358 20995
rect 13300 20955 13358 20961
rect 18300 20995 18358 21001
rect 18300 20961 18312 20995
rect 18346 20992 18358 20995
rect 18506 20992 18512 21004
rect 18346 20964 18512 20992
rect 18346 20961 18358 20964
rect 18300 20955 18358 20961
rect 18506 20952 18512 20964
rect 18564 20952 18570 21004
rect 8570 20924 8576 20936
rect 8483 20896 8576 20924
rect 8570 20884 8576 20896
rect 8628 20924 8634 20936
rect 9815 20927 9873 20933
rect 9815 20924 9827 20927
rect 8628 20896 9827 20924
rect 8628 20884 8634 20896
rect 9815 20893 9827 20896
rect 9861 20893 9873 20927
rect 16574 20924 16580 20936
rect 16535 20896 16580 20924
rect 9815 20887 9873 20893
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20924 20039 20927
rect 20070 20924 20076 20936
rect 20027 20896 20076 20924
rect 20027 20893 20039 20896
rect 19981 20887 20039 20893
rect 20070 20884 20076 20896
rect 20128 20884 20134 20936
rect 1535 20791 1593 20797
rect 1535 20757 1547 20791
rect 1581 20788 1593 20791
rect 1946 20788 1952 20800
rect 1581 20760 1952 20788
rect 1581 20757 1593 20760
rect 1535 20751 1593 20757
rect 1946 20748 1952 20760
rect 2004 20748 2010 20800
rect 13403 20791 13461 20797
rect 13403 20757 13415 20791
rect 13449 20788 13461 20791
rect 13906 20788 13912 20800
rect 13449 20760 13912 20788
rect 13449 20757 13461 20760
rect 13403 20751 13461 20757
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 18371 20791 18429 20797
rect 18371 20757 18383 20791
rect 18417 20788 18429 20791
rect 19518 20788 19524 20800
rect 18417 20760 19524 20788
rect 18417 20757 18429 20760
rect 18371 20751 18429 20757
rect 19518 20748 19524 20760
rect 19576 20748 19582 20800
rect 1104 20698 21436 20720
rect 1104 20646 4739 20698
rect 4791 20646 4803 20698
rect 4855 20646 4867 20698
rect 4919 20646 4931 20698
rect 4983 20646 12255 20698
rect 12307 20646 12319 20698
rect 12371 20646 12383 20698
rect 12435 20646 12447 20698
rect 12499 20646 19770 20698
rect 19822 20646 19834 20698
rect 19886 20646 19898 20698
rect 19950 20646 19962 20698
rect 20014 20646 21436 20698
rect 1104 20624 21436 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 1946 20584 1952 20596
rect 1907 20556 1952 20584
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 8570 20584 8576 20596
rect 8531 20556 8576 20584
rect 8570 20544 8576 20556
rect 8628 20544 8634 20596
rect 12986 20544 12992 20596
rect 13044 20584 13050 20596
rect 13265 20587 13323 20593
rect 13265 20584 13277 20587
rect 13044 20556 13277 20584
rect 13044 20544 13050 20556
rect 13265 20553 13277 20556
rect 13311 20553 13323 20587
rect 13906 20584 13912 20596
rect 13867 20556 13912 20584
rect 13265 20547 13323 20553
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 16390 20544 16396 20596
rect 16448 20584 16454 20596
rect 16669 20587 16727 20593
rect 16669 20584 16681 20587
rect 16448 20556 16681 20584
rect 16448 20544 16454 20556
rect 16669 20553 16681 20556
rect 16715 20553 16727 20587
rect 16669 20547 16727 20553
rect 18325 20587 18383 20593
rect 18325 20553 18337 20587
rect 18371 20584 18383 20587
rect 18506 20584 18512 20596
rect 18371 20556 18512 20584
rect 18371 20553 18383 20556
rect 18325 20547 18383 20553
rect 18506 20544 18512 20556
rect 18564 20544 18570 20596
rect 19334 20584 19340 20596
rect 19295 20556 19340 20584
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 1964 20448 1992 20544
rect 2225 20451 2283 20457
rect 2225 20448 2237 20451
rect 1964 20420 2237 20448
rect 2225 20417 2237 20420
rect 2271 20417 2283 20451
rect 13924 20448 13952 20544
rect 14737 20519 14795 20525
rect 14737 20485 14749 20519
rect 14783 20516 14795 20519
rect 17034 20516 17040 20528
rect 14783 20488 17040 20516
rect 14783 20485 14795 20488
rect 14737 20479 14795 20485
rect 17034 20476 17040 20488
rect 17092 20516 17098 20528
rect 17092 20488 19932 20516
rect 17092 20476 17098 20488
rect 14185 20451 14243 20457
rect 14185 20448 14197 20451
rect 13924 20420 14197 20448
rect 2225 20411 2283 20417
rect 14185 20417 14197 20420
rect 14231 20417 14243 20451
rect 14185 20411 14243 20417
rect 16393 20451 16451 20457
rect 16393 20417 16405 20451
rect 16439 20448 16451 20451
rect 16574 20448 16580 20460
rect 16439 20420 16580 20448
rect 16439 20417 16451 20420
rect 16393 20411 16451 20417
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 18969 20451 19027 20457
rect 18969 20417 18981 20451
rect 19015 20448 19027 20451
rect 19610 20448 19616 20460
rect 19015 20420 19616 20448
rect 19015 20417 19027 20420
rect 18969 20411 19027 20417
rect 19610 20408 19616 20420
rect 19668 20408 19674 20460
rect 19904 20457 19932 20488
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20417 19947 20451
rect 19889 20411 19947 20417
rect 2866 20312 2872 20324
rect 2827 20284 2872 20312
rect 2866 20272 2872 20284
rect 2924 20272 2930 20324
rect 9582 20272 9588 20324
rect 9640 20312 9646 20324
rect 9769 20315 9827 20321
rect 9769 20312 9781 20315
rect 9640 20284 9781 20312
rect 9640 20272 9646 20284
rect 9769 20281 9781 20284
rect 9815 20312 9827 20315
rect 15749 20315 15807 20321
rect 9815 20284 13814 20312
rect 9815 20281 9827 20284
rect 9769 20275 9827 20281
rect 12066 20204 12072 20256
rect 12124 20244 12130 20256
rect 12161 20247 12219 20253
rect 12161 20244 12173 20247
rect 12124 20216 12173 20244
rect 12124 20204 12130 20216
rect 12161 20213 12173 20216
rect 12207 20213 12219 20247
rect 13786 20244 13814 20284
rect 15749 20281 15761 20315
rect 15795 20281 15807 20315
rect 15749 20275 15807 20281
rect 15010 20244 15016 20256
rect 13786 20216 15016 20244
rect 12161 20207 12219 20213
rect 15010 20204 15016 20216
rect 15068 20204 15074 20256
rect 15470 20244 15476 20256
rect 15431 20216 15476 20244
rect 15470 20204 15476 20216
rect 15528 20244 15534 20256
rect 15764 20244 15792 20275
rect 15528 20216 15792 20244
rect 15528 20204 15534 20216
rect 1104 20154 21436 20176
rect 1104 20102 8497 20154
rect 8549 20102 8561 20154
rect 8613 20102 8625 20154
rect 8677 20102 8689 20154
rect 8741 20102 16012 20154
rect 16064 20102 16076 20154
rect 16128 20102 16140 20154
rect 16192 20102 16204 20154
rect 16256 20102 21436 20154
rect 1104 20080 21436 20102
rect 14090 20040 14096 20052
rect 14051 20012 14096 20040
rect 14090 20000 14096 20012
rect 14148 20000 14154 20052
rect 15010 19932 15016 19984
rect 15068 19972 15074 19984
rect 16025 19975 16083 19981
rect 16025 19972 16037 19975
rect 15068 19944 16037 19972
rect 15068 19932 15074 19944
rect 16025 19941 16037 19944
rect 16071 19941 16083 19975
rect 16025 19935 16083 19941
rect 16298 19932 16304 19984
rect 16356 19972 16362 19984
rect 16942 19972 16948 19984
rect 16356 19944 16948 19972
rect 16356 19932 16362 19944
rect 16942 19932 16948 19944
rect 17000 19932 17006 19984
rect 17589 19975 17647 19981
rect 17589 19941 17601 19975
rect 17635 19972 17647 19975
rect 17862 19972 17868 19984
rect 17635 19944 17868 19972
rect 17635 19941 17647 19944
rect 17589 19935 17647 19941
rect 17862 19932 17868 19944
rect 17920 19972 17926 19984
rect 19981 19975 20039 19981
rect 19981 19972 19993 19975
rect 17920 19944 19993 19972
rect 17920 19932 17926 19944
rect 19981 19941 19993 19944
rect 20027 19972 20039 19975
rect 20070 19972 20076 19984
rect 20027 19944 20076 19972
rect 20027 19941 20039 19944
rect 19981 19935 20039 19941
rect 20070 19932 20076 19944
rect 20128 19932 20134 19984
rect 15381 19839 15439 19845
rect 15381 19805 15393 19839
rect 15427 19836 15439 19839
rect 15838 19836 15844 19848
rect 15427 19808 15844 19836
rect 15427 19805 15439 19808
rect 15381 19799 15439 19805
rect 15838 19796 15844 19808
rect 15896 19836 15902 19848
rect 16574 19836 16580 19848
rect 15896 19808 16580 19836
rect 15896 19796 15902 19808
rect 16574 19796 16580 19808
rect 16632 19796 16638 19848
rect 19334 19836 19340 19848
rect 19295 19808 19340 19836
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 1104 19610 21436 19632
rect 1104 19558 4739 19610
rect 4791 19558 4803 19610
rect 4855 19558 4867 19610
rect 4919 19558 4931 19610
rect 4983 19558 12255 19610
rect 12307 19558 12319 19610
rect 12371 19558 12383 19610
rect 12435 19558 12447 19610
rect 12499 19558 19770 19610
rect 19822 19558 19834 19610
rect 19886 19558 19898 19610
rect 19950 19558 19962 19610
rect 20014 19558 21436 19610
rect 1104 19536 21436 19558
rect 15059 19499 15117 19505
rect 15059 19465 15071 19499
rect 15105 19496 15117 19499
rect 15470 19496 15476 19508
rect 15105 19468 15476 19496
rect 15105 19465 15117 19468
rect 15059 19459 15117 19465
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 15838 19496 15844 19508
rect 15799 19468 15844 19496
rect 15838 19456 15844 19468
rect 15896 19456 15902 19508
rect 16942 19496 16948 19508
rect 16903 19468 16948 19496
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 17862 19496 17868 19508
rect 17823 19468 17868 19496
rect 17862 19456 17868 19468
rect 17920 19456 17926 19508
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19360 15531 19363
rect 15654 19360 15660 19372
rect 15519 19332 15660 19360
rect 15519 19329 15531 19332
rect 15473 19323 15531 19329
rect 15010 19301 15016 19304
rect 14988 19295 15016 19301
rect 14988 19292 15000 19295
rect 14923 19264 15000 19292
rect 14988 19261 15000 19264
rect 15068 19292 15074 19304
rect 15488 19292 15516 19323
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 17880 19360 17908 19456
rect 18141 19363 18199 19369
rect 18141 19360 18153 19363
rect 17880 19332 18153 19360
rect 18141 19329 18153 19332
rect 18187 19329 18199 19363
rect 18414 19360 18420 19372
rect 18375 19332 18420 19360
rect 18141 19323 18199 19329
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 19518 19320 19524 19372
rect 19576 19360 19582 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19576 19332 19717 19360
rect 19576 19320 19582 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 15068 19264 15516 19292
rect 14988 19255 15016 19261
rect 15010 19252 15016 19255
rect 15068 19252 15074 19264
rect 19426 19184 19432 19236
rect 19484 19224 19490 19236
rect 20349 19227 20407 19233
rect 20349 19224 20361 19227
rect 19484 19196 20361 19224
rect 19484 19184 19490 19196
rect 20349 19193 20361 19196
rect 20395 19193 20407 19227
rect 20349 19187 20407 19193
rect 19334 19156 19340 19168
rect 19295 19128 19340 19156
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 1104 19066 21436 19088
rect 1104 19014 8497 19066
rect 8549 19014 8561 19066
rect 8613 19014 8625 19066
rect 8677 19014 8689 19066
rect 8741 19014 16012 19066
rect 16064 19014 16076 19066
rect 16128 19014 16140 19066
rect 16192 19014 16204 19066
rect 16256 19014 21436 19066
rect 1104 18992 21436 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 19751 18955 19809 18961
rect 19751 18952 19763 18955
rect 19392 18924 19763 18952
rect 19392 18912 19398 18924
rect 19751 18921 19763 18924
rect 19797 18921 19809 18955
rect 19751 18915 19809 18921
rect 19518 18844 19524 18896
rect 19576 18884 19582 18896
rect 20073 18887 20131 18893
rect 20073 18884 20085 18887
rect 19576 18856 20085 18884
rect 19576 18844 19582 18856
rect 20073 18853 20085 18856
rect 20119 18853 20131 18887
rect 20073 18847 20131 18853
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 6549 18819 6607 18825
rect 6549 18785 6561 18819
rect 6595 18816 6607 18819
rect 6638 18816 6644 18828
rect 6595 18788 6644 18816
rect 6595 18785 6607 18788
rect 6549 18779 6607 18785
rect 6638 18776 6644 18788
rect 6696 18776 6702 18828
rect 19680 18819 19738 18825
rect 19680 18785 19692 18819
rect 19726 18816 19738 18819
rect 20346 18816 20352 18828
rect 19726 18788 20352 18816
rect 19726 18785 19738 18788
rect 19680 18779 19738 18785
rect 20346 18776 20352 18788
rect 20404 18776 20410 18828
rect 6086 18572 6092 18624
rect 6144 18612 6150 18624
rect 6687 18615 6745 18621
rect 6687 18612 6699 18615
rect 6144 18584 6699 18612
rect 6144 18572 6150 18584
rect 6687 18581 6699 18584
rect 6733 18581 6745 18615
rect 6687 18575 6745 18581
rect 1104 18522 21436 18544
rect 1104 18470 4739 18522
rect 4791 18470 4803 18522
rect 4855 18470 4867 18522
rect 4919 18470 4931 18522
rect 4983 18470 12255 18522
rect 12307 18470 12319 18522
rect 12371 18470 12383 18522
rect 12435 18470 12447 18522
rect 12499 18470 19770 18522
rect 19822 18470 19834 18522
rect 19886 18470 19898 18522
rect 19950 18470 19962 18522
rect 20014 18470 21436 18522
rect 1104 18448 21436 18470
rect 1394 18368 1400 18420
rect 1452 18408 1458 18420
rect 1581 18411 1639 18417
rect 1581 18408 1593 18411
rect 1452 18380 1593 18408
rect 1452 18368 1458 18380
rect 1581 18377 1593 18380
rect 1627 18377 1639 18411
rect 7466 18408 7472 18420
rect 7427 18380 7472 18408
rect 1581 18371 1639 18377
rect 7466 18368 7472 18380
rect 7524 18368 7530 18420
rect 19705 18411 19763 18417
rect 19705 18377 19717 18411
rect 19751 18408 19763 18411
rect 20346 18408 20352 18420
rect 19751 18380 20352 18408
rect 19751 18377 19763 18380
rect 19705 18371 19763 18377
rect 20346 18368 20352 18380
rect 20404 18368 20410 18420
rect 6638 18272 6644 18284
rect 6551 18244 6644 18272
rect 6638 18232 6644 18244
rect 6696 18272 6702 18284
rect 11698 18272 11704 18284
rect 6696 18244 11704 18272
rect 6696 18232 6702 18244
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 7098 18164 7104 18216
rect 7156 18204 7162 18216
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 7156 18176 7297 18204
rect 7156 18164 7162 18176
rect 7285 18173 7297 18176
rect 7331 18204 7343 18207
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7331 18176 7849 18204
rect 7331 18173 7343 18176
rect 7285 18167 7343 18173
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 8389 18207 8447 18213
rect 8389 18173 8401 18207
rect 8435 18204 8447 18207
rect 8435 18176 9076 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 8573 18071 8631 18077
rect 8573 18037 8585 18071
rect 8619 18068 8631 18071
rect 8846 18068 8852 18080
rect 8619 18040 8852 18068
rect 8619 18037 8631 18040
rect 8573 18031 8631 18037
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 9048 18077 9076 18176
rect 9033 18071 9091 18077
rect 9033 18037 9045 18071
rect 9079 18068 9091 18071
rect 9490 18068 9496 18080
rect 9079 18040 9496 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 1104 17978 21436 18000
rect 1104 17926 8497 17978
rect 8549 17926 8561 17978
rect 8613 17926 8625 17978
rect 8677 17926 8689 17978
rect 8741 17926 16012 17978
rect 16064 17926 16076 17978
rect 16128 17926 16140 17978
rect 16192 17926 16204 17978
rect 16256 17926 21436 17978
rect 1104 17904 21436 17926
rect 1394 17824 1400 17876
rect 1452 17864 1458 17876
rect 1811 17867 1869 17873
rect 1811 17864 1823 17867
rect 1452 17836 1823 17864
rect 1452 17824 1458 17836
rect 1811 17833 1823 17836
rect 1857 17833 1869 17867
rect 6270 17864 6276 17876
rect 6231 17836 6276 17864
rect 1811 17827 1869 17833
rect 6270 17824 6276 17836
rect 6328 17824 6334 17876
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17728 1731 17731
rect 1762 17728 1768 17740
rect 1719 17700 1768 17728
rect 1719 17697 1731 17700
rect 1673 17691 1731 17697
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 6086 17728 6092 17740
rect 6047 17700 6092 17728
rect 6086 17688 6092 17700
rect 6144 17688 6150 17740
rect 7650 17660 7656 17672
rect 7611 17632 7656 17660
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 1104 17434 21436 17456
rect 1104 17382 4739 17434
rect 4791 17382 4803 17434
rect 4855 17382 4867 17434
rect 4919 17382 4931 17434
rect 4983 17382 12255 17434
rect 12307 17382 12319 17434
rect 12371 17382 12383 17434
rect 12435 17382 12447 17434
rect 12499 17382 19770 17434
rect 19822 17382 19834 17434
rect 19886 17382 19898 17434
rect 19950 17382 19962 17434
rect 20014 17382 21436 17434
rect 1104 17360 21436 17382
rect 2866 17280 2872 17332
rect 2924 17320 2930 17332
rect 3053 17323 3111 17329
rect 3053 17320 3065 17323
rect 2924 17292 3065 17320
rect 2924 17280 2930 17292
rect 3053 17289 3065 17292
rect 3099 17289 3111 17323
rect 6086 17320 6092 17332
rect 6047 17292 6092 17320
rect 3053 17283 3111 17289
rect 3068 17184 3096 17283
rect 6086 17280 6092 17292
rect 6144 17280 6150 17332
rect 7098 17320 7104 17332
rect 7059 17292 7104 17320
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 7650 17320 7656 17332
rect 7611 17292 7656 17320
rect 7650 17280 7656 17292
rect 7708 17320 7714 17332
rect 7708 17292 7972 17320
rect 7708 17280 7714 17292
rect 3329 17187 3387 17193
rect 3329 17184 3341 17187
rect 3068 17156 3341 17184
rect 3329 17153 3341 17156
rect 3375 17184 3387 17187
rect 7742 17184 7748 17196
rect 3375 17156 7748 17184
rect 3375 17153 3387 17156
rect 3329 17147 3387 17153
rect 7742 17144 7748 17156
rect 7800 17144 7806 17196
rect 7944 17193 7972 17292
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17153 7987 17187
rect 8386 17184 8392 17196
rect 8347 17156 8392 17184
rect 7929 17147 7987 17153
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 6892 17119 6950 17125
rect 6892 17085 6904 17119
rect 6938 17116 6950 17119
rect 6938 17088 7420 17116
rect 6938 17085 6950 17088
rect 6892 17079 6950 17085
rect 3973 17051 4031 17057
rect 3973 17048 3985 17051
rect 2700 17020 3985 17048
rect 2700 16992 2728 17020
rect 3973 17017 3985 17020
rect 4019 17017 4031 17051
rect 3973 17011 4031 17017
rect 1762 16980 1768 16992
rect 1675 16952 1768 16980
rect 1762 16940 1768 16952
rect 1820 16980 1826 16992
rect 2682 16980 2688 16992
rect 1820 16952 2688 16980
rect 1820 16940 1826 16952
rect 2682 16940 2688 16952
rect 2740 16940 2746 16992
rect 7392 16989 7420 17088
rect 7377 16983 7435 16989
rect 7377 16949 7389 16983
rect 7423 16980 7435 16983
rect 8386 16980 8392 16992
rect 7423 16952 8392 16980
rect 7423 16949 7435 16952
rect 7377 16943 7435 16949
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 1104 16890 21436 16912
rect 1104 16838 8497 16890
rect 8549 16838 8561 16890
rect 8613 16838 8625 16890
rect 8677 16838 8689 16890
rect 8741 16838 16012 16890
rect 16064 16838 16076 16890
rect 16128 16838 16140 16890
rect 16192 16838 16204 16890
rect 16256 16838 21436 16890
rect 1104 16816 21436 16838
rect 9861 16779 9919 16785
rect 9861 16745 9873 16779
rect 9907 16776 9919 16779
rect 19242 16776 19248 16788
rect 9907 16748 19248 16776
rect 9907 16745 9919 16748
rect 9861 16739 9919 16745
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 19794 16776 19800 16788
rect 19755 16748 19800 16776
rect 19794 16736 19800 16748
rect 19852 16736 19858 16788
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19613 16643 19671 16649
rect 19613 16640 19625 16643
rect 19484 16612 19625 16640
rect 19484 16600 19490 16612
rect 19613 16609 19625 16612
rect 19659 16609 19671 16643
rect 19613 16603 19671 16609
rect 8110 16572 8116 16584
rect 8071 16544 8116 16572
rect 8110 16532 8116 16544
rect 8168 16532 8174 16584
rect 8386 16572 8392 16584
rect 8347 16544 8392 16572
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 1104 16346 21436 16368
rect 1104 16294 4739 16346
rect 4791 16294 4803 16346
rect 4855 16294 4867 16346
rect 4919 16294 4931 16346
rect 4983 16294 12255 16346
rect 12307 16294 12319 16346
rect 12371 16294 12383 16346
rect 12435 16294 12447 16346
rect 12499 16294 19770 16346
rect 19822 16294 19834 16346
rect 19886 16294 19898 16346
rect 19950 16294 19962 16346
rect 20014 16294 21436 16346
rect 1104 16272 21436 16294
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 19576 16068 19993 16096
rect 19576 16056 19582 16068
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 8018 15960 8024 15972
rect 7931 15932 8024 15960
rect 8018 15920 8024 15932
rect 8076 15960 8082 15972
rect 8205 15963 8263 15969
rect 8205 15960 8217 15963
rect 8076 15932 8217 15960
rect 8076 15920 8082 15932
rect 8205 15929 8217 15932
rect 8251 15929 8263 15963
rect 8205 15923 8263 15929
rect 8849 15963 8907 15969
rect 8849 15929 8861 15963
rect 8895 15960 8907 15963
rect 9122 15960 9128 15972
rect 8895 15932 9128 15960
rect 8895 15929 8907 15932
rect 8849 15923 8907 15929
rect 7653 15895 7711 15901
rect 7653 15861 7665 15895
rect 7699 15892 7711 15895
rect 8110 15892 8116 15904
rect 7699 15864 8116 15892
rect 7699 15861 7711 15864
rect 7653 15855 7711 15861
rect 8110 15852 8116 15864
rect 8168 15892 8174 15904
rect 8864 15892 8892 15923
rect 9122 15920 9128 15932
rect 9180 15920 9186 15972
rect 19153 15963 19211 15969
rect 19153 15929 19165 15963
rect 19199 15960 19211 15963
rect 19518 15960 19524 15972
rect 19199 15932 19524 15960
rect 19199 15929 19211 15932
rect 19153 15923 19211 15929
rect 19518 15920 19524 15932
rect 19576 15960 19582 15972
rect 19705 15963 19763 15969
rect 19705 15960 19717 15963
rect 19576 15932 19717 15960
rect 19576 15920 19582 15932
rect 19705 15929 19717 15932
rect 19751 15929 19763 15963
rect 19705 15923 19763 15929
rect 9674 15892 9680 15904
rect 8168 15864 8892 15892
rect 9635 15864 9680 15892
rect 8168 15852 8174 15864
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 19426 15892 19432 15904
rect 19387 15864 19432 15892
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 1104 15802 21436 15824
rect 1104 15750 8497 15802
rect 8549 15750 8561 15802
rect 8613 15750 8625 15802
rect 8677 15750 8689 15802
rect 8741 15750 16012 15802
rect 16064 15750 16076 15802
rect 16128 15750 16140 15802
rect 16192 15750 16204 15802
rect 16256 15750 21436 15802
rect 1104 15728 21436 15750
rect 7883 15691 7941 15697
rect 7883 15657 7895 15691
rect 7929 15688 7941 15691
rect 8018 15688 8024 15700
rect 7929 15660 8024 15688
rect 7929 15657 7941 15660
rect 7883 15651 7941 15657
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 19518 15580 19524 15632
rect 19576 15620 19582 15632
rect 19751 15623 19809 15629
rect 19751 15620 19763 15623
rect 19576 15592 19763 15620
rect 19576 15580 19582 15592
rect 19751 15589 19763 15592
rect 19797 15589 19809 15623
rect 19751 15583 19809 15589
rect 7374 15512 7380 15564
rect 7432 15552 7438 15564
rect 7780 15555 7838 15561
rect 7780 15552 7792 15555
rect 7432 15524 7792 15552
rect 7432 15512 7438 15524
rect 7780 15521 7792 15524
rect 7826 15552 7838 15555
rect 9674 15552 9680 15564
rect 7826 15524 9680 15552
rect 7826 15521 7838 15524
rect 7780 15515 7838 15521
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 19664 15555 19722 15561
rect 19664 15521 19676 15555
rect 19710 15552 19722 15555
rect 20070 15552 20076 15564
rect 19710 15524 20076 15552
rect 19710 15521 19722 15524
rect 19664 15515 19722 15521
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 1104 15258 21436 15280
rect 1104 15206 4739 15258
rect 4791 15206 4803 15258
rect 4855 15206 4867 15258
rect 4919 15206 4931 15258
rect 4983 15206 12255 15258
rect 12307 15206 12319 15258
rect 12371 15206 12383 15258
rect 12435 15206 12447 15258
rect 12499 15206 19770 15258
rect 19822 15206 19834 15258
rect 19886 15206 19898 15258
rect 19950 15206 19962 15258
rect 20014 15206 21436 15258
rect 1104 15184 21436 15206
rect 14550 15144 14556 15156
rect 14511 15116 14556 15144
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 15010 15144 15016 15156
rect 14971 15116 15016 15144
rect 15010 15104 15016 15116
rect 15068 15144 15074 15156
rect 15933 15147 15991 15153
rect 15933 15144 15945 15147
rect 15068 15116 15945 15144
rect 15068 15104 15074 15116
rect 9122 15008 9128 15020
rect 9083 14980 9128 15008
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 15555 14949 15583 15116
rect 15933 15113 15945 15116
rect 15979 15113 15991 15147
rect 15933 15107 15991 15113
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 19567 15147 19625 15153
rect 19567 15144 19579 15147
rect 19484 15116 19579 15144
rect 19484 15104 19490 15116
rect 19567 15113 19579 15116
rect 19613 15113 19625 15147
rect 19567 15107 19625 15113
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14940 14427 14943
rect 15540 14943 15598 14949
rect 15540 14940 15552 14943
rect 14415 14912 15552 14940
rect 14415 14909 14427 14912
rect 14369 14903 14427 14909
rect 15540 14909 15552 14912
rect 15586 14909 15598 14943
rect 15540 14903 15598 14909
rect 19496 14943 19554 14949
rect 19496 14909 19508 14943
rect 19542 14940 19554 14943
rect 20254 14940 20260 14952
rect 19542 14912 20260 14940
rect 19542 14909 19554 14912
rect 19496 14903 19554 14909
rect 20254 14900 20260 14912
rect 20312 14900 20318 14952
rect 8665 14875 8723 14881
rect 8665 14841 8677 14875
rect 8711 14872 8723 14875
rect 8846 14872 8852 14884
rect 8711 14844 8852 14872
rect 8711 14841 8723 14844
rect 8665 14835 8723 14841
rect 8846 14832 8852 14844
rect 8904 14832 8910 14884
rect 19981 14875 20039 14881
rect 19981 14841 19993 14875
rect 20027 14872 20039 14875
rect 20070 14872 20076 14884
rect 20027 14844 20076 14872
rect 20027 14841 20039 14844
rect 19981 14835 20039 14841
rect 20070 14832 20076 14844
rect 20128 14872 20134 14884
rect 20714 14872 20720 14884
rect 20128 14844 20720 14872
rect 20128 14832 20134 14844
rect 20714 14832 20720 14844
rect 20772 14832 20778 14884
rect 7374 14764 7380 14816
rect 7432 14804 7438 14816
rect 7745 14807 7803 14813
rect 7745 14804 7757 14807
rect 7432 14776 7757 14804
rect 7432 14764 7438 14776
rect 7745 14773 7757 14776
rect 7791 14773 7803 14807
rect 7745 14767 7803 14773
rect 15611 14807 15669 14813
rect 15611 14773 15623 14807
rect 15657 14804 15669 14807
rect 15838 14804 15844 14816
rect 15657 14776 15844 14804
rect 15657 14773 15669 14776
rect 15611 14767 15669 14773
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 1104 14714 21436 14736
rect 1104 14662 8497 14714
rect 8549 14662 8561 14714
rect 8613 14662 8625 14714
rect 8677 14662 8689 14714
rect 8741 14662 16012 14714
rect 16064 14662 16076 14714
rect 16128 14662 16140 14714
rect 16192 14662 16204 14714
rect 16256 14662 21436 14714
rect 1104 14640 21436 14662
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 9815 14603 9873 14609
rect 9815 14600 9827 14603
rect 8904 14572 9827 14600
rect 8904 14560 8910 14572
rect 9815 14569 9827 14572
rect 9861 14569 9873 14603
rect 9815 14563 9873 14569
rect 13446 14560 13452 14612
rect 13504 14600 13510 14612
rect 13817 14603 13875 14609
rect 13817 14600 13829 14603
rect 13504 14572 13829 14600
rect 13504 14560 13510 14572
rect 13817 14569 13829 14572
rect 13863 14569 13875 14603
rect 13817 14563 13875 14569
rect 15838 14492 15844 14544
rect 15896 14532 15902 14544
rect 16117 14535 16175 14541
rect 16117 14532 16129 14535
rect 15896 14504 16129 14532
rect 15896 14492 15902 14504
rect 16117 14501 16129 14504
rect 16163 14501 16175 14535
rect 16117 14495 16175 14501
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 9766 14464 9772 14476
rect 9631 14436 9772 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 13630 14464 13636 14476
rect 13591 14436 13636 14464
rect 13630 14424 13636 14436
rect 13688 14424 13694 14476
rect 16666 14328 16672 14340
rect 16627 14300 16672 14328
rect 16666 14288 16672 14300
rect 16724 14288 16730 14340
rect 1104 14170 21436 14192
rect 1104 14118 4739 14170
rect 4791 14118 4803 14170
rect 4855 14118 4867 14170
rect 4919 14118 4931 14170
rect 4983 14118 12255 14170
rect 12307 14118 12319 14170
rect 12371 14118 12383 14170
rect 12435 14118 12447 14170
rect 12499 14118 19770 14170
rect 19822 14118 19834 14170
rect 19886 14118 19898 14170
rect 19950 14118 19962 14170
rect 20014 14118 21436 14170
rect 1104 14096 21436 14118
rect 9766 14056 9772 14068
rect 9727 14028 9772 14056
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10505 14059 10563 14065
rect 10505 14025 10517 14059
rect 10551 14056 10563 14059
rect 10870 14056 10876 14068
rect 10551 14028 10876 14056
rect 10551 14025 10563 14028
rect 10505 14019 10563 14025
rect 10020 13855 10078 13861
rect 10020 13821 10032 13855
rect 10066 13852 10078 13855
rect 10520 13852 10548 14019
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 13630 14056 13636 14068
rect 13591 14028 13636 14056
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 15838 14016 15844 14068
rect 15896 14056 15902 14068
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 15896 14028 15945 14056
rect 15896 14016 15902 14028
rect 15933 14025 15945 14028
rect 15979 14025 15991 14059
rect 15933 14019 15991 14025
rect 18230 13948 18236 14000
rect 18288 13988 18294 14000
rect 20254 13988 20260 14000
rect 18288 13960 20260 13988
rect 18288 13948 18294 13960
rect 16666 13920 16672 13932
rect 16627 13892 16672 13920
rect 16666 13880 16672 13892
rect 16724 13920 16730 13932
rect 19061 13923 19119 13929
rect 19061 13920 19073 13923
rect 16724 13892 19073 13920
rect 16724 13880 16730 13892
rect 19061 13889 19073 13892
rect 19107 13920 19119 13923
rect 19150 13920 19156 13932
rect 19107 13892 19156 13920
rect 19107 13889 19119 13892
rect 19061 13883 19119 13889
rect 19150 13880 19156 13892
rect 19208 13880 19214 13932
rect 19628 13929 19656 13960
rect 20254 13948 20260 13960
rect 20312 13948 20318 14000
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 10066 13824 10548 13852
rect 10066 13821 10078 13824
rect 10020 13815 10078 13821
rect 16209 13787 16267 13793
rect 16209 13753 16221 13787
rect 16255 13784 16267 13787
rect 16298 13784 16304 13796
rect 16255 13756 16304 13784
rect 16255 13753 16267 13756
rect 16209 13747 16267 13753
rect 16298 13744 16304 13756
rect 16356 13744 16362 13796
rect 19150 13744 19156 13796
rect 19208 13784 19214 13796
rect 19337 13787 19395 13793
rect 19337 13784 19349 13787
rect 19208 13756 19349 13784
rect 19208 13744 19214 13756
rect 19337 13753 19349 13756
rect 19383 13784 19395 13787
rect 19426 13784 19432 13796
rect 19383 13756 19432 13784
rect 19383 13753 19395 13756
rect 19337 13747 19395 13753
rect 19426 13744 19432 13756
rect 19484 13744 19490 13796
rect 10042 13676 10048 13728
rect 10100 13716 10106 13728
rect 10229 13719 10287 13725
rect 10229 13716 10241 13719
rect 10100 13688 10241 13716
rect 10100 13676 10106 13688
rect 10229 13685 10241 13688
rect 10275 13685 10287 13719
rect 10229 13679 10287 13685
rect 1104 13626 21436 13648
rect 1104 13574 8497 13626
rect 8549 13574 8561 13626
rect 8613 13574 8625 13626
rect 8677 13574 8689 13626
rect 8741 13574 16012 13626
rect 16064 13574 16076 13626
rect 16128 13574 16140 13626
rect 16192 13574 16204 13626
rect 16256 13574 21436 13626
rect 1104 13552 21436 13574
rect 15795 13515 15853 13521
rect 15795 13481 15807 13515
rect 15841 13512 15853 13515
rect 16209 13515 16267 13521
rect 16209 13512 16221 13515
rect 15841 13484 16221 13512
rect 15841 13481 15853 13484
rect 15795 13475 15853 13481
rect 16209 13481 16221 13484
rect 16255 13512 16267 13515
rect 16298 13512 16304 13524
rect 16255 13484 16304 13512
rect 16255 13481 16267 13484
rect 16209 13475 16267 13481
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 13630 13336 13636 13388
rect 13688 13376 13694 13388
rect 15654 13376 15660 13388
rect 13688 13348 15660 13376
rect 13688 13336 13694 13348
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 10042 13308 10048 13320
rect 10003 13280 10048 13308
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 10410 13308 10416 13320
rect 10371 13280 10416 13308
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 1104 13082 21436 13104
rect 1104 13030 4739 13082
rect 4791 13030 4803 13082
rect 4855 13030 4867 13082
rect 4919 13030 4931 13082
rect 4983 13030 12255 13082
rect 12307 13030 12319 13082
rect 12371 13030 12383 13082
rect 12435 13030 12447 13082
rect 12499 13030 19770 13082
rect 19822 13030 19834 13082
rect 19886 13030 19898 13082
rect 19950 13030 19962 13082
rect 20014 13030 21436 13082
rect 1104 13008 21436 13030
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10781 12971 10839 12977
rect 10781 12968 10793 12971
rect 10100 12940 10793 12968
rect 10100 12928 10106 12940
rect 10781 12937 10793 12940
rect 10827 12937 10839 12971
rect 10781 12931 10839 12937
rect 10410 12900 10416 12912
rect 10371 12872 10416 12900
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 19705 12835 19763 12841
rect 19705 12832 19717 12835
rect 19484 12804 19717 12832
rect 19484 12792 19490 12804
rect 19705 12801 19717 12804
rect 19751 12801 19763 12835
rect 19705 12795 19763 12801
rect 9677 12699 9735 12705
rect 9677 12665 9689 12699
rect 9723 12696 9735 12699
rect 9858 12696 9864 12708
rect 9723 12668 9864 12696
rect 9723 12665 9735 12668
rect 9677 12659 9735 12665
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 19245 12699 19303 12705
rect 19245 12665 19257 12699
rect 19291 12696 19303 12699
rect 19426 12696 19432 12708
rect 19291 12668 19432 12696
rect 19291 12665 19303 12668
rect 19245 12659 19303 12665
rect 19426 12656 19432 12668
rect 19484 12656 19490 12708
rect 15654 12628 15660 12640
rect 15615 12600 15660 12628
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 1104 12538 21436 12560
rect 1104 12486 8497 12538
rect 8549 12486 8561 12538
rect 8613 12486 8625 12538
rect 8677 12486 8689 12538
rect 8741 12486 16012 12538
rect 16064 12486 16076 12538
rect 16128 12486 16140 12538
rect 16192 12486 16204 12538
rect 16256 12486 21436 12538
rect 1104 12464 21436 12486
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19751 12427 19809 12433
rect 19751 12424 19763 12427
rect 19484 12396 19763 12424
rect 19484 12384 19490 12396
rect 19751 12393 19763 12396
rect 19797 12393 19809 12427
rect 19751 12387 19809 12393
rect 9766 12356 9772 12368
rect 9679 12328 9772 12356
rect 9766 12316 9772 12328
rect 9824 12356 9830 12368
rect 10410 12356 10416 12368
rect 9824 12328 10416 12356
rect 9824 12316 9830 12328
rect 10410 12316 10416 12328
rect 10468 12316 10474 12368
rect 19610 12288 19616 12300
rect 19571 12260 19616 12288
rect 19610 12248 19616 12260
rect 19668 12248 19674 12300
rect 8478 12220 8484 12232
rect 8439 12192 8484 12220
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 10045 12223 10103 12229
rect 10045 12220 10057 12223
rect 9456 12192 10057 12220
rect 9456 12180 9462 12192
rect 10045 12189 10057 12192
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 1104 11994 21436 12016
rect 1104 11942 4739 11994
rect 4791 11942 4803 11994
rect 4855 11942 4867 11994
rect 4919 11942 4931 11994
rect 4983 11942 12255 11994
rect 12307 11942 12319 11994
rect 12371 11942 12383 11994
rect 12435 11942 12447 11994
rect 12499 11942 19770 11994
rect 19822 11942 19834 11994
rect 19886 11942 19898 11994
rect 19950 11942 19962 11994
rect 20014 11942 21436 11994
rect 1104 11920 21436 11942
rect 8478 11880 8484 11892
rect 8439 11852 8484 11880
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 9766 11880 9772 11892
rect 9727 11852 9772 11880
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 10367 11883 10425 11889
rect 10367 11880 10379 11883
rect 9916 11852 10379 11880
rect 9916 11840 9922 11852
rect 10367 11849 10379 11852
rect 10413 11849 10425 11883
rect 12618 11880 12624 11892
rect 12579 11852 12624 11880
rect 10367 11843 10425 11849
rect 12618 11840 12624 11852
rect 12676 11840 12682 11892
rect 8496 11744 8524 11840
rect 8757 11747 8815 11753
rect 8757 11744 8769 11747
rect 8496 11716 8769 11744
rect 8757 11713 8769 11716
rect 8803 11713 8815 11747
rect 9398 11744 9404 11756
rect 9359 11716 9404 11744
rect 8757 11707 8815 11713
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 16393 11747 16451 11753
rect 16393 11744 16405 11747
rect 15891 11716 16405 11744
rect 7720 11679 7778 11685
rect 7720 11645 7732 11679
rect 7766 11645 7778 11679
rect 7720 11639 7778 11645
rect 7735 11608 7763 11639
rect 8205 11611 8263 11617
rect 8205 11608 8217 11611
rect 7735 11580 8217 11608
rect 8205 11577 8217 11580
rect 8251 11608 8263 11611
rect 9416 11608 9444 11704
rect 10296 11679 10354 11685
rect 10296 11645 10308 11679
rect 10342 11676 10354 11679
rect 10686 11676 10692 11688
rect 10342 11648 10692 11676
rect 10342 11645 10354 11648
rect 10296 11639 10354 11645
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11676 12495 11679
rect 12618 11676 12624 11688
rect 12483 11648 12624 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 12618 11636 12624 11648
rect 12676 11676 12682 11688
rect 12989 11679 13047 11685
rect 12989 11676 13001 11679
rect 12676 11648 13001 11676
rect 12676 11636 12682 11648
rect 12989 11645 13001 11648
rect 13035 11645 13047 11679
rect 12989 11639 13047 11645
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15654 11676 15660 11688
rect 15344 11648 15660 11676
rect 15344 11636 15350 11648
rect 15654 11636 15660 11648
rect 15712 11676 15718 11688
rect 15891 11685 15919 11716
rect 16393 11713 16405 11716
rect 16439 11713 16451 11747
rect 16393 11707 16451 11713
rect 15876 11679 15934 11685
rect 15876 11676 15888 11679
rect 15712 11648 15888 11676
rect 15712 11636 15718 11648
rect 15876 11645 15888 11648
rect 15922 11645 15934 11679
rect 15876 11639 15934 11645
rect 15979 11679 16037 11685
rect 15979 11645 15991 11679
rect 16025 11676 16037 11679
rect 16298 11676 16304 11688
rect 16025 11648 16304 11676
rect 16025 11645 16037 11648
rect 15979 11639 16037 11645
rect 16298 11636 16304 11648
rect 16356 11636 16362 11688
rect 16888 11679 16946 11685
rect 16888 11645 16900 11679
rect 16934 11645 16946 11679
rect 19096 11679 19154 11685
rect 19096 11676 19108 11679
rect 16888 11639 16946 11645
rect 18892 11648 19108 11676
rect 8251 11580 9444 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 10870 11568 10876 11620
rect 10928 11608 10934 11620
rect 16903 11608 16931 11639
rect 17313 11611 17371 11617
rect 17313 11608 17325 11611
rect 10928 11580 17325 11608
rect 10928 11568 10934 11580
rect 17313 11577 17325 11580
rect 17359 11577 17371 11611
rect 17313 11571 17371 11577
rect 7791 11543 7849 11549
rect 7791 11509 7803 11543
rect 7837 11540 7849 11543
rect 7926 11540 7932 11552
rect 7837 11512 7932 11540
rect 7837 11509 7849 11512
rect 7791 11503 7849 11509
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 16991 11543 17049 11549
rect 16991 11540 17003 11543
rect 16448 11512 17003 11540
rect 16448 11500 16454 11512
rect 16991 11509 17003 11512
rect 17037 11509 17049 11543
rect 18046 11540 18052 11552
rect 18007 11512 18052 11540
rect 16991 11503 17049 11509
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18690 11500 18696 11552
rect 18748 11540 18754 11552
rect 18892 11549 18920 11648
rect 19096 11645 19108 11648
rect 19142 11645 19154 11679
rect 19096 11639 19154 11645
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 18748 11512 18889 11540
rect 18748 11500 18754 11512
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18877 11503 18935 11509
rect 19199 11543 19257 11549
rect 19199 11509 19211 11543
rect 19245 11540 19257 11543
rect 19518 11540 19524 11552
rect 19245 11512 19524 11540
rect 19245 11509 19257 11512
rect 19199 11503 19257 11509
rect 19518 11500 19524 11512
rect 19576 11500 19582 11552
rect 19610 11500 19616 11552
rect 19668 11540 19674 11552
rect 19705 11543 19763 11549
rect 19705 11540 19717 11543
rect 19668 11512 19717 11540
rect 19668 11500 19674 11512
rect 19705 11509 19717 11512
rect 19751 11540 19763 11543
rect 20622 11540 20628 11552
rect 19751 11512 20628 11540
rect 19751 11509 19763 11512
rect 19705 11503 19763 11509
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 1104 11450 21436 11472
rect 1104 11398 8497 11450
rect 8549 11398 8561 11450
rect 8613 11398 8625 11450
rect 8677 11398 8689 11450
rect 8741 11398 16012 11450
rect 16064 11398 16076 11450
rect 16128 11398 16140 11450
rect 16192 11398 16204 11450
rect 16256 11398 21436 11450
rect 1104 11376 21436 11398
rect 12618 11336 12624 11348
rect 12579 11308 12624 11336
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 19794 11336 19800 11348
rect 19755 11308 19800 11336
rect 19794 11296 19800 11308
rect 19852 11296 19858 11348
rect 16390 11268 16396 11280
rect 16351 11240 16396 11268
rect 16390 11228 16396 11240
rect 16448 11228 16454 11280
rect 7926 11200 7932 11212
rect 7887 11172 7932 11200
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 12504 11203 12562 11209
rect 12504 11169 12516 11203
rect 12550 11200 12562 11203
rect 12894 11200 12900 11212
rect 12550 11172 12900 11200
rect 12550 11169 12562 11172
rect 12504 11163 12562 11169
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 19518 11160 19524 11212
rect 19576 11200 19582 11212
rect 19613 11203 19671 11209
rect 19613 11200 19625 11203
rect 19576 11172 19625 11200
rect 19576 11160 19582 11172
rect 19613 11169 19625 11172
rect 19659 11169 19671 11203
rect 19613 11163 19671 11169
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 17957 11135 18015 11141
rect 17957 11132 17969 11135
rect 16960 11104 17969 11132
rect 16960 11076 16988 11104
rect 17957 11101 17969 11104
rect 18003 11101 18015 11135
rect 17957 11095 18015 11101
rect 18601 11135 18659 11141
rect 18601 11101 18613 11135
rect 18647 11132 18659 11135
rect 18782 11132 18788 11144
rect 18647 11104 18788 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 8110 11064 8116 11076
rect 8071 11036 8116 11064
rect 8110 11024 8116 11036
rect 8168 11024 8174 11076
rect 16942 11064 16948 11076
rect 16903 11036 16948 11064
rect 16942 11024 16948 11036
rect 17000 11024 17006 11076
rect 1104 10906 21436 10928
rect 1104 10854 4739 10906
rect 4791 10854 4803 10906
rect 4855 10854 4867 10906
rect 4919 10854 4931 10906
rect 4983 10854 12255 10906
rect 12307 10854 12319 10906
rect 12371 10854 12383 10906
rect 12435 10854 12447 10906
rect 12499 10854 19770 10906
rect 19822 10854 19834 10906
rect 19886 10854 19898 10906
rect 19950 10854 19962 10906
rect 20014 10854 21436 10906
rect 1104 10832 21436 10854
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 8389 10795 8447 10801
rect 8389 10792 8401 10795
rect 7984 10764 8401 10792
rect 7984 10752 7990 10764
rect 8389 10761 8401 10764
rect 8435 10761 8447 10795
rect 12894 10792 12900 10804
rect 12855 10764 12900 10792
rect 8389 10755 8447 10761
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 16298 10792 16304 10804
rect 16259 10764 16304 10792
rect 16298 10752 16304 10764
rect 16356 10792 16362 10804
rect 16356 10764 16528 10792
rect 16356 10752 16362 10764
rect 15933 10727 15991 10733
rect 15933 10693 15945 10727
rect 15979 10724 15991 10727
rect 16390 10724 16396 10736
rect 15979 10696 16396 10724
rect 15979 10693 15991 10696
rect 15933 10687 15991 10693
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 16500 10665 16528 10764
rect 18046 10752 18052 10804
rect 18104 10792 18110 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 18104 10764 18245 10792
rect 18104 10752 18110 10764
rect 18233 10761 18245 10764
rect 18279 10792 18291 10795
rect 18279 10764 18552 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7340 10628 7757 10656
rect 7340 10616 7346 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 16485 10659 16543 10665
rect 16485 10625 16497 10659
rect 16531 10625 16543 10659
rect 16942 10656 16948 10668
rect 16903 10628 16948 10656
rect 16485 10619 16543 10625
rect 16942 10616 16948 10628
rect 17000 10656 17006 10668
rect 18524 10665 18552 10764
rect 19518 10752 19524 10804
rect 19576 10792 19582 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 19576 10764 19625 10792
rect 19576 10752 19582 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 19613 10755 19671 10761
rect 20165 10727 20223 10733
rect 20165 10693 20177 10727
rect 20211 10724 20223 10727
rect 22094 10724 22100 10736
rect 20211 10696 22100 10724
rect 20211 10693 20223 10696
rect 20165 10687 20223 10693
rect 22094 10684 22100 10696
rect 22152 10684 22158 10736
rect 17773 10659 17831 10665
rect 17773 10656 17785 10659
rect 17000 10628 17785 10656
rect 17000 10616 17006 10628
rect 17773 10625 17785 10628
rect 17819 10625 17831 10659
rect 17773 10619 17831 10625
rect 18509 10659 18567 10665
rect 18509 10625 18521 10659
rect 18555 10625 18567 10659
rect 18782 10656 18788 10668
rect 18743 10628 18788 10656
rect 18509 10619 18567 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 106 10548 112 10600
rect 164 10588 170 10600
rect 1432 10591 1490 10597
rect 1432 10588 1444 10591
rect 164 10560 1444 10588
rect 164 10548 170 10560
rect 1432 10557 1444 10560
rect 1478 10588 1490 10591
rect 1857 10591 1915 10597
rect 1857 10588 1869 10591
rect 1478 10560 1869 10588
rect 1478 10557 1490 10560
rect 1432 10551 1490 10557
rect 1857 10557 1869 10560
rect 1903 10588 1915 10591
rect 2444 10591 2502 10597
rect 2444 10588 2456 10591
rect 1903 10560 2456 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2444 10557 2456 10560
rect 2490 10588 2502 10591
rect 2869 10591 2927 10597
rect 2869 10588 2881 10591
rect 2490 10560 2881 10588
rect 2490 10557 2502 10560
rect 2444 10551 2502 10557
rect 2869 10557 2881 10560
rect 2915 10557 2927 10591
rect 2869 10551 2927 10557
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 20070 10588 20076 10600
rect 20027 10560 20076 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 20070 10548 20076 10560
rect 20128 10588 20134 10600
rect 20533 10591 20591 10597
rect 20533 10588 20545 10591
rect 20128 10560 20545 10588
rect 20128 10548 20134 10560
rect 20533 10557 20545 10560
rect 20579 10557 20591 10591
rect 20533 10551 20591 10557
rect 1535 10523 1593 10529
rect 1535 10489 1547 10523
rect 1581 10520 1593 10523
rect 1946 10520 1952 10532
rect 1581 10492 1952 10520
rect 1581 10489 1593 10492
rect 1535 10483 1593 10489
rect 1946 10480 1952 10492
rect 2004 10480 2010 10532
rect 7285 10523 7343 10529
rect 7285 10489 7297 10523
rect 7331 10520 7343 10523
rect 7466 10520 7472 10532
rect 7331 10492 7472 10520
rect 7331 10489 7343 10492
rect 7285 10483 7343 10489
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 1854 10412 1860 10464
rect 1912 10452 1918 10464
rect 2547 10455 2605 10461
rect 2547 10452 2559 10455
rect 1912 10424 2559 10452
rect 1912 10412 1918 10424
rect 2547 10421 2559 10424
rect 2593 10421 2605 10455
rect 12434 10452 12440 10464
rect 12395 10424 12440 10452
rect 2547 10415 2605 10421
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 1104 10362 21436 10384
rect 1104 10310 8497 10362
rect 8549 10310 8561 10362
rect 8613 10310 8625 10362
rect 8677 10310 8689 10362
rect 8741 10310 16012 10362
rect 16064 10310 16076 10362
rect 16128 10310 16140 10362
rect 16192 10310 16204 10362
rect 16256 10310 21436 10362
rect 1104 10288 21436 10310
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 6178 10248 6184 10260
rect 5675 10220 6184 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 8251 10251 8309 10257
rect 8251 10248 8263 10251
rect 7524 10220 8263 10248
rect 7524 10208 7530 10220
rect 8251 10217 8263 10220
rect 8297 10217 8309 10251
rect 8251 10211 8309 10217
rect 7282 10180 7288 10192
rect 7243 10152 7288 10180
rect 7282 10140 7288 10152
rect 7340 10140 7346 10192
rect 12434 10140 12440 10192
rect 12492 10180 12498 10192
rect 12802 10180 12808 10192
rect 12492 10152 12808 10180
rect 12492 10140 12498 10152
rect 12802 10140 12808 10152
rect 12860 10140 12866 10192
rect 5442 10112 5448 10124
rect 5403 10084 5448 10112
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 8110 10112 8116 10124
rect 8071 10084 8116 10112
rect 8110 10072 8116 10084
rect 8168 10112 8174 10124
rect 10870 10112 10876 10124
rect 8168 10084 10876 10112
rect 8168 10072 8174 10084
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 1946 10044 1952 10056
rect 1627 10016 1952 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 6638 10044 6644 10056
rect 6599 10016 6644 10044
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 12894 10004 12900 10056
rect 12952 10044 12958 10056
rect 13081 10047 13139 10053
rect 13081 10044 13093 10047
rect 12952 10016 13093 10044
rect 12952 10004 12958 10016
rect 13081 10013 13093 10016
rect 13127 10013 13139 10047
rect 13081 10007 13139 10013
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10044 17371 10047
rect 18414 10044 18420 10056
rect 17359 10016 18420 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 18414 10004 18420 10016
rect 18472 10004 18478 10056
rect 18690 10044 18696 10056
rect 18651 10016 18696 10044
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 2130 9976 2136 9988
rect 2091 9948 2136 9976
rect 2130 9936 2136 9948
rect 2188 9936 2194 9988
rect 1104 9818 21436 9840
rect 1104 9766 4739 9818
rect 4791 9766 4803 9818
rect 4855 9766 4867 9818
rect 4919 9766 4931 9818
rect 4983 9766 12255 9818
rect 12307 9766 12319 9818
rect 12371 9766 12383 9818
rect 12435 9766 12447 9818
rect 12499 9766 19770 9818
rect 19822 9766 19834 9818
rect 19886 9766 19898 9818
rect 19950 9766 19962 9818
rect 20014 9766 21436 9818
rect 1104 9744 21436 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 2869 9707 2927 9713
rect 2869 9704 2881 9707
rect 1452 9676 2881 9704
rect 1452 9664 1458 9676
rect 2869 9673 2881 9676
rect 2915 9704 2927 9707
rect 3142 9704 3148 9716
rect 2915 9676 3148 9704
rect 2915 9673 2927 9676
rect 2869 9667 2927 9673
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 5859 9707 5917 9713
rect 5859 9673 5871 9707
rect 5905 9704 5917 9707
rect 6638 9704 6644 9716
rect 5905 9676 6644 9704
rect 5905 9673 5917 9676
rect 5859 9667 5917 9673
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 8110 9704 8116 9716
rect 8071 9676 8116 9704
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 12802 9704 12808 9716
rect 12763 9676 12808 9704
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 18414 9664 18420 9716
rect 18472 9704 18478 9716
rect 19061 9707 19119 9713
rect 19061 9704 19073 9707
rect 18472 9676 19073 9704
rect 18472 9664 18478 9676
rect 19061 9673 19073 9676
rect 19107 9673 19119 9707
rect 19061 9667 19119 9673
rect 19150 9664 19156 9716
rect 19208 9704 19214 9716
rect 19797 9707 19855 9713
rect 19797 9704 19809 9707
rect 19208 9676 19809 9704
rect 19208 9664 19214 9676
rect 19797 9673 19809 9676
rect 19843 9673 19855 9707
rect 19797 9667 19855 9673
rect 2130 9636 2136 9648
rect 2091 9608 2136 9636
rect 2130 9596 2136 9608
rect 2188 9636 2194 9648
rect 2188 9608 3464 9636
rect 2188 9596 2194 9608
rect 3142 9568 3148 9580
rect 3103 9540 3148 9568
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3436 9577 3464 9608
rect 5442 9596 5448 9648
rect 5500 9636 5506 9648
rect 5537 9639 5595 9645
rect 5537 9636 5549 9639
rect 5500 9608 5549 9636
rect 5500 9596 5506 9608
rect 5537 9605 5549 9608
rect 5583 9636 5595 9639
rect 8711 9639 8769 9645
rect 8711 9636 8723 9639
rect 5583 9608 8723 9636
rect 5583 9605 5595 9608
rect 5537 9599 5595 9605
rect 8711 9605 8723 9608
rect 8757 9605 8769 9639
rect 18690 9636 18696 9648
rect 18651 9608 18696 9636
rect 8711 9599 8769 9605
rect 18690 9596 18696 9608
rect 18748 9596 18754 9648
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9568 7159 9571
rect 7282 9568 7288 9580
rect 7147 9540 7288 9568
rect 7147 9537 7159 9540
rect 7101 9531 7159 9537
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 8220 9540 9536 9568
rect 5788 9503 5846 9509
rect 5788 9469 5800 9503
rect 5834 9500 5846 9503
rect 5834 9472 6316 9500
rect 5834 9469 5846 9472
rect 5788 9463 5846 9469
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 1670 9432 1676 9444
rect 1627 9404 1676 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 1670 9392 1676 9404
rect 1728 9392 1734 9444
rect 6288 9373 6316 9472
rect 7745 9435 7803 9441
rect 7745 9401 7757 9435
rect 7791 9432 7803 9435
rect 7926 9432 7932 9444
rect 7791 9404 7932 9432
rect 7791 9401 7803 9404
rect 7745 9395 7803 9401
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 8220 9432 8248 9540
rect 9508 9512 9536 9540
rect 12894 9528 12900 9580
rect 12952 9568 12958 9580
rect 13633 9571 13691 9577
rect 13633 9568 13645 9571
rect 12952 9540 13645 9568
rect 12952 9528 12958 9540
rect 13633 9537 13645 9540
rect 13679 9537 13691 9571
rect 13633 9531 13691 9537
rect 16868 9540 19656 9568
rect 8640 9503 8698 9509
rect 8640 9469 8652 9503
rect 8686 9500 8698 9503
rect 8686 9472 9076 9500
rect 8686 9469 8698 9472
rect 8640 9463 8698 9469
rect 8036 9404 8248 9432
rect 6273 9367 6331 9373
rect 6273 9333 6285 9367
rect 6319 9364 6331 9367
rect 8036 9364 8064 9404
rect 9048 9376 9076 9472
rect 9490 9460 9496 9512
rect 9548 9500 9554 9512
rect 9620 9503 9678 9509
rect 9620 9500 9632 9503
rect 9548 9472 9632 9500
rect 9548 9460 9554 9472
rect 9620 9469 9632 9472
rect 9666 9500 9678 9503
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9666 9472 10057 9500
rect 9666 9469 9678 9472
rect 9620 9463 9678 9469
rect 10045 9469 10057 9472
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 14550 9460 14556 9512
rect 14608 9500 14614 9512
rect 16868 9509 16896 9540
rect 19628 9509 19656 9540
rect 16428 9503 16486 9509
rect 16428 9500 16440 9503
rect 14608 9472 16440 9500
rect 14608 9460 14614 9472
rect 16428 9469 16440 9472
rect 16474 9500 16486 9503
rect 16853 9503 16911 9509
rect 16853 9500 16865 9503
rect 16474 9472 16865 9500
rect 16474 9469 16486 9472
rect 16428 9463 16486 9469
rect 16853 9469 16865 9472
rect 16899 9469 16911 9503
rect 16853 9463 16911 9469
rect 19613 9503 19671 9509
rect 19613 9469 19625 9503
rect 19659 9500 19671 9503
rect 20165 9503 20223 9509
rect 20165 9500 20177 9503
rect 19659 9472 20177 9500
rect 19659 9469 19671 9472
rect 19613 9463 19671 9469
rect 20165 9469 20177 9472
rect 20211 9469 20223 9503
rect 20165 9463 20223 9469
rect 13173 9435 13231 9441
rect 13173 9401 13185 9435
rect 13219 9432 13231 9435
rect 13357 9435 13415 9441
rect 13357 9432 13369 9435
rect 13219 9404 13369 9432
rect 13219 9401 13231 9404
rect 13173 9395 13231 9401
rect 13357 9401 13369 9404
rect 13403 9432 13415 9435
rect 14090 9432 14096 9444
rect 13403 9404 14096 9432
rect 13403 9401 13415 9404
rect 13357 9395 13415 9401
rect 14090 9392 14096 9404
rect 14148 9392 14154 9444
rect 18141 9435 18199 9441
rect 18141 9432 18153 9435
rect 17788 9404 18153 9432
rect 9030 9364 9036 9376
rect 6319 9336 8064 9364
rect 8991 9336 9036 9364
rect 6319 9333 6331 9336
rect 6273 9327 6331 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 9723 9367 9781 9373
rect 9723 9364 9735 9367
rect 9180 9336 9735 9364
rect 9180 9324 9186 9336
rect 9723 9333 9735 9336
rect 9769 9333 9781 9367
rect 9723 9327 9781 9333
rect 16531 9367 16589 9373
rect 16531 9333 16543 9367
rect 16577 9364 16589 9367
rect 16666 9364 16672 9376
rect 16577 9336 16672 9364
rect 16577 9333 16589 9336
rect 16531 9327 16589 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 17126 9324 17132 9376
rect 17184 9364 17190 9376
rect 17788 9373 17816 9404
rect 18141 9401 18153 9404
rect 18187 9401 18199 9435
rect 18141 9395 18199 9401
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17184 9336 17785 9364
rect 17184 9324 17190 9336
rect 17773 9333 17785 9336
rect 17819 9333 17831 9367
rect 17773 9327 17831 9333
rect 1104 9274 21436 9296
rect 1104 9222 8497 9274
rect 8549 9222 8561 9274
rect 8613 9222 8625 9274
rect 8677 9222 8689 9274
rect 8741 9222 16012 9274
rect 16064 9222 16076 9274
rect 16128 9222 16140 9274
rect 16192 9222 16204 9274
rect 16256 9222 21436 9274
rect 1104 9200 21436 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 7101 9163 7159 9169
rect 7101 9160 7113 9163
rect 2188 9132 2268 9160
rect 2188 9120 2194 9132
rect 2240 9101 2268 9132
rect 6472 9132 7113 9160
rect 6472 9101 6500 9132
rect 7101 9129 7113 9132
rect 7147 9160 7159 9163
rect 7282 9160 7288 9172
rect 7147 9132 7288 9160
rect 7147 9129 7159 9132
rect 7101 9123 7159 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 19751 9163 19809 9169
rect 19751 9129 19763 9163
rect 19797 9160 19809 9163
rect 20070 9160 20076 9172
rect 19797 9132 20076 9160
rect 19797 9129 19809 9132
rect 19751 9123 19809 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 2225 9095 2283 9101
rect 2225 9061 2237 9095
rect 2271 9061 2283 9095
rect 2225 9055 2283 9061
rect 6457 9095 6515 9101
rect 6457 9061 6469 9095
rect 6503 9061 6515 9095
rect 6457 9055 6515 9061
rect 7377 9095 7435 9101
rect 7377 9061 7389 9095
rect 7423 9092 7435 9095
rect 7466 9092 7472 9104
rect 7423 9064 7472 9092
rect 7423 9061 7435 9064
rect 7377 9055 7435 9061
rect 7466 9052 7472 9064
rect 7524 9092 7530 9104
rect 9122 9092 9128 9104
rect 7524 9064 9128 9092
rect 7524 9052 7530 9064
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 16577 9095 16635 9101
rect 16577 9061 16589 9095
rect 16623 9092 16635 9095
rect 16666 9092 16672 9104
rect 16623 9064 16672 9092
rect 16623 9061 16635 9064
rect 16577 9055 16635 9061
rect 16666 9052 16672 9064
rect 16724 9052 16730 9104
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 4100 9027 4158 9033
rect 4100 9024 4112 9027
rect 4028 8996 4112 9024
rect 4028 8984 4034 8996
rect 4100 8993 4112 8996
rect 4146 8993 4158 9027
rect 4100 8987 4158 8993
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 9712 9027 9770 9033
rect 9712 9024 9724 9027
rect 9548 8996 9724 9024
rect 9548 8984 9554 8996
rect 9712 8993 9724 8996
rect 9758 8993 9770 9027
rect 9712 8987 9770 8993
rect 12066 8984 12072 9036
rect 12124 9024 12130 9036
rect 12380 9027 12438 9033
rect 12380 9024 12392 9027
rect 12124 8996 12392 9024
rect 12124 8984 12130 8996
rect 12380 8993 12392 8996
rect 12426 8993 12438 9027
rect 12380 8987 12438 8993
rect 18782 8984 18788 9036
rect 18840 9024 18846 9036
rect 19426 9024 19432 9036
rect 18840 8996 19432 9024
rect 18840 8984 18846 8996
rect 19426 8984 19432 8996
rect 19484 9024 19490 9036
rect 19648 9027 19706 9033
rect 19648 9024 19660 9027
rect 19484 8996 19660 9024
rect 19484 8984 19490 8996
rect 19648 8993 19660 8996
rect 19694 8993 19706 9027
rect 19648 8987 19706 8993
rect 2682 8956 2688 8968
rect 2643 8928 2688 8956
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 5813 8959 5871 8965
rect 5813 8925 5825 8959
rect 5859 8925 5871 8959
rect 7742 8956 7748 8968
rect 7703 8928 7748 8956
rect 5813 8919 5871 8925
rect 5718 8848 5724 8900
rect 5776 8888 5782 8900
rect 5828 8888 5856 8919
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 12483 8959 12541 8965
rect 12483 8925 12495 8959
rect 12529 8956 12541 8959
rect 13446 8956 13452 8968
rect 12529 8928 13452 8956
rect 12529 8925 12541 8928
rect 12483 8919 12541 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 14090 8956 14096 8968
rect 14051 8928 14096 8956
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 18138 8956 18144 8968
rect 18099 8928 18144 8956
rect 18138 8916 18144 8928
rect 18196 8916 18202 8968
rect 5776 8860 5856 8888
rect 5776 8848 5782 8860
rect 7926 8848 7932 8900
rect 7984 8888 7990 8900
rect 11698 8888 11704 8900
rect 7984 8860 11704 8888
rect 7984 8848 7990 8860
rect 11698 8848 11704 8860
rect 11756 8888 11762 8900
rect 17126 8888 17132 8900
rect 11756 8860 13814 8888
rect 17087 8860 17132 8888
rect 11756 8848 11762 8860
rect 1670 8820 1676 8832
rect 1631 8792 1676 8820
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 4203 8823 4261 8829
rect 4203 8820 4215 8823
rect 2280 8792 4215 8820
rect 2280 8780 2286 8792
rect 4203 8789 4215 8792
rect 4249 8789 4261 8823
rect 4203 8783 4261 8789
rect 9398 8780 9404 8832
rect 9456 8820 9462 8832
rect 9815 8823 9873 8829
rect 9815 8820 9827 8823
rect 9456 8792 9827 8820
rect 9456 8780 9462 8792
rect 9815 8789 9827 8792
rect 9861 8789 9873 8823
rect 13786 8820 13814 8860
rect 17126 8848 17132 8860
rect 17184 8848 17190 8900
rect 18693 8891 18751 8897
rect 18693 8888 18705 8891
rect 17696 8860 18705 8888
rect 17696 8820 17724 8860
rect 18693 8857 18705 8860
rect 18739 8857 18751 8891
rect 18693 8851 18751 8857
rect 13786 8792 17724 8820
rect 9815 8783 9873 8789
rect 1104 8730 21436 8752
rect 1104 8678 4739 8730
rect 4791 8678 4803 8730
rect 4855 8678 4867 8730
rect 4919 8678 4931 8730
rect 4983 8678 12255 8730
rect 12307 8678 12319 8730
rect 12371 8678 12383 8730
rect 12435 8678 12447 8730
rect 12499 8678 19770 8730
rect 19822 8678 19834 8730
rect 19886 8678 19898 8730
rect 19950 8678 19962 8730
rect 20014 8678 21436 8730
rect 1104 8656 21436 8678
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 2777 8619 2835 8625
rect 2777 8616 2789 8619
rect 2188 8588 2789 8616
rect 2188 8576 2194 8588
rect 2777 8585 2789 8588
rect 2823 8585 2835 8619
rect 2777 8579 2835 8585
rect 7377 8619 7435 8625
rect 7377 8585 7389 8619
rect 7423 8616 7435 8619
rect 7466 8616 7472 8628
rect 7423 8588 7472 8616
rect 7423 8585 7435 8588
rect 7377 8579 7435 8585
rect 7466 8576 7472 8588
rect 7524 8576 7530 8628
rect 9490 8616 9496 8628
rect 9451 8588 9496 8616
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 12066 8576 12072 8628
rect 12124 8616 12130 8628
rect 12618 8616 12624 8628
rect 12124 8588 12624 8616
rect 12124 8576 12130 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16666 8616 16672 8628
rect 16347 8588 16672 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 19426 8616 19432 8628
rect 19387 8588 19432 8616
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 1854 8480 1860 8492
rect 1719 8452 1860 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 2682 8440 2688 8492
rect 2740 8480 2746 8492
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 2740 8452 4537 8480
rect 2740 8440 2746 8452
rect 4525 8449 4537 8452
rect 4571 8449 4583 8483
rect 7742 8480 7748 8492
rect 7703 8452 7748 8480
rect 4525 8443 4583 8449
rect 7742 8440 7748 8452
rect 7800 8480 7806 8492
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 7800 8452 8677 8480
rect 7800 8440 7806 8452
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 9950 8480 9956 8492
rect 9911 8452 9956 8480
rect 8665 8443 8723 8449
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 14090 8440 14096 8492
rect 14148 8480 14154 8492
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 14148 8452 14381 8480
rect 14148 8440 14154 8452
rect 14369 8449 14381 8452
rect 14415 8449 14427 8483
rect 17126 8480 17132 8492
rect 17087 8452 17132 8480
rect 14369 8443 14427 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8480 17555 8483
rect 18138 8480 18144 8492
rect 17543 8452 18144 8480
rect 17543 8449 17555 8452
rect 17497 8443 17555 8449
rect 18138 8440 18144 8452
rect 18196 8480 18202 8492
rect 18417 8483 18475 8489
rect 18417 8480 18429 8483
rect 18196 8452 18429 8480
rect 18196 8440 18202 8452
rect 18417 8449 18429 8452
rect 18463 8480 18475 8483
rect 19150 8480 19156 8492
rect 18463 8452 19156 8480
rect 18463 8449 18475 8452
rect 18417 8443 18475 8449
rect 19150 8440 19156 8452
rect 19208 8480 19214 8492
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19208 8452 19993 8480
rect 19208 8440 19214 8452
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 2498 8344 2504 8356
rect 2459 8316 2504 8344
rect 2498 8304 2504 8316
rect 2556 8304 2562 8356
rect 3697 8347 3755 8353
rect 3697 8313 3709 8347
rect 3743 8344 3755 8347
rect 4249 8347 4307 8353
rect 4249 8344 4261 8347
rect 3743 8316 4261 8344
rect 3743 8313 3755 8316
rect 3697 8307 3755 8313
rect 4249 8313 4261 8316
rect 4295 8344 4307 8347
rect 5442 8344 5448 8356
rect 4295 8316 5448 8344
rect 4295 8313 4307 8316
rect 4249 8307 4307 8313
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 8389 8347 8447 8353
rect 8389 8313 8401 8347
rect 8435 8313 8447 8347
rect 8389 8307 8447 8313
rect 9125 8347 9183 8353
rect 9125 8313 9137 8347
rect 9171 8344 9183 8347
rect 9674 8344 9680 8356
rect 9171 8316 9680 8344
rect 9171 8313 9183 8316
rect 9125 8307 9183 8313
rect 1854 8236 1860 8288
rect 1912 8276 1918 8288
rect 3970 8276 3976 8288
rect 1912 8248 3976 8276
rect 1912 8236 1918 8248
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 5718 8276 5724 8288
rect 5679 8248 5724 8276
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 8404 8276 8432 8307
rect 9674 8304 9680 8316
rect 9732 8304 9738 8356
rect 13909 8347 13967 8353
rect 13909 8313 13921 8347
rect 13955 8344 13967 8347
rect 14090 8344 14096 8356
rect 13955 8316 14096 8344
rect 13955 8313 13967 8316
rect 13909 8307 13967 8313
rect 14090 8304 14096 8316
rect 14148 8304 14154 8356
rect 16485 8347 16543 8353
rect 16485 8313 16497 8347
rect 16531 8313 16543 8347
rect 18141 8347 18199 8353
rect 18141 8344 18153 8347
rect 16485 8307 16543 8313
rect 17788 8316 18153 8344
rect 9030 8276 9036 8288
rect 8404 8248 9036 8276
rect 9030 8236 9036 8248
rect 9088 8276 9094 8288
rect 10042 8276 10048 8288
rect 9088 8248 10048 8276
rect 9088 8236 9094 8248
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 16390 8236 16396 8288
rect 16448 8276 16454 8288
rect 16500 8276 16528 8307
rect 17788 8288 17816 8316
rect 18141 8313 18153 8316
rect 18187 8313 18199 8347
rect 19705 8347 19763 8353
rect 19705 8344 19717 8347
rect 18141 8307 18199 8313
rect 19076 8316 19717 8344
rect 19076 8288 19104 8316
rect 19705 8313 19717 8316
rect 19751 8313 19763 8347
rect 19705 8307 19763 8313
rect 17770 8276 17776 8288
rect 16448 8248 16528 8276
rect 17731 8248 17776 8276
rect 16448 8236 16454 8248
rect 17770 8236 17776 8248
rect 17828 8236 17834 8288
rect 19058 8276 19064 8288
rect 19019 8248 19064 8276
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 1104 8186 21436 8208
rect 1104 8134 8497 8186
rect 8549 8134 8561 8186
rect 8613 8134 8625 8186
rect 8677 8134 8689 8186
rect 8741 8134 16012 8186
rect 16064 8134 16076 8186
rect 16128 8134 16140 8186
rect 16192 8134 16204 8186
rect 16256 8134 21436 8186
rect 1104 8112 21436 8134
rect 4847 8075 4905 8081
rect 4847 8041 4859 8075
rect 4893 8072 4905 8075
rect 5718 8072 5724 8084
rect 4893 8044 5724 8072
rect 4893 8041 4905 8044
rect 4847 8035 4905 8041
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 11379 8075 11437 8081
rect 11379 8072 11391 8075
rect 9732 8044 11391 8072
rect 9732 8032 9738 8044
rect 11379 8041 11391 8044
rect 11425 8041 11437 8075
rect 11379 8035 11437 8041
rect 14090 8032 14096 8084
rect 14148 8072 14154 8084
rect 15427 8075 15485 8081
rect 15427 8072 15439 8075
rect 14148 8044 15439 8072
rect 14148 8032 14154 8044
rect 15427 8041 15439 8044
rect 15473 8041 15485 8075
rect 15427 8035 15485 8041
rect 16761 8075 16819 8081
rect 16761 8041 16773 8075
rect 16807 8072 16819 8075
rect 17770 8072 17776 8084
rect 16807 8044 17776 8072
rect 16807 8041 16819 8044
rect 16761 8035 16819 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 1857 8007 1915 8013
rect 1857 7973 1869 8007
rect 1903 8004 1915 8007
rect 1946 8004 1952 8016
rect 1903 7976 1952 8004
rect 1903 7973 1915 7976
rect 1857 7967 1915 7973
rect 1946 7964 1952 7976
rect 2004 8004 2010 8016
rect 2222 8004 2228 8016
rect 2004 7976 2228 8004
rect 2004 7964 2010 7976
rect 2222 7964 2228 7976
rect 2280 7964 2286 8016
rect 2498 8004 2504 8016
rect 2459 7976 2504 8004
rect 2498 7964 2504 7976
rect 2556 7964 2562 8016
rect 4614 7936 4620 7948
rect 4575 7908 4620 7936
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 10686 7896 10692 7948
rect 10744 7936 10750 7948
rect 11276 7939 11334 7945
rect 11276 7936 11288 7939
rect 10744 7908 11288 7936
rect 10744 7896 10750 7908
rect 11276 7905 11288 7908
rect 11322 7936 11334 7939
rect 11698 7936 11704 7948
rect 11322 7908 11704 7936
rect 11322 7905 11334 7908
rect 11276 7899 11334 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 12748 7939 12806 7945
rect 12748 7936 12760 7939
rect 12676 7908 12760 7936
rect 12676 7896 12682 7908
rect 12748 7905 12760 7908
rect 12794 7905 12806 7939
rect 12748 7899 12806 7905
rect 15356 7939 15414 7945
rect 15356 7905 15368 7939
rect 15402 7936 15414 7939
rect 15562 7936 15568 7948
rect 15402 7908 15568 7936
rect 15402 7905 15414 7908
rect 15356 7899 15414 7905
rect 15562 7896 15568 7908
rect 15620 7896 15626 7948
rect 17773 7939 17831 7945
rect 17773 7905 17785 7939
rect 17819 7936 17831 7939
rect 17862 7936 17868 7948
rect 17819 7908 17868 7936
rect 17819 7905 17831 7908
rect 17773 7899 17831 7905
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 7650 7868 7656 7880
rect 7611 7840 7656 7868
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7800 7840 7941 7868
rect 7800 7828 7806 7840
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 9766 7868 9772 7880
rect 8444 7840 9772 7868
rect 8444 7828 8450 7840
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 10042 7868 10048 7880
rect 10003 7840 10048 7868
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 18874 7868 18880 7880
rect 18835 7840 18880 7868
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 19150 7868 19156 7880
rect 19111 7840 19156 7868
rect 19150 7828 19156 7840
rect 19208 7828 19214 7880
rect 12851 7735 12909 7741
rect 12851 7701 12863 7735
rect 12897 7732 12909 7735
rect 12986 7732 12992 7744
rect 12897 7704 12992 7732
rect 12897 7701 12909 7704
rect 12851 7695 12909 7701
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 16390 7732 16396 7744
rect 16351 7704 16396 7732
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 17911 7735 17969 7741
rect 17911 7701 17923 7735
rect 17957 7732 17969 7735
rect 19242 7732 19248 7744
rect 17957 7704 19248 7732
rect 17957 7701 17969 7704
rect 17911 7695 17969 7701
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 1104 7642 21436 7664
rect 1104 7590 4739 7642
rect 4791 7590 4803 7642
rect 4855 7590 4867 7642
rect 4919 7590 4931 7642
rect 4983 7590 12255 7642
rect 12307 7590 12319 7642
rect 12371 7590 12383 7642
rect 12435 7590 12447 7642
rect 12499 7590 19770 7642
rect 19822 7590 19834 7642
rect 19886 7590 19898 7642
rect 19950 7590 19962 7642
rect 20014 7590 21436 7642
rect 1104 7568 21436 7590
rect 1535 7531 1593 7537
rect 1535 7497 1547 7531
rect 1581 7528 1593 7531
rect 1670 7528 1676 7540
rect 1581 7500 1676 7528
rect 1581 7497 1593 7500
rect 1535 7491 1593 7497
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 4614 7528 4620 7540
rect 4575 7500 4620 7528
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 9824 7500 10333 7528
rect 9824 7488 9830 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 11698 7528 11704 7540
rect 11659 7500 11704 7528
rect 10321 7491 10379 7497
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 12713 7531 12771 7537
rect 12713 7528 12725 7531
rect 12676 7500 12725 7528
rect 12676 7488 12682 7500
rect 12713 7497 12725 7500
rect 12759 7497 12771 7531
rect 16482 7528 16488 7540
rect 16443 7500 16488 7528
rect 12713 7491 12771 7497
rect 16482 7488 16488 7500
rect 16540 7488 16546 7540
rect 17862 7528 17868 7540
rect 17775 7500 17868 7528
rect 17862 7488 17868 7500
rect 17920 7528 17926 7540
rect 18690 7528 18696 7540
rect 17920 7500 18696 7528
rect 17920 7488 17926 7500
rect 8386 7460 8392 7472
rect 8347 7432 8392 7460
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 9950 7460 9956 7472
rect 8496 7432 9956 7460
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2556 7364 2789 7392
rect 2556 7352 2562 7364
rect 2777 7361 2789 7364
rect 2823 7392 2835 7395
rect 4154 7392 4160 7404
rect 2823 7364 4160 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 4338 7392 4344 7404
rect 4295 7364 4344 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 4338 7352 4344 7364
rect 4396 7392 4402 7404
rect 4801 7395 4859 7401
rect 4801 7392 4813 7395
rect 4396 7364 4813 7392
rect 4396 7352 4402 7364
rect 4801 7361 4813 7364
rect 4847 7361 4859 7395
rect 5442 7392 5448 7404
rect 5355 7364 5448 7392
rect 4801 7355 4859 7361
rect 5442 7352 5448 7364
rect 5500 7392 5506 7404
rect 8496 7392 8524 7432
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 11716 7460 11744 7488
rect 16117 7463 16175 7469
rect 11716 7432 13814 7460
rect 5500 7364 8524 7392
rect 9217 7395 9275 7401
rect 5500 7352 5506 7364
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 9398 7392 9404 7404
rect 9263 7364 9404 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7392 12311 7395
rect 12986 7392 12992 7404
rect 12299 7364 12992 7392
rect 12299 7361 12311 7364
rect 12253 7355 12311 7361
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 1464 7327 1522 7333
rect 1464 7293 1476 7327
rect 1510 7324 1522 7327
rect 1854 7324 1860 7336
rect 1510 7296 1860 7324
rect 1510 7293 1522 7296
rect 1464 7287 1522 7293
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 10908 7327 10966 7333
rect 10908 7293 10920 7327
rect 10954 7324 10966 7327
rect 11333 7327 11391 7333
rect 11333 7324 11345 7327
rect 10954 7296 11345 7324
rect 10954 7293 10966 7296
rect 10908 7287 10966 7293
rect 11333 7293 11345 7296
rect 11379 7293 11391 7327
rect 13786 7324 13814 7432
rect 16117 7429 16129 7463
rect 16163 7460 16175 7463
rect 16574 7460 16580 7472
rect 16163 7432 16580 7460
rect 16163 7429 16175 7432
rect 16117 7423 16175 7429
rect 16574 7420 16580 7432
rect 16632 7420 16638 7472
rect 15933 7327 15991 7333
rect 15933 7324 15945 7327
rect 13786 7296 15945 7324
rect 11333 7287 11391 7293
rect 15933 7293 15945 7296
rect 15979 7324 15991 7327
rect 16482 7324 16488 7336
rect 15979 7296 16488 7324
rect 15979 7293 15991 7296
rect 15933 7287 15991 7293
rect 2501 7259 2559 7265
rect 2501 7225 2513 7259
rect 2547 7225 2559 7259
rect 4614 7256 4620 7268
rect 2501 7219 2559 7225
rect 4126 7228 4620 7256
rect 2222 7188 2228 7200
rect 2183 7160 2228 7188
rect 2222 7148 2228 7160
rect 2280 7188 2286 7200
rect 2516 7188 2544 7219
rect 2280 7160 2544 7188
rect 2280 7148 2286 7160
rect 2590 7148 2596 7200
rect 2648 7188 2654 7200
rect 4126 7188 4154 7228
rect 4614 7216 4620 7228
rect 4672 7216 4678 7268
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 7653 7259 7711 7265
rect 7653 7256 7665 7259
rect 7616 7228 7665 7256
rect 7616 7216 7622 7228
rect 7653 7225 7665 7228
rect 7699 7256 7711 7259
rect 7837 7259 7895 7265
rect 7837 7256 7849 7259
rect 7699 7228 7849 7256
rect 7699 7225 7711 7228
rect 7653 7219 7711 7225
rect 7837 7225 7849 7228
rect 7883 7225 7895 7259
rect 7837 7219 7895 7225
rect 7926 7216 7932 7268
rect 7984 7256 7990 7268
rect 10923 7256 10951 7287
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 18191 7333 18219 7500
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 18322 7352 18328 7404
rect 18380 7392 18386 7404
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 18380 7364 19533 7392
rect 18380 7352 18386 7364
rect 19521 7361 19533 7364
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 18176 7327 18234 7333
rect 18176 7293 18188 7327
rect 18222 7293 18234 7327
rect 18176 7287 18234 7293
rect 13630 7256 13636 7268
rect 7984 7228 10951 7256
rect 13591 7228 13636 7256
rect 7984 7216 7990 7228
rect 13630 7216 13636 7228
rect 13688 7216 13694 7268
rect 18279 7259 18337 7265
rect 18279 7225 18291 7259
rect 18325 7256 18337 7259
rect 18874 7256 18880 7268
rect 18325 7228 18880 7256
rect 18325 7225 18337 7228
rect 18279 7219 18337 7225
rect 18874 7216 18880 7228
rect 18932 7216 18938 7268
rect 19245 7259 19303 7265
rect 19245 7225 19257 7259
rect 19291 7225 19303 7259
rect 19245 7219 19303 7225
rect 2648 7160 4154 7188
rect 7285 7191 7343 7197
rect 2648 7148 2654 7160
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 7742 7188 7748 7200
rect 7331 7160 7748 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 11011 7191 11069 7197
rect 11011 7157 11023 7191
rect 11057 7188 11069 7191
rect 11146 7188 11152 7200
rect 11057 7160 11152 7188
rect 11057 7157 11069 7160
rect 11011 7151 11069 7157
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 15381 7191 15439 7197
rect 15381 7157 15393 7191
rect 15427 7188 15439 7191
rect 15562 7188 15568 7200
rect 15427 7160 15568 7188
rect 15427 7157 15439 7160
rect 15381 7151 15439 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 18782 7148 18788 7200
rect 18840 7188 18846 7200
rect 18969 7191 19027 7197
rect 18969 7188 18981 7191
rect 18840 7160 18981 7188
rect 18840 7148 18846 7160
rect 18969 7157 18981 7160
rect 19015 7188 19027 7191
rect 19260 7188 19288 7219
rect 19015 7160 19288 7188
rect 19015 7157 19027 7160
rect 18969 7151 19027 7157
rect 1104 7098 21436 7120
rect 1104 7046 8497 7098
rect 8549 7046 8561 7098
rect 8613 7046 8625 7098
rect 8677 7046 8689 7098
rect 8741 7046 16012 7098
rect 16064 7046 16076 7098
rect 16128 7046 16140 7098
rect 16192 7046 16204 7098
rect 16256 7046 21436 7098
rect 1104 7024 21436 7046
rect 1397 6987 1455 6993
rect 1397 6953 1409 6987
rect 1443 6984 1455 6987
rect 2222 6984 2228 6996
rect 1443 6956 2228 6984
rect 1443 6953 1455 6956
rect 1397 6947 1455 6953
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 7558 6984 7564 6996
rect 7519 6956 7564 6984
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 8711 6987 8769 6993
rect 8711 6984 8723 6987
rect 7800 6956 8723 6984
rect 7800 6944 7806 6956
rect 8711 6953 8723 6956
rect 8757 6953 8769 6987
rect 8711 6947 8769 6953
rect 16255 6987 16313 6993
rect 16255 6953 16267 6987
rect 16301 6984 16313 6987
rect 16390 6984 16396 6996
rect 16301 6956 16396 6984
rect 16301 6953 16313 6956
rect 16255 6947 16313 6953
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 18874 6984 18880 6996
rect 18835 6956 18880 6984
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 1946 6916 1952 6928
rect 1907 6888 1952 6916
rect 1946 6876 1952 6888
rect 2004 6876 2010 6928
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 4212 6888 4257 6916
rect 4212 6876 4218 6888
rect 11146 6876 11152 6928
rect 11204 6916 11210 6928
rect 11333 6919 11391 6925
rect 11333 6916 11345 6919
rect 11204 6888 11345 6916
rect 11204 6876 11210 6888
rect 11333 6885 11345 6888
rect 11379 6885 11391 6919
rect 19242 6916 19248 6928
rect 19203 6888 19248 6916
rect 11333 6879 11391 6885
rect 19242 6876 19248 6888
rect 19300 6876 19306 6928
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2498 6848 2504 6860
rect 2455 6820 2504 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 8640 6851 8698 6857
rect 8640 6817 8652 6851
rect 8686 6848 8698 6851
rect 8846 6848 8852 6860
rect 8686 6820 8852 6848
rect 8686 6817 8698 6820
rect 8640 6811 8698 6817
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 12872 6851 12930 6857
rect 12872 6817 12884 6851
rect 12918 6848 12930 6851
rect 13078 6848 13084 6860
rect 12918 6820 13084 6848
rect 12918 6817 12930 6820
rect 12872 6811 12930 6817
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 13884 6851 13942 6857
rect 13884 6817 13896 6851
rect 13930 6848 13942 6851
rect 14550 6848 14556 6860
rect 13930 6820 14556 6848
rect 13930 6817 13942 6820
rect 13884 6811 13942 6817
rect 14550 6808 14556 6820
rect 14608 6808 14614 6860
rect 16184 6851 16242 6857
rect 16184 6817 16196 6851
rect 16230 6848 16242 6851
rect 16482 6848 16488 6860
rect 16230 6820 16488 6848
rect 16230 6817 16242 6820
rect 16184 6811 16242 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 5718 6780 5724 6792
rect 5679 6752 5724 6780
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12710 6780 12716 6792
rect 12023 6752 12716 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 17678 6780 17684 6792
rect 17639 6752 17684 6780
rect 17678 6740 17684 6752
rect 17736 6780 17742 6792
rect 19521 6783 19579 6789
rect 17736 6752 18920 6780
rect 17736 6740 17742 6752
rect 4709 6715 4767 6721
rect 4709 6681 4721 6715
rect 4755 6712 4767 6715
rect 6270 6712 6276 6724
rect 4755 6684 6276 6712
rect 4755 6681 4767 6684
rect 4709 6675 4767 6681
rect 6270 6672 6276 6684
rect 6328 6672 6334 6724
rect 18230 6712 18236 6724
rect 18191 6684 18236 6712
rect 18230 6672 18236 6684
rect 18288 6672 18294 6724
rect 18892 6712 18920 6752
rect 19521 6749 19533 6783
rect 19567 6749 19579 6783
rect 19521 6743 19579 6749
rect 19426 6712 19432 6724
rect 18892 6684 19432 6712
rect 19426 6672 19432 6684
rect 19484 6712 19490 6724
rect 19536 6712 19564 6743
rect 19484 6684 19564 6712
rect 19484 6672 19490 6684
rect 2547 6647 2605 6653
rect 2547 6613 2559 6647
rect 2593 6644 2605 6647
rect 2774 6644 2780 6656
rect 2593 6616 2780 6644
rect 2593 6613 2605 6616
rect 2547 6607 2605 6613
rect 2774 6604 2780 6616
rect 2832 6644 2838 6656
rect 2869 6647 2927 6653
rect 2869 6644 2881 6647
rect 2832 6616 2881 6644
rect 2832 6604 2838 6616
rect 2869 6613 2881 6616
rect 2915 6613 2927 6647
rect 2869 6607 2927 6613
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 12943 6647 13001 6653
rect 12943 6644 12955 6647
rect 11756 6616 12955 6644
rect 11756 6604 11762 6616
rect 12943 6613 12955 6616
rect 12989 6613 13001 6647
rect 12943 6607 13001 6613
rect 13446 6604 13452 6656
rect 13504 6644 13510 6656
rect 13955 6647 14013 6653
rect 13955 6644 13967 6647
rect 13504 6616 13967 6644
rect 13504 6604 13510 6616
rect 13955 6613 13967 6616
rect 14001 6613 14013 6647
rect 13955 6607 14013 6613
rect 1104 6554 21436 6576
rect 1104 6502 4739 6554
rect 4791 6502 4803 6554
rect 4855 6502 4867 6554
rect 4919 6502 4931 6554
rect 4983 6502 12255 6554
rect 12307 6502 12319 6554
rect 12371 6502 12383 6554
rect 12435 6502 12447 6554
rect 12499 6502 19770 6554
rect 19822 6502 19834 6554
rect 19886 6502 19898 6554
rect 19950 6502 19962 6554
rect 20014 6502 21436 6554
rect 1104 6480 21436 6502
rect 2498 6440 2504 6452
rect 2459 6412 2504 6440
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4212 6412 4257 6440
rect 4212 6400 4218 6412
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 11241 6443 11299 6449
rect 11241 6440 11253 6443
rect 11204 6412 11253 6440
rect 11204 6400 11210 6412
rect 11241 6409 11253 6412
rect 11287 6409 11299 6443
rect 11241 6403 11299 6409
rect 12897 6443 12955 6449
rect 12897 6409 12909 6443
rect 12943 6440 12955 6443
rect 13078 6440 13084 6452
rect 12943 6412 13084 6440
rect 12943 6409 12955 6412
rect 12897 6403 12955 6409
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 17678 6440 17684 6452
rect 17639 6412 17684 6440
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 18187 6443 18245 6449
rect 18187 6409 18199 6443
rect 18233 6440 18245 6443
rect 19058 6440 19064 6452
rect 18233 6412 19064 6440
rect 18233 6409 18245 6412
rect 18187 6403 18245 6409
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 20073 6443 20131 6449
rect 20073 6440 20085 6443
rect 19300 6412 20085 6440
rect 19300 6400 19306 6412
rect 20073 6409 20085 6412
rect 20119 6409 20131 6443
rect 20073 6403 20131 6409
rect 2225 6375 2283 6381
rect 2225 6341 2237 6375
rect 2271 6372 2283 6375
rect 2682 6372 2688 6384
rect 2271 6344 2688 6372
rect 2271 6341 2283 6344
rect 2225 6335 2283 6341
rect 1724 6239 1782 6245
rect 1724 6205 1736 6239
rect 1770 6236 1782 6239
rect 2240 6236 2268 6335
rect 2682 6332 2688 6344
rect 2740 6332 2746 6384
rect 5718 6372 5724 6384
rect 5631 6344 5724 6372
rect 5718 6332 5724 6344
rect 5776 6372 5782 6384
rect 5776 6344 13676 6372
rect 5776 6332 5782 6344
rect 13648 6316 13676 6344
rect 2774 6304 2780 6316
rect 2735 6276 2780 6304
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 4338 6264 4344 6316
rect 4396 6304 4402 6316
rect 4571 6307 4629 6313
rect 4571 6304 4583 6307
rect 4396 6276 4583 6304
rect 4396 6264 4402 6276
rect 4571 6273 4583 6276
rect 4617 6273 4629 6307
rect 4571 6267 4629 6273
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 8573 6307 8631 6313
rect 8573 6304 8585 6307
rect 8444 6276 8585 6304
rect 8444 6264 8450 6276
rect 8573 6273 8585 6276
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6304 13323 6307
rect 13446 6304 13452 6316
rect 13311 6276 13452 6304
rect 13311 6273 13323 6276
rect 13265 6267 13323 6273
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 13630 6264 13636 6316
rect 13688 6304 13694 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 13688 6276 13737 6304
rect 13688 6264 13694 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 19426 6304 19432 6316
rect 19387 6276 19432 6304
rect 13725 6267 13783 6273
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 1770 6208 2268 6236
rect 4484 6239 4542 6245
rect 1770 6205 1782 6208
rect 1724 6199 1782 6205
rect 4484 6205 4496 6239
rect 4530 6236 4542 6239
rect 18116 6239 18174 6245
rect 4530 6208 5028 6236
rect 4530 6205 4542 6208
rect 4484 6199 4542 6205
rect 1811 6171 1869 6177
rect 1811 6137 1823 6171
rect 1857 6168 1869 6171
rect 3234 6168 3240 6180
rect 1857 6140 3240 6168
rect 1857 6137 1869 6140
rect 1811 6131 1869 6137
rect 3234 6128 3240 6140
rect 3292 6128 3298 6180
rect 3418 6168 3424 6180
rect 3379 6140 3424 6168
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 5000 6109 5028 6208
rect 18116 6205 18128 6239
rect 18162 6236 18174 6239
rect 18162 6208 18644 6236
rect 18162 6205 18174 6208
rect 18116 6199 18174 6205
rect 8297 6171 8355 6177
rect 8297 6137 8309 6171
rect 8343 6137 8355 6171
rect 10137 6171 10195 6177
rect 10137 6168 10149 6171
rect 8297 6131 8355 6137
rect 9876 6140 10149 6168
rect 4985 6103 5043 6109
rect 4985 6069 4997 6103
rect 5031 6100 5043 6103
rect 5074 6100 5080 6112
rect 5031 6072 5080 6100
rect 5031 6069 5043 6072
rect 4985 6063 5043 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 8018 6100 8024 6112
rect 7979 6072 8024 6100
rect 8018 6060 8024 6072
rect 8076 6100 8082 6112
rect 8312 6100 8340 6131
rect 9876 6112 9904 6140
rect 10137 6137 10149 6140
rect 10183 6137 10195 6171
rect 10137 6131 10195 6137
rect 10781 6171 10839 6177
rect 10781 6137 10793 6171
rect 10827 6168 10839 6171
rect 11054 6168 11060 6180
rect 10827 6140 11060 6168
rect 10827 6137 10839 6140
rect 10781 6131 10839 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 18616 6112 18644 6208
rect 18969 6171 19027 6177
rect 18969 6137 18981 6171
rect 19015 6168 19027 6171
rect 19150 6168 19156 6180
rect 19015 6140 19156 6168
rect 19015 6137 19027 6140
rect 18969 6131 19027 6137
rect 19150 6128 19156 6140
rect 19208 6128 19214 6180
rect 8076 6072 8340 6100
rect 8076 6060 8082 6072
rect 8846 6060 8852 6112
rect 8904 6100 8910 6112
rect 9217 6103 9275 6109
rect 9217 6100 9229 6103
rect 8904 6072 9229 6100
rect 8904 6060 8910 6072
rect 9217 6069 9229 6072
rect 9263 6069 9275 6103
rect 9858 6100 9864 6112
rect 9819 6072 9864 6100
rect 9217 6063 9275 6069
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 14461 6103 14519 6109
rect 14461 6069 14473 6103
rect 14507 6100 14519 6103
rect 14550 6100 14556 6112
rect 14507 6072 14556 6100
rect 14507 6069 14519 6072
rect 14461 6063 14519 6069
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 16209 6103 16267 6109
rect 16209 6069 16221 6103
rect 16255 6100 16267 6103
rect 16482 6100 16488 6112
rect 16255 6072 16488 6100
rect 16255 6069 16267 6072
rect 16209 6063 16267 6069
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 18598 6100 18604 6112
rect 18559 6072 18604 6100
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 1104 6010 21436 6032
rect 1104 5958 8497 6010
rect 8549 5958 8561 6010
rect 8613 5958 8625 6010
rect 8677 5958 8689 6010
rect 8741 5958 16012 6010
rect 16064 5958 16076 6010
rect 16128 5958 16140 6010
rect 16192 5958 16204 6010
rect 16256 5958 21436 6010
rect 1104 5936 21436 5958
rect 7699 5899 7757 5905
rect 7699 5865 7711 5899
rect 7745 5896 7757 5899
rect 8018 5896 8024 5908
rect 7745 5868 8024 5896
rect 7745 5865 7757 5868
rect 7699 5859 7757 5865
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 8711 5899 8769 5905
rect 8711 5865 8723 5899
rect 8757 5896 8769 5899
rect 9858 5896 9864 5908
rect 8757 5868 9864 5896
rect 8757 5865 8769 5868
rect 8711 5859 8769 5865
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 3418 5828 3424 5840
rect 2823 5800 3424 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 3418 5788 3424 5800
rect 3476 5788 3482 5840
rect 5261 5831 5319 5837
rect 5261 5797 5273 5831
rect 5307 5828 5319 5831
rect 5718 5828 5724 5840
rect 5307 5800 5724 5828
rect 5307 5797 5319 5800
rect 5261 5791 5319 5797
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 10137 5831 10195 5837
rect 10137 5828 10149 5831
rect 9824 5800 10149 5828
rect 9824 5788 9830 5800
rect 10137 5797 10149 5800
rect 10183 5797 10195 5831
rect 11698 5828 11704 5840
rect 11659 5800 11704 5828
rect 10137 5791 10195 5797
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 5350 5720 5356 5772
rect 5408 5760 5414 5772
rect 6546 5760 6552 5772
rect 6604 5769 6610 5772
rect 6604 5763 6642 5769
rect 5408 5732 6552 5760
rect 5408 5720 5414 5732
rect 6546 5720 6552 5732
rect 6630 5729 6642 5763
rect 6604 5723 6642 5729
rect 7628 5763 7686 5769
rect 7628 5729 7640 5763
rect 7674 5760 7686 5763
rect 7834 5760 7840 5772
rect 7674 5732 7840 5760
rect 7674 5729 7686 5732
rect 7628 5723 7686 5729
rect 6604 5720 6610 5723
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 8608 5763 8666 5769
rect 8608 5760 8620 5763
rect 7984 5732 8620 5760
rect 7984 5720 7990 5732
rect 8608 5729 8620 5732
rect 8654 5760 8666 5763
rect 9122 5760 9128 5772
rect 8654 5732 9128 5760
rect 8654 5729 8666 5732
rect 8608 5723 8666 5729
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 13078 5720 13084 5772
rect 13136 5760 13142 5772
rect 13208 5763 13266 5769
rect 13208 5760 13220 5763
rect 13136 5732 13220 5760
rect 13136 5720 13142 5732
rect 13208 5729 13220 5732
rect 13254 5729 13266 5763
rect 13208 5723 13266 5729
rect 15816 5763 15874 5769
rect 15816 5729 15828 5763
rect 15862 5760 15874 5763
rect 16666 5760 16672 5772
rect 15862 5732 16672 5760
rect 15862 5729 15874 5732
rect 15816 5723 15874 5729
rect 16666 5720 16672 5732
rect 16724 5720 16730 5772
rect 2130 5692 2136 5704
rect 2091 5664 2136 5692
rect 2130 5652 2136 5664
rect 2188 5652 2194 5704
rect 4614 5692 4620 5704
rect 4575 5664 4620 5692
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 11054 5692 11060 5704
rect 10827 5664 11060 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 11054 5652 11060 5664
rect 11112 5692 11118 5704
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 11112 5664 11989 5692
rect 11112 5652 11118 5664
rect 11977 5661 11989 5664
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 17865 5695 17923 5701
rect 17865 5661 17877 5695
rect 17911 5692 17923 5695
rect 18966 5692 18972 5704
rect 17911 5664 18972 5692
rect 17911 5661 17923 5664
rect 17865 5655 17923 5661
rect 18966 5652 18972 5664
rect 19024 5652 19030 5704
rect 19426 5692 19432 5704
rect 19387 5664 19432 5692
rect 19426 5652 19432 5664
rect 19484 5652 19490 5704
rect 6687 5559 6745 5565
rect 6687 5525 6699 5559
rect 6733 5556 6745 5559
rect 7650 5556 7656 5568
rect 6733 5528 7656 5556
rect 6733 5525 6745 5528
rect 6687 5519 6745 5525
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 12618 5516 12624 5568
rect 12676 5556 12682 5568
rect 13311 5559 13369 5565
rect 13311 5556 13323 5559
rect 12676 5528 13323 5556
rect 12676 5516 12682 5528
rect 13311 5525 13323 5528
rect 13357 5525 13369 5559
rect 13311 5519 13369 5525
rect 15654 5516 15660 5568
rect 15712 5556 15718 5568
rect 15887 5559 15945 5565
rect 15887 5556 15899 5559
rect 15712 5528 15899 5556
rect 15712 5516 15718 5528
rect 15887 5525 15899 5528
rect 15933 5525 15945 5559
rect 15887 5519 15945 5525
rect 1104 5466 21436 5488
rect 1104 5414 4739 5466
rect 4791 5414 4803 5466
rect 4855 5414 4867 5466
rect 4919 5414 4931 5466
rect 4983 5414 12255 5466
rect 12307 5414 12319 5466
rect 12371 5414 12383 5466
rect 12435 5414 12447 5466
rect 12499 5414 19770 5466
rect 19822 5414 19834 5466
rect 19886 5414 19898 5466
rect 19950 5414 19962 5466
rect 20014 5414 21436 5466
rect 1104 5392 21436 5414
rect 1535 5355 1593 5361
rect 1535 5321 1547 5355
rect 1581 5352 1593 5355
rect 2130 5352 2136 5364
rect 1581 5324 2136 5352
rect 1581 5321 1593 5324
rect 1535 5315 1593 5321
rect 2130 5312 2136 5324
rect 2188 5352 2194 5364
rect 2225 5355 2283 5361
rect 2225 5352 2237 5355
rect 2188 5324 2237 5352
rect 2188 5312 2194 5324
rect 2225 5321 2237 5324
rect 2271 5321 2283 5355
rect 2225 5315 2283 5321
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 3605 5355 3663 5361
rect 3605 5352 3617 5355
rect 3292 5324 3617 5352
rect 3292 5312 3298 5324
rect 3605 5321 3617 5324
rect 3651 5352 3663 5355
rect 3878 5352 3884 5364
rect 3651 5324 3884 5352
rect 3651 5321 3663 5324
rect 3605 5315 3663 5321
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 6546 5352 6552 5364
rect 6507 5324 6552 5352
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 9122 5352 9128 5364
rect 9083 5324 9128 5352
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 9861 5355 9919 5361
rect 9861 5352 9873 5355
rect 9824 5324 9873 5352
rect 9824 5312 9830 5324
rect 9861 5321 9873 5324
rect 9907 5321 9919 5355
rect 11054 5352 11060 5364
rect 11015 5324 11060 5352
rect 9861 5315 9919 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11698 5352 11704 5364
rect 11659 5324 11704 5352
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 13078 5312 13084 5364
rect 13136 5352 13142 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 13136 5324 13461 5352
rect 13136 5312 13142 5324
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 16666 5352 16672 5364
rect 16627 5324 16672 5352
rect 13449 5315 13507 5321
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 18966 5312 18972 5364
rect 19024 5352 19030 5364
rect 19705 5355 19763 5361
rect 19705 5352 19717 5355
rect 19024 5324 19717 5352
rect 19024 5312 19030 5324
rect 19705 5321 19717 5324
rect 19751 5321 19763 5355
rect 19705 5315 19763 5321
rect 3145 5287 3203 5293
rect 3145 5284 3157 5287
rect 2751 5256 3157 5284
rect 1210 5176 1216 5228
rect 1268 5216 1274 5228
rect 1857 5219 1915 5225
rect 1857 5216 1869 5219
rect 1268 5188 1869 5216
rect 1268 5176 1274 5188
rect 1479 5157 1507 5188
rect 1857 5185 1869 5188
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 2751 5157 2779 5256
rect 3145 5253 3157 5256
rect 3191 5284 3203 5287
rect 3326 5284 3332 5296
rect 3191 5256 3332 5284
rect 3191 5253 3203 5256
rect 3145 5247 3203 5253
rect 3326 5244 3332 5256
rect 3384 5244 3390 5296
rect 11072 5284 11100 5312
rect 10152 5256 11100 5284
rect 19429 5287 19487 5293
rect 10152 5225 10180 5256
rect 19429 5253 19441 5287
rect 19475 5284 19487 5287
rect 20162 5284 20168 5296
rect 19475 5256 20168 5284
rect 19475 5253 19487 5256
rect 19429 5247 19487 5253
rect 2823 5219 2881 5225
rect 2823 5185 2835 5219
rect 2869 5216 2881 5219
rect 6181 5219 6239 5225
rect 6181 5216 6193 5219
rect 2869 5188 6193 5216
rect 2869 5185 2881 5188
rect 2823 5179 2881 5185
rect 6181 5185 6193 5188
rect 6227 5216 6239 5219
rect 6917 5219 6975 5225
rect 6917 5216 6929 5219
rect 6227 5188 6929 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6917 5185 6929 5188
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10410 5216 10416 5228
rect 10371 5188 10416 5216
rect 10137 5179 10195 5185
rect 10410 5176 10416 5188
rect 10468 5176 10474 5228
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 12529 5219 12587 5225
rect 12529 5216 12541 5219
rect 12299 5188 12541 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12529 5185 12541 5188
rect 12575 5216 12587 5219
rect 12618 5216 12624 5228
rect 12575 5188 12624 5216
rect 12575 5185 12587 5188
rect 12529 5179 12587 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 12805 5219 12863 5225
rect 12805 5216 12817 5219
rect 12768 5188 12817 5216
rect 12768 5176 12774 5188
rect 12805 5185 12817 5188
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 15473 5219 15531 5225
rect 15473 5185 15485 5219
rect 15519 5216 15531 5219
rect 15654 5216 15660 5228
rect 15519 5188 15660 5216
rect 15519 5185 15531 5188
rect 15473 5179 15531 5185
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 19015 5219 19073 5225
rect 19015 5185 19027 5219
rect 19061 5216 19073 5219
rect 19150 5216 19156 5228
rect 19061 5188 19156 5216
rect 19061 5185 19073 5188
rect 19015 5179 19073 5185
rect 19150 5176 19156 5188
rect 19208 5176 19214 5228
rect 1464 5151 1522 5157
rect 1464 5117 1476 5151
rect 1510 5117 1522 5151
rect 1464 5111 1522 5117
rect 2736 5151 2794 5157
rect 2736 5117 2748 5151
rect 2782 5117 2794 5151
rect 2736 5111 2794 5117
rect 5074 5108 5080 5160
rect 5132 5148 5138 5160
rect 5420 5151 5478 5157
rect 5420 5148 5432 5151
rect 5132 5120 5432 5148
rect 5132 5108 5138 5120
rect 5420 5117 5432 5120
rect 5466 5148 5478 5151
rect 8732 5151 8790 5157
rect 5466 5120 5856 5148
rect 5466 5117 5478 5120
rect 5420 5111 5478 5117
rect 3878 5080 3884 5092
rect 3839 5052 3884 5080
rect 3878 5040 3884 5052
rect 3936 5040 3942 5092
rect 4522 5080 4528 5092
rect 4483 5052 4528 5080
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 5828 5024 5856 5120
rect 8732 5117 8744 5151
rect 8778 5148 8790 5151
rect 14068 5151 14126 5157
rect 14068 5148 14080 5151
rect 8778 5120 9444 5148
rect 8778 5117 8790 5120
rect 8732 5111 8790 5117
rect 7561 5083 7619 5089
rect 7561 5049 7573 5083
rect 7607 5080 7619 5083
rect 7926 5080 7932 5092
rect 7607 5052 7932 5080
rect 7607 5049 7619 5052
rect 7561 5043 7619 5049
rect 7926 5040 7932 5052
rect 7984 5040 7990 5092
rect 9416 5024 9444 5120
rect 13786 5120 14080 5148
rect 4798 5012 4804 5024
rect 4759 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 5491 5015 5549 5021
rect 5491 4981 5503 5015
rect 5537 5012 5549 5015
rect 5718 5012 5724 5024
rect 5537 4984 5724 5012
rect 5537 4981 5549 4984
rect 5491 4975 5549 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 7834 5012 7840 5024
rect 5868 4984 5913 5012
rect 7795 4984 7840 5012
rect 5868 4972 5874 4984
rect 7834 4972 7840 4984
rect 7892 4972 7898 5024
rect 8803 5015 8861 5021
rect 8803 4981 8815 5015
rect 8849 5012 8861 5015
rect 8938 5012 8944 5024
rect 8849 4984 8944 5012
rect 8849 4981 8861 4984
rect 8803 4975 8861 4981
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 9398 4972 9404 5024
rect 9456 5012 9462 5024
rect 9493 5015 9551 5021
rect 9493 5012 9505 5015
rect 9456 4984 9505 5012
rect 9456 4972 9462 4984
rect 9493 4981 9505 4984
rect 9539 4981 9551 5015
rect 9493 4975 9551 4981
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 13786 5012 13814 5120
rect 14068 5117 14080 5120
rect 14114 5148 14126 5151
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 14114 5120 14473 5148
rect 14114 5117 14126 5120
rect 14068 5111 14126 5117
rect 14461 5117 14473 5120
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 18598 5108 18604 5160
rect 18656 5148 18662 5160
rect 18928 5151 18986 5157
rect 18928 5148 18940 5151
rect 18656 5120 18940 5148
rect 18656 5108 18662 5120
rect 18928 5117 18940 5120
rect 18974 5148 18986 5151
rect 19444 5148 19472 5247
rect 20162 5244 20168 5256
rect 20220 5244 20226 5296
rect 18974 5120 19472 5148
rect 18974 5117 18986 5120
rect 18928 5111 18986 5117
rect 16298 5080 16304 5092
rect 16259 5052 16304 5080
rect 16298 5040 16304 5052
rect 16356 5040 16362 5092
rect 10744 4984 13814 5012
rect 14139 5015 14197 5021
rect 10744 4972 10750 4984
rect 14139 4981 14151 5015
rect 14185 5012 14197 5015
rect 15378 5012 15384 5024
rect 14185 4984 15384 5012
rect 14185 4981 14197 4984
rect 14139 4975 14197 4981
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 1104 4922 21436 4944
rect 1104 4870 8497 4922
rect 8549 4870 8561 4922
rect 8613 4870 8625 4922
rect 8677 4870 8689 4922
rect 8741 4870 16012 4922
rect 16064 4870 16076 4922
rect 16128 4870 16140 4922
rect 16192 4870 16204 4922
rect 16256 4870 21436 4922
rect 1104 4848 21436 4870
rect 3099 4811 3157 4817
rect 3099 4777 3111 4811
rect 3145 4808 3157 4811
rect 4798 4808 4804 4820
rect 3145 4780 4804 4808
rect 3145 4777 3157 4780
rect 3099 4771 3157 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 6546 4768 6552 4820
rect 6604 4808 6610 4820
rect 10686 4808 10692 4820
rect 6604 4780 10692 4808
rect 6604 4768 6610 4780
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 6089 4743 6147 4749
rect 6089 4740 6101 4743
rect 5776 4712 6101 4740
rect 5776 4700 5782 4712
rect 6089 4709 6101 4712
rect 6135 4740 6147 4743
rect 6178 4740 6184 4752
rect 6135 4712 6184 4740
rect 6135 4709 6147 4712
rect 6089 4703 6147 4709
rect 6178 4700 6184 4712
rect 6236 4700 6242 4752
rect 7650 4740 7656 4752
rect 7611 4712 7656 4740
rect 7650 4700 7656 4712
rect 7708 4700 7714 4752
rect 10410 4740 10416 4752
rect 10371 4712 10416 4740
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 12621 4743 12679 4749
rect 12621 4709 12633 4743
rect 12667 4740 12679 4743
rect 12710 4740 12716 4752
rect 12667 4712 12716 4740
rect 12667 4709 12679 4712
rect 12621 4703 12679 4709
rect 12710 4700 12716 4712
rect 12768 4740 12774 4752
rect 12897 4743 12955 4749
rect 12897 4740 12909 4743
rect 12768 4712 12909 4740
rect 12768 4700 12774 4712
rect 12897 4709 12909 4712
rect 12943 4709 12955 4743
rect 15378 4740 15384 4752
rect 15339 4712 15384 4740
rect 12897 4703 12955 4709
rect 15378 4700 15384 4712
rect 15436 4700 15442 4752
rect 15746 4700 15752 4752
rect 15804 4740 15810 4752
rect 16025 4743 16083 4749
rect 16025 4740 16037 4743
rect 15804 4712 16037 4740
rect 15804 4700 15810 4712
rect 16025 4709 16037 4712
rect 16071 4740 16083 4743
rect 16298 4740 16304 4752
rect 16071 4712 16304 4740
rect 16071 4709 16083 4712
rect 16025 4703 16083 4709
rect 16298 4700 16304 4712
rect 16356 4700 16362 4752
rect 18782 4700 18788 4752
rect 18840 4740 18846 4752
rect 19981 4743 20039 4749
rect 19981 4740 19993 4743
rect 18840 4712 19993 4740
rect 18840 4700 18846 4712
rect 19981 4709 19993 4712
rect 20027 4709 20039 4743
rect 19981 4703 20039 4709
rect 16888 4675 16946 4681
rect 16888 4641 16900 4675
rect 16934 4641 16946 4675
rect 16888 4635 16946 4641
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 3050 4604 3056 4616
rect 2915 4576 3056 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4604 4583 4607
rect 4614 4604 4620 4616
rect 4571 4576 4620 4604
rect 4571 4573 4583 4576
rect 4525 4567 4583 4573
rect 4614 4564 4620 4576
rect 4672 4604 4678 4616
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 4672 4576 6377 4604
rect 4672 4564 4678 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 7926 4604 7932 4616
rect 7887 4576 7932 4604
rect 6365 4567 6423 4573
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 9766 4604 9772 4616
rect 9727 4576 9772 4604
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 11974 4604 11980 4616
rect 11887 4576 11980 4604
rect 11974 4564 11980 4576
rect 12032 4604 12038 4616
rect 13449 4607 13507 4613
rect 13449 4604 13461 4607
rect 12032 4576 13461 4604
rect 12032 4564 12038 4576
rect 13449 4573 13461 4576
rect 13495 4573 13507 4607
rect 13449 4567 13507 4573
rect 16903 4548 16931 4635
rect 19334 4604 19340 4616
rect 19295 4576 19340 4604
rect 19334 4564 19340 4576
rect 19392 4564 19398 4616
rect 5074 4536 5080 4548
rect 5035 4508 5080 4536
rect 5074 4496 5080 4508
rect 5132 4496 5138 4548
rect 16850 4496 16856 4548
rect 16908 4508 16931 4548
rect 16908 4496 16914 4508
rect 16298 4428 16304 4480
rect 16356 4468 16362 4480
rect 16991 4471 17049 4477
rect 16991 4468 17003 4471
rect 16356 4440 17003 4468
rect 16356 4428 16362 4440
rect 16991 4437 17003 4440
rect 17037 4437 17049 4471
rect 16991 4431 17049 4437
rect 1104 4378 21436 4400
rect 1104 4326 4739 4378
rect 4791 4326 4803 4378
rect 4855 4326 4867 4378
rect 4919 4326 4931 4378
rect 4983 4326 12255 4378
rect 12307 4326 12319 4378
rect 12371 4326 12383 4378
rect 12435 4326 12447 4378
rect 12499 4326 19770 4378
rect 19822 4326 19834 4378
rect 19886 4326 19898 4378
rect 19950 4326 19962 4378
rect 20014 4326 21436 4378
rect 1104 4304 21436 4326
rect 4614 4224 4620 4276
rect 4672 4264 4678 4276
rect 4801 4267 4859 4273
rect 4801 4264 4813 4267
rect 4672 4236 4813 4264
rect 4672 4224 4678 4236
rect 4801 4233 4813 4236
rect 4847 4233 4859 4267
rect 6178 4264 6184 4276
rect 6139 4236 6184 4264
rect 4801 4227 4859 4233
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 7650 4224 7656 4276
rect 7708 4264 7714 4276
rect 8021 4267 8079 4273
rect 8021 4264 8033 4267
rect 7708 4236 8033 4264
rect 7708 4224 7714 4236
rect 8021 4233 8033 4236
rect 8067 4233 8079 4267
rect 9677 4267 9735 4273
rect 9677 4264 9689 4267
rect 8021 4227 8079 4233
rect 9048 4236 9689 4264
rect 4433 4199 4491 4205
rect 4433 4165 4445 4199
rect 4479 4196 4491 4199
rect 4632 4196 4660 4224
rect 4479 4168 4660 4196
rect 4479 4165 4491 4168
rect 4433 4159 4491 4165
rect 7926 4156 7932 4208
rect 7984 4196 7990 4208
rect 9048 4196 9076 4236
rect 9677 4233 9689 4236
rect 9723 4264 9735 4267
rect 9766 4264 9772 4276
rect 9723 4236 9772 4264
rect 9723 4233 9735 4236
rect 9677 4227 9735 4233
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 11974 4264 11980 4276
rect 11935 4236 11980 4264
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 15378 4264 15384 4276
rect 15339 4236 15384 4264
rect 15378 4224 15384 4236
rect 15436 4224 15442 4276
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 19429 4267 19487 4273
rect 19429 4264 19441 4267
rect 19392 4236 19441 4264
rect 19392 4224 19398 4236
rect 19429 4233 19441 4236
rect 19475 4264 19487 4267
rect 19751 4267 19809 4273
rect 19751 4264 19763 4267
rect 19475 4236 19763 4264
rect 19475 4233 19487 4236
rect 19429 4227 19487 4233
rect 19751 4233 19763 4236
rect 19797 4233 19809 4267
rect 19751 4227 19809 4233
rect 7984 4168 9076 4196
rect 7984 4156 7990 4168
rect 1854 4128 1860 4140
rect 1815 4100 1860 4128
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 9048 4137 9076 4168
rect 10873 4199 10931 4205
rect 10873 4165 10885 4199
rect 10919 4196 10931 4199
rect 11698 4196 11704 4208
rect 10919 4168 11704 4196
rect 10919 4165 10931 4168
rect 10873 4159 10931 4165
rect 11698 4156 11704 4168
rect 11756 4156 11762 4208
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 9011 4100 9045 4128
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 12710 4128 12716 4140
rect 12575 4100 12716 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 14458 4128 14464 4140
rect 14083 4100 14464 4128
rect 1464 4063 1522 4069
rect 1464 4029 1476 4063
rect 1510 4060 1522 4063
rect 1872 4060 1900 4088
rect 7282 4069 7288 4072
rect 7260 4063 7288 4069
rect 7260 4060 7272 4063
rect 1510 4032 1900 4060
rect 7195 4032 7272 4060
rect 1510 4029 1522 4032
rect 1464 4023 1522 4029
rect 7260 4029 7272 4032
rect 7340 4060 7346 4072
rect 10686 4060 10692 4072
rect 7340 4032 7788 4060
rect 10599 4032 10692 4060
rect 7260 4023 7288 4029
rect 7282 4020 7288 4023
rect 7340 4020 7346 4032
rect 3881 3995 3939 4001
rect 3881 3992 3893 3995
rect 3620 3964 3893 3992
rect 3620 3936 3648 3964
rect 3881 3961 3893 3964
rect 3927 3961 3939 3995
rect 3881 3955 3939 3961
rect 7760 3936 7788 4032
rect 10686 4020 10692 4032
rect 10744 4060 10750 4072
rect 14083 4069 14111 4100
rect 14458 4088 14464 4100
rect 14516 4088 14522 4140
rect 19153 4131 19211 4137
rect 19153 4128 19165 4131
rect 18683 4100 19165 4128
rect 18683 4069 18711 4100
rect 19153 4097 19165 4100
rect 19199 4128 19211 4131
rect 20254 4128 20260 4140
rect 19199 4100 20260 4128
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 11241 4063 11299 4069
rect 11241 4060 11253 4063
rect 10744 4032 11253 4060
rect 10744 4020 10750 4032
rect 11241 4029 11253 4032
rect 11287 4029 11299 4063
rect 11241 4023 11299 4029
rect 14068 4063 14126 4069
rect 14068 4029 14080 4063
rect 14114 4029 14126 4063
rect 14068 4023 14126 4029
rect 18668 4063 18726 4069
rect 18668 4029 18680 4063
rect 18714 4029 18726 4063
rect 18668 4023 18726 4029
rect 19680 4063 19738 4069
rect 19680 4029 19692 4063
rect 19726 4060 19738 4063
rect 19726 4032 20208 4060
rect 19726 4029 19738 4032
rect 19680 4023 19738 4029
rect 8573 3995 8631 4001
rect 8573 3961 8585 3995
rect 8619 3992 8631 3995
rect 8757 3995 8815 4001
rect 8757 3992 8769 3995
rect 8619 3964 8769 3992
rect 8619 3961 8631 3964
rect 8573 3955 8631 3961
rect 8757 3961 8769 3964
rect 8803 3992 8815 3995
rect 8938 3992 8944 4004
rect 8803 3964 8944 3992
rect 8803 3961 8815 3964
rect 8757 3955 8815 3961
rect 8938 3952 8944 3964
rect 8996 3952 9002 4004
rect 13170 3992 13176 4004
rect 13131 3964 13176 3992
rect 13170 3952 13176 3964
rect 13228 3952 13234 4004
rect 15013 3995 15071 4001
rect 15013 3961 15025 3995
rect 15059 3992 15071 3995
rect 15746 3992 15752 4004
rect 15059 3964 15752 3992
rect 15059 3961 15071 3964
rect 15013 3955 15071 3961
rect 15746 3952 15752 3964
rect 15804 3952 15810 4004
rect 16393 3995 16451 4001
rect 16393 3961 16405 3995
rect 16439 3992 16451 3995
rect 16850 3992 16856 4004
rect 16439 3964 16856 3992
rect 16439 3961 16451 3964
rect 16393 3955 16451 3961
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 20180 3936 20208 4032
rect 1535 3927 1593 3933
rect 1535 3893 1547 3927
rect 1581 3924 1593 3927
rect 2130 3924 2136 3936
rect 1581 3896 2136 3924
rect 1581 3893 1593 3896
rect 1535 3887 1593 3893
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 3050 3924 3056 3936
rect 3011 3896 3056 3924
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 3602 3924 3608 3936
rect 3563 3896 3608 3924
rect 3602 3884 3608 3896
rect 3660 3884 3666 3936
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 7331 3927 7389 3933
rect 7331 3893 7343 3927
rect 7377 3924 7389 3927
rect 7558 3924 7564 3936
rect 7377 3896 7564 3924
rect 7377 3893 7389 3896
rect 7331 3887 7389 3893
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 7742 3924 7748 3936
rect 7703 3896 7748 3924
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 14139 3927 14197 3933
rect 14139 3924 14151 3927
rect 11296 3896 14151 3924
rect 11296 3884 11302 3896
rect 14139 3893 14151 3896
rect 14185 3893 14197 3927
rect 14139 3887 14197 3893
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 18739 3927 18797 3933
rect 18739 3924 18751 3927
rect 18564 3896 18751 3924
rect 18564 3884 18570 3896
rect 18739 3893 18751 3896
rect 18785 3893 18797 3927
rect 20162 3924 20168 3936
rect 20123 3896 20168 3924
rect 18739 3887 18797 3893
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 1104 3834 21436 3856
rect 1104 3782 8497 3834
rect 8549 3782 8561 3834
rect 8613 3782 8625 3834
rect 8677 3782 8689 3834
rect 8741 3782 16012 3834
rect 16064 3782 16076 3834
rect 16128 3782 16140 3834
rect 16192 3782 16204 3834
rect 16256 3782 21436 3834
rect 1104 3760 21436 3782
rect 2130 3652 2136 3664
rect 2091 3624 2136 3652
rect 2130 3612 2136 3624
rect 2188 3612 2194 3664
rect 7558 3652 7564 3664
rect 7519 3624 7564 3652
rect 7558 3612 7564 3624
rect 7616 3612 7622 3664
rect 10410 3652 10416 3664
rect 10371 3624 10416 3652
rect 10410 3612 10416 3624
rect 10468 3652 10474 3664
rect 10468 3624 12664 3652
rect 10468 3612 10474 3624
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 4522 3584 4528 3596
rect 4479 3556 4528 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 6362 3584 6368 3596
rect 6323 3556 6368 3584
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 11238 3584 11244 3596
rect 11199 3556 11244 3584
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11974 3544 11980 3596
rect 12032 3584 12038 3596
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 12032 3556 12357 3584
rect 12032 3544 12038 3556
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12636 3584 12664 3624
rect 13446 3584 13452 3596
rect 13504 3593 13510 3596
rect 13504 3587 13542 3593
rect 12636 3556 13452 3584
rect 12345 3547 12403 3553
rect 13446 3544 13452 3556
rect 13530 3553 13542 3587
rect 13504 3547 13542 3553
rect 13504 3544 13510 3547
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 19648 3587 19706 3593
rect 19648 3584 19660 3587
rect 19576 3556 19660 3584
rect 19576 3544 19582 3556
rect 19648 3553 19660 3556
rect 19694 3553 19706 3587
rect 19648 3547 19706 3553
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3516 2835 3519
rect 5442 3516 5448 3528
rect 2823 3488 5448 3516
rect 2823 3485 2835 3488
rect 2777 3479 2835 3485
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5994 3476 6000 3528
rect 6052 3516 6058 3528
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 6052 3488 7849 3516
rect 6052 3476 6058 3488
rect 7837 3485 7849 3488
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3516 9827 3519
rect 10042 3516 10048 3528
rect 9815 3488 10048 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 7852 3448 7880 3479
rect 10042 3476 10048 3488
rect 10100 3516 10106 3528
rect 15378 3516 15384 3528
rect 10100 3488 13814 3516
rect 15339 3488 15384 3516
rect 10100 3476 10106 3488
rect 12618 3448 12624 3460
rect 7852 3420 12624 3448
rect 12618 3408 12624 3420
rect 12676 3448 12682 3460
rect 12897 3451 12955 3457
rect 12897 3448 12909 3451
rect 12676 3420 12909 3448
rect 12676 3408 12682 3420
rect 12897 3417 12909 3420
rect 12943 3417 12955 3451
rect 13786 3448 13814 3488
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 15657 3519 15715 3525
rect 15657 3516 15669 3519
rect 15488 3488 15669 3516
rect 15488 3448 15516 3488
rect 15657 3485 15669 3488
rect 15703 3485 15715 3519
rect 16942 3516 16948 3528
rect 16903 3488 16948 3516
rect 15657 3479 15715 3485
rect 16942 3476 16948 3488
rect 17000 3476 17006 3528
rect 17218 3516 17224 3528
rect 17179 3488 17224 3516
rect 17218 3476 17224 3488
rect 17276 3476 17282 3528
rect 18414 3516 18420 3528
rect 18375 3488 18420 3516
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 13786 3420 15516 3448
rect 12897 3411 12955 3417
rect 4614 3389 4620 3392
rect 4571 3383 4620 3389
rect 4571 3380 4583 3383
rect 4527 3352 4583 3380
rect 4571 3349 4583 3352
rect 4617 3349 4620 3383
rect 4571 3343 4620 3349
rect 4614 3340 4620 3343
rect 4672 3380 4678 3392
rect 4893 3383 4951 3389
rect 4893 3380 4905 3383
rect 4672 3352 4905 3380
rect 4672 3340 4678 3352
rect 4893 3349 4905 3352
rect 4939 3349 4951 3383
rect 4893 3343 4951 3349
rect 6549 3383 6607 3389
rect 6549 3349 6561 3383
rect 6595 3380 6607 3383
rect 7006 3380 7012 3392
rect 6595 3352 7012 3380
rect 6595 3349 6607 3352
rect 6549 3343 6607 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 11425 3383 11483 3389
rect 11425 3349 11437 3383
rect 11471 3380 11483 3383
rect 12066 3380 12072 3392
rect 11471 3352 12072 3380
rect 11471 3349 11483 3352
rect 11425 3343 11483 3349
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 12529 3383 12587 3389
rect 12529 3349 12541 3383
rect 12575 3380 12587 3383
rect 12802 3380 12808 3392
rect 12575 3352 12808 3380
rect 12575 3349 12587 3352
rect 12529 3343 12587 3349
rect 12802 3340 12808 3352
rect 12860 3340 12866 3392
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 13587 3383 13645 3389
rect 13587 3380 13599 3383
rect 13044 3352 13599 3380
rect 13044 3340 13050 3352
rect 13587 3349 13599 3352
rect 13633 3349 13645 3383
rect 13587 3343 13645 3349
rect 19610 3340 19616 3392
rect 19668 3380 19674 3392
rect 19751 3383 19809 3389
rect 19751 3380 19763 3383
rect 19668 3352 19763 3380
rect 19668 3340 19674 3352
rect 19751 3349 19763 3352
rect 19797 3349 19809 3383
rect 19751 3343 19809 3349
rect 1104 3290 21436 3312
rect 1104 3238 4739 3290
rect 4791 3238 4803 3290
rect 4855 3238 4867 3290
rect 4919 3238 4931 3290
rect 4983 3238 12255 3290
rect 12307 3238 12319 3290
rect 12371 3238 12383 3290
rect 12435 3238 12447 3290
rect 12499 3238 19770 3290
rect 19822 3238 19834 3290
rect 19886 3238 19898 3290
rect 19950 3238 19962 3290
rect 20014 3238 21436 3290
rect 1104 3216 21436 3238
rect 2130 3176 2136 3188
rect 2091 3148 2136 3176
rect 2130 3136 2136 3148
rect 2188 3136 2194 3188
rect 3467 3179 3525 3185
rect 3467 3145 3479 3179
rect 3513 3176 3525 3179
rect 3602 3176 3608 3188
rect 3513 3148 3608 3176
rect 3513 3145 3525 3148
rect 3467 3139 3525 3145
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 5776 3148 6561 3176
rect 5776 3136 5782 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 2455 3111 2513 3117
rect 2455 3077 2467 3111
rect 2501 3108 2513 3111
rect 6181 3111 6239 3117
rect 6181 3108 6193 3111
rect 2501 3080 6193 3108
rect 2501 3077 2513 3080
rect 2455 3071 2513 3077
rect 6181 3077 6193 3080
rect 6227 3108 6239 3111
rect 6362 3108 6368 3120
rect 6227 3080 6368 3108
rect 6227 3077 6239 3080
rect 6181 3071 6239 3077
rect 6362 3068 6368 3080
rect 6420 3068 6426 3120
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 2399 3012 2881 3040
rect 2399 2981 2427 3012
rect 2869 3009 2881 3012
rect 2915 3040 2927 3043
rect 2915 3012 4154 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 2384 2975 2442 2981
rect 2384 2941 2396 2975
rect 2430 2941 2442 2975
rect 2384 2935 2442 2941
rect 3396 2975 3454 2981
rect 3396 2941 3408 2975
rect 3442 2972 3454 2975
rect 3442 2944 3924 2972
rect 3442 2941 3454 2944
rect 3396 2935 3454 2941
rect 3896 2848 3924 2944
rect 4126 2904 4154 3012
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 4672 3012 4813 3040
rect 4672 3000 4678 3012
rect 4801 3009 4813 3012
rect 4847 3009 4859 3043
rect 6564 3040 6592 3139
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7616 3148 7849 3176
rect 7616 3136 7622 3148
rect 7837 3145 7849 3148
rect 7883 3145 7895 3179
rect 10042 3176 10048 3188
rect 10003 3148 10048 3176
rect 7837 3139 7895 3145
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 11241 3179 11299 3185
rect 11241 3145 11253 3179
rect 11287 3176 11299 3179
rect 12986 3176 12992 3188
rect 11287 3148 12992 3176
rect 11287 3145 11299 3148
rect 11241 3139 11299 3145
rect 6638 3068 6644 3120
rect 6696 3108 6702 3120
rect 10060 3108 10088 3136
rect 6696 3080 10088 3108
rect 6696 3068 6702 3080
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6564 3012 6929 3040
rect 4801 3003 4859 3009
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 5442 2932 5448 2984
rect 5500 2972 5506 2984
rect 6638 2972 6644 2984
rect 5500 2944 6644 2972
rect 5500 2932 5506 2944
rect 6638 2932 6644 2944
rect 6696 2932 6702 2984
rect 10597 2975 10655 2981
rect 10597 2941 10609 2975
rect 10643 2972 10655 2975
rect 11256 2972 11284 3139
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 14507 3179 14565 3185
rect 14507 3145 14519 3179
rect 14553 3176 14565 3179
rect 15378 3176 15384 3188
rect 14553 3148 15384 3176
rect 14553 3145 14565 3148
rect 14507 3139 14565 3145
rect 15378 3136 15384 3148
rect 15436 3176 15442 3188
rect 15841 3179 15899 3185
rect 15841 3176 15853 3179
rect 15436 3148 15853 3176
rect 15436 3136 15442 3148
rect 15841 3145 15853 3148
rect 15887 3145 15899 3179
rect 15841 3139 15899 3145
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 17000 3148 17509 3176
rect 17000 3136 17006 3148
rect 17497 3145 17509 3148
rect 17543 3176 17555 3179
rect 17543 3148 19840 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 11517 3111 11575 3117
rect 11517 3108 11529 3111
rect 11388 3080 11529 3108
rect 11388 3068 11394 3080
rect 11517 3077 11529 3080
rect 11563 3077 11575 3111
rect 14918 3108 14924 3120
rect 14879 3080 14924 3108
rect 11517 3071 11575 3077
rect 14918 3068 14924 3080
rect 14976 3068 14982 3120
rect 15289 3111 15347 3117
rect 15289 3077 15301 3111
rect 15335 3108 15347 3111
rect 17218 3108 17224 3120
rect 15335 3080 17224 3108
rect 15335 3077 15347 3080
rect 15289 3071 15347 3077
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3040 12587 3043
rect 12618 3040 12624 3052
rect 12575 3012 12624 3040
rect 12575 3009 12587 3012
rect 12529 3003 12587 3009
rect 12618 3000 12624 3012
rect 12676 3000 12682 3052
rect 13170 3040 13176 3052
rect 13131 3012 13176 3040
rect 13170 3000 13176 3012
rect 13228 3040 13234 3052
rect 15463 3040 15491 3080
rect 17218 3068 17224 3080
rect 17276 3068 17282 3120
rect 19610 3068 19616 3120
rect 19668 3108 19674 3120
rect 19668 3080 19748 3108
rect 19668 3068 19674 3080
rect 16850 3040 16856 3052
rect 13228 3012 15491 3040
rect 16811 3012 16856 3040
rect 13228 3000 13234 3012
rect 10643 2944 11284 2972
rect 14436 2975 14494 2981
rect 10643 2941 10655 2944
rect 10597 2935 10655 2941
rect 14436 2941 14448 2975
rect 14482 2972 14494 2975
rect 14918 2972 14924 2984
rect 14482 2944 14924 2972
rect 14482 2941 14494 2944
rect 14436 2935 14494 2941
rect 14918 2932 14924 2944
rect 14976 2932 14982 2984
rect 15463 2981 15491 3012
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3040 17923 3043
rect 18141 3043 18199 3049
rect 18141 3040 18153 3043
rect 17911 3012 18153 3040
rect 17911 3009 17923 3012
rect 17865 3003 17923 3009
rect 18141 3009 18153 3012
rect 18187 3040 18199 3043
rect 18414 3040 18420 3052
rect 18187 3012 18420 3040
rect 18187 3009 18199 3012
rect 18141 3003 18199 3009
rect 18414 3000 18420 3012
rect 18472 3000 18478 3052
rect 19720 3049 19748 3080
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3009 19763 3043
rect 19812 3040 19840 3148
rect 19981 3043 20039 3049
rect 19981 3040 19993 3043
rect 19812 3012 19993 3040
rect 19705 3003 19763 3009
rect 19981 3009 19993 3012
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 15448 2975 15506 2981
rect 15448 2941 15460 2975
rect 15494 2941 15506 2975
rect 15448 2935 15506 2941
rect 7561 2907 7619 2913
rect 4126 2876 5396 2904
rect 3878 2836 3884 2848
rect 3839 2808 3884 2836
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 4525 2839 4583 2845
rect 4525 2805 4537 2839
rect 4571 2836 4583 2839
rect 4614 2836 4620 2848
rect 4571 2808 4620 2836
rect 4571 2805 4583 2808
rect 4525 2799 4583 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 5368 2836 5396 2876
rect 7561 2873 7573 2907
rect 7607 2873 7619 2907
rect 7561 2867 7619 2873
rect 9125 2907 9183 2913
rect 9125 2873 9137 2907
rect 9171 2873 9183 2907
rect 9125 2867 9183 2873
rect 9769 2907 9827 2913
rect 9769 2873 9781 2907
rect 9815 2904 9827 2907
rect 10134 2904 10140 2916
rect 9815 2876 10140 2904
rect 9815 2873 9827 2876
rect 9769 2867 9827 2873
rect 7576 2836 7604 2867
rect 8202 2836 8208 2848
rect 5368 2808 8208 2836
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 8849 2839 8907 2845
rect 8849 2836 8861 2839
rect 8444 2808 8861 2836
rect 8444 2796 8450 2808
rect 8849 2805 8861 2808
rect 8895 2836 8907 2839
rect 9140 2836 9168 2867
rect 10134 2864 10140 2876
rect 10192 2864 10198 2916
rect 10226 2864 10232 2916
rect 10284 2904 10290 2916
rect 11974 2904 11980 2916
rect 10284 2876 11980 2904
rect 10284 2864 10290 2876
rect 11974 2864 11980 2876
rect 12032 2904 12038 2916
rect 12161 2907 12219 2913
rect 12161 2904 12173 2907
rect 12032 2876 12173 2904
rect 12032 2864 12038 2876
rect 12161 2873 12173 2876
rect 12207 2904 12219 2907
rect 13446 2904 13452 2916
rect 12207 2876 13452 2904
rect 12207 2873 12219 2876
rect 12161 2867 12219 2873
rect 13446 2864 13452 2876
rect 13504 2864 13510 2916
rect 16301 2907 16359 2913
rect 16301 2873 16313 2907
rect 16347 2904 16359 2907
rect 16485 2907 16543 2913
rect 16485 2904 16497 2907
rect 16347 2876 16497 2904
rect 16347 2873 16359 2876
rect 16301 2867 16359 2873
rect 16485 2873 16497 2876
rect 16531 2904 16543 2907
rect 18782 2904 18788 2916
rect 16531 2876 18788 2904
rect 16531 2873 16543 2876
rect 16485 2867 16543 2873
rect 18782 2864 18788 2876
rect 18840 2864 18846 2916
rect 8895 2808 9168 2836
rect 10781 2839 10839 2845
rect 8895 2805 8907 2808
rect 8849 2799 8907 2805
rect 10781 2805 10793 2839
rect 10827 2836 10839 2839
rect 10962 2836 10968 2848
rect 10827 2808 10968 2836
rect 10827 2805 10839 2808
rect 10781 2799 10839 2805
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 15519 2839 15577 2845
rect 15519 2805 15531 2839
rect 15565 2836 15577 2839
rect 17310 2836 17316 2848
rect 15565 2808 17316 2836
rect 15565 2805 15577 2808
rect 15519 2799 15577 2805
rect 17310 2796 17316 2808
rect 17368 2796 17374 2848
rect 19518 2836 19524 2848
rect 19431 2808 19524 2836
rect 19518 2796 19524 2808
rect 19576 2836 19582 2848
rect 21726 2836 21732 2848
rect 19576 2808 21732 2836
rect 19576 2796 19582 2808
rect 21726 2796 21732 2808
rect 21784 2796 21790 2848
rect 1104 2746 21436 2768
rect 1104 2694 8497 2746
rect 8549 2694 8561 2746
rect 8613 2694 8625 2746
rect 8677 2694 8689 2746
rect 8741 2694 16012 2746
rect 16064 2694 16076 2746
rect 16128 2694 16140 2746
rect 16192 2694 16204 2746
rect 16256 2694 21436 2746
rect 1104 2672 21436 2694
rect 2087 2635 2145 2641
rect 2087 2601 2099 2635
rect 2133 2632 2145 2635
rect 8386 2632 8392 2644
rect 2133 2604 8392 2632
rect 2133 2601 2145 2604
rect 2087 2595 2145 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 9398 2632 9404 2644
rect 9311 2604 9404 2632
rect 9398 2592 9404 2604
rect 9456 2632 9462 2644
rect 11977 2635 12035 2641
rect 11977 2632 11989 2635
rect 9456 2604 11989 2632
rect 9456 2592 9462 2604
rect 3237 2567 3295 2573
rect 3237 2533 3249 2567
rect 3283 2564 3295 2567
rect 7377 2567 7435 2573
rect 3283 2536 7328 2564
rect 3283 2533 3295 2536
rect 3237 2527 3295 2533
rect 2016 2499 2074 2505
rect 2016 2465 2028 2499
rect 2062 2496 2074 2499
rect 2498 2496 2504 2508
rect 2062 2468 2504 2496
rect 2062 2465 2074 2468
rect 2016 2459 2074 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 3028 2499 3086 2505
rect 3028 2465 3040 2499
rect 3074 2496 3086 2499
rect 3421 2499 3479 2505
rect 3421 2496 3433 2499
rect 3074 2468 3433 2496
rect 3074 2465 3086 2468
rect 3028 2459 3086 2465
rect 3421 2465 3433 2468
rect 3467 2465 3479 2499
rect 3421 2459 3479 2465
rect 4316 2499 4374 2505
rect 4316 2465 4328 2499
rect 4362 2496 4374 2499
rect 4614 2496 4620 2508
rect 4362 2468 4620 2496
rect 4362 2465 4374 2468
rect 4316 2459 4374 2465
rect 3436 2428 3464 2459
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6052 2468 6097 2496
rect 6052 2456 6058 2468
rect 4985 2431 5043 2437
rect 4985 2428 4997 2431
rect 3436 2400 4997 2428
rect 4985 2397 4997 2400
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2397 5411 2431
rect 7300 2428 7328 2536
rect 7377 2533 7389 2567
rect 7423 2564 7435 2567
rect 7561 2567 7619 2573
rect 7561 2564 7573 2567
rect 7423 2536 7573 2564
rect 7423 2533 7435 2536
rect 7377 2527 7435 2533
rect 7561 2533 7573 2536
rect 7607 2564 7619 2567
rect 10134 2564 10140 2576
rect 7607 2536 10140 2564
rect 7607 2533 7619 2536
rect 7561 2527 7619 2533
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 11440 2505 11468 2604
rect 11977 2601 11989 2604
rect 12023 2632 12035 2635
rect 12161 2635 12219 2641
rect 12161 2632 12173 2635
rect 12023 2604 12173 2632
rect 12023 2601 12035 2604
rect 11977 2595 12035 2601
rect 12161 2601 12173 2604
rect 12207 2601 12219 2635
rect 12161 2595 12219 2601
rect 12618 2592 12624 2644
rect 12676 2632 12682 2644
rect 16117 2635 16175 2641
rect 12676 2604 13400 2632
rect 12676 2592 12682 2604
rect 13372 2573 13400 2604
rect 16117 2601 16129 2635
rect 16163 2632 16175 2635
rect 16298 2632 16304 2644
rect 16163 2604 16304 2632
rect 16163 2601 16175 2604
rect 16117 2595 16175 2601
rect 13357 2567 13415 2573
rect 13357 2533 13369 2567
rect 13403 2533 13415 2567
rect 13357 2527 13415 2533
rect 13446 2524 13452 2576
rect 13504 2564 13510 2576
rect 13504 2536 13814 2564
rect 13504 2524 13510 2536
rect 11425 2499 11483 2505
rect 8260 2468 8305 2496
rect 8260 2456 8266 2468
rect 11425 2465 11437 2499
rect 11471 2465 11483 2499
rect 13786 2496 13814 2536
rect 14236 2499 14294 2505
rect 14236 2496 14248 2499
rect 13786 2468 14248 2496
rect 11425 2459 11483 2465
rect 14236 2465 14248 2468
rect 14282 2496 14294 2499
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 14282 2468 14657 2496
rect 14282 2465 14294 2468
rect 14236 2459 14294 2465
rect 14645 2465 14657 2468
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 16132 2496 16160 2595
rect 16298 2592 16304 2604
rect 16356 2592 16362 2644
rect 17310 2592 17316 2644
rect 17368 2632 17374 2644
rect 19610 2632 19616 2644
rect 17368 2604 19104 2632
rect 19571 2604 19616 2632
rect 17368 2592 17374 2604
rect 18141 2567 18199 2573
rect 18141 2533 18153 2567
rect 18187 2564 18199 2567
rect 18417 2567 18475 2573
rect 18417 2564 18429 2567
rect 18187 2536 18429 2564
rect 18187 2533 18199 2536
rect 18141 2527 18199 2533
rect 18417 2533 18429 2536
rect 18463 2564 18475 2567
rect 18506 2564 18512 2576
rect 18463 2536 18512 2564
rect 18463 2533 18475 2536
rect 18417 2527 18475 2533
rect 18506 2524 18512 2536
rect 18564 2524 18570 2576
rect 15519 2468 16160 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 16482 2456 16488 2508
rect 16540 2496 16546 2508
rect 16577 2499 16635 2505
rect 16577 2496 16589 2499
rect 16540 2468 16589 2496
rect 16540 2456 16546 2468
rect 16577 2465 16589 2468
rect 16623 2496 16635 2499
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 16623 2468 17141 2496
rect 16623 2465 16635 2468
rect 16577 2459 16635 2465
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 19076 2496 19104 2604
rect 19610 2592 19616 2604
rect 19668 2592 19674 2644
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19076 2468 19901 2496
rect 17129 2459 17187 2465
rect 19889 2465 19901 2468
rect 19935 2496 19947 2499
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 19935 2468 20453 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 20441 2459 20499 2465
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 7300 2400 9505 2428
rect 5353 2391 5411 2397
rect 9493 2397 9505 2400
rect 9539 2428 9551 2431
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9539 2400 9873 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 10134 2428 10140 2440
rect 10095 2400 10140 2428
rect 9861 2391 9919 2397
rect 4387 2363 4445 2369
rect 4387 2329 4399 2363
rect 4433 2360 4445 2363
rect 5077 2363 5135 2369
rect 5077 2360 5089 2363
rect 4433 2332 5089 2360
rect 4433 2329 4445 2332
rect 4387 2323 4445 2329
rect 5077 2329 5089 2332
rect 5123 2360 5135 2363
rect 5368 2360 5396 2391
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12483 2400 12725 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 12713 2397 12725 2400
rect 12759 2428 12771 2431
rect 14323 2431 14381 2437
rect 14323 2428 14335 2431
rect 12759 2400 14335 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 14323 2397 14335 2400
rect 14369 2397 14381 2431
rect 18782 2428 18788 2440
rect 18743 2400 18788 2428
rect 14323 2391 14381 2397
rect 18782 2388 18788 2400
rect 18840 2388 18846 2440
rect 5123 2332 5396 2360
rect 11609 2363 11667 2369
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 13170 2360 13176 2372
rect 11655 2332 13176 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 13170 2320 13176 2332
rect 13228 2320 13234 2372
rect 16761 2363 16819 2369
rect 16761 2329 16773 2363
rect 16807 2360 16819 2363
rect 17310 2360 17316 2372
rect 16807 2332 17316 2360
rect 16807 2329 16819 2332
rect 16761 2323 16819 2329
rect 17310 2320 17316 2332
rect 17368 2320 17374 2372
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 4614 2252 4620 2304
rect 4672 2292 4678 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4672 2264 4721 2292
rect 4672 2252 4678 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 4985 2295 5043 2301
rect 4985 2261 4997 2295
rect 5031 2292 5043 2295
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 5031 2264 9413 2292
rect 5031 2261 5043 2264
rect 4985 2255 5043 2261
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 9401 2255 9459 2261
rect 12161 2295 12219 2301
rect 12161 2261 12173 2295
rect 12207 2292 12219 2295
rect 13814 2292 13820 2304
rect 12207 2264 13820 2292
rect 12207 2261 12219 2264
rect 12161 2255 12219 2261
rect 13814 2252 13820 2264
rect 13872 2252 13878 2304
rect 14274 2252 14280 2304
rect 14332 2292 14338 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 14332 2264 15669 2292
rect 14332 2252 14338 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 19426 2252 19432 2304
rect 19484 2292 19490 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 19484 2264 20085 2292
rect 19484 2252 19490 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 1104 2202 21436 2224
rect 1104 2150 4739 2202
rect 4791 2150 4803 2202
rect 4855 2150 4867 2202
rect 4919 2150 4931 2202
rect 4983 2150 12255 2202
rect 12307 2150 12319 2202
rect 12371 2150 12383 2202
rect 12435 2150 12447 2202
rect 12499 2150 19770 2202
rect 19822 2150 19834 2202
rect 19886 2150 19898 2202
rect 19950 2150 19962 2202
rect 20014 2150 21436 2202
rect 1104 2128 21436 2150
rect 12802 76 12808 128
rect 12860 116 12866 128
rect 18414 116 18420 128
rect 12860 88 18420 116
rect 12860 76 12866 88
rect 18414 76 18420 88
rect 18472 76 18478 128
rect 20714 76 20720 128
rect 20772 116 20778 128
rect 21358 116 21364 128
rect 20772 88 21364 116
rect 20772 76 20778 88
rect 21358 76 21364 88
rect 21416 76 21422 128
<< via1 >>
rect 2780 24216 2832 24268
rect 4068 24216 4120 24268
rect 5264 24216 5316 24268
rect 7840 24216 7892 24268
rect 8497 22278 8549 22330
rect 8561 22278 8613 22330
rect 8625 22278 8677 22330
rect 8689 22278 8741 22330
rect 16012 22278 16064 22330
rect 16076 22278 16128 22330
rect 16140 22278 16192 22330
rect 16204 22278 16256 22330
rect 20 22040 72 22092
rect 15568 22040 15620 22092
rect 20168 22040 20220 22092
rect 112 21972 164 22024
rect 12992 21972 13044 22024
rect 19616 21836 19668 21888
rect 4739 21734 4791 21786
rect 4803 21734 4855 21786
rect 4867 21734 4919 21786
rect 4931 21734 4983 21786
rect 12255 21734 12307 21786
rect 12319 21734 12371 21786
rect 12383 21734 12435 21786
rect 12447 21734 12499 21786
rect 19770 21734 19822 21786
rect 19834 21734 19886 21786
rect 19898 21734 19950 21786
rect 19962 21734 20014 21786
rect 10324 21496 10376 21548
rect 10968 21496 11020 21548
rect 15568 21428 15620 21480
rect 15016 21403 15068 21412
rect 14096 21335 14148 21344
rect 14096 21301 14105 21335
rect 14105 21301 14139 21335
rect 14139 21301 14148 21335
rect 15016 21369 15025 21403
rect 15025 21369 15059 21403
rect 15059 21369 15068 21403
rect 15016 21360 15068 21369
rect 18420 21632 18472 21684
rect 20168 21632 20220 21684
rect 20260 21564 20312 21616
rect 21548 21632 21600 21684
rect 14096 21292 14148 21301
rect 16304 21292 16356 21344
rect 16396 21292 16448 21344
rect 19708 21292 19760 21344
rect 8497 21190 8549 21242
rect 8561 21190 8613 21242
rect 8625 21190 8677 21242
rect 8689 21190 8741 21242
rect 16012 21190 16064 21242
rect 16076 21190 16128 21242
rect 16140 21190 16192 21242
rect 16204 21190 16256 21242
rect 8944 21088 8996 21140
rect 12072 21088 12124 21140
rect 1584 20952 1636 21004
rect 9588 20995 9640 21004
rect 9588 20961 9597 20995
rect 9597 20961 9631 20995
rect 9631 20961 9640 20995
rect 9588 20952 9640 20961
rect 12072 20952 12124 21004
rect 14832 21020 14884 21072
rect 16396 21020 16448 21072
rect 19340 21063 19392 21072
rect 19340 21029 19349 21063
rect 19349 21029 19383 21063
rect 19383 21029 19392 21063
rect 19340 21020 19392 21029
rect 19708 21020 19760 21072
rect 12992 20952 13044 21004
rect 18512 20952 18564 21004
rect 8576 20884 8628 20936
rect 16580 20927 16632 20936
rect 16580 20893 16589 20927
rect 16589 20893 16623 20927
rect 16623 20893 16632 20927
rect 16580 20884 16632 20893
rect 20076 20884 20128 20936
rect 1952 20748 2004 20800
rect 13912 20748 13964 20800
rect 19524 20748 19576 20800
rect 4739 20646 4791 20698
rect 4803 20646 4855 20698
rect 4867 20646 4919 20698
rect 4931 20646 4983 20698
rect 12255 20646 12307 20698
rect 12319 20646 12371 20698
rect 12383 20646 12435 20698
rect 12447 20646 12499 20698
rect 19770 20646 19822 20698
rect 19834 20646 19886 20698
rect 19898 20646 19950 20698
rect 19962 20646 20014 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 1952 20587 2004 20596
rect 1952 20553 1961 20587
rect 1961 20553 1995 20587
rect 1995 20553 2004 20587
rect 1952 20544 2004 20553
rect 8576 20587 8628 20596
rect 8576 20553 8585 20587
rect 8585 20553 8619 20587
rect 8619 20553 8628 20587
rect 8576 20544 8628 20553
rect 12992 20544 13044 20596
rect 13912 20587 13964 20596
rect 13912 20553 13921 20587
rect 13921 20553 13955 20587
rect 13955 20553 13964 20587
rect 13912 20544 13964 20553
rect 16396 20544 16448 20596
rect 18512 20544 18564 20596
rect 19340 20587 19392 20596
rect 19340 20553 19349 20587
rect 19349 20553 19383 20587
rect 19383 20553 19392 20587
rect 19340 20544 19392 20553
rect 17040 20476 17092 20528
rect 16580 20408 16632 20460
rect 19616 20451 19668 20460
rect 19616 20417 19625 20451
rect 19625 20417 19659 20451
rect 19659 20417 19668 20451
rect 19616 20408 19668 20417
rect 2872 20315 2924 20324
rect 2872 20281 2881 20315
rect 2881 20281 2915 20315
rect 2915 20281 2924 20315
rect 2872 20272 2924 20281
rect 9588 20272 9640 20324
rect 12072 20204 12124 20256
rect 15016 20204 15068 20256
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 8497 20102 8549 20154
rect 8561 20102 8613 20154
rect 8625 20102 8677 20154
rect 8689 20102 8741 20154
rect 16012 20102 16064 20154
rect 16076 20102 16128 20154
rect 16140 20102 16192 20154
rect 16204 20102 16256 20154
rect 14096 20043 14148 20052
rect 14096 20009 14105 20043
rect 14105 20009 14139 20043
rect 14139 20009 14148 20043
rect 14096 20000 14148 20009
rect 15016 19932 15068 19984
rect 16304 19932 16356 19984
rect 16948 19975 17000 19984
rect 16948 19941 16957 19975
rect 16957 19941 16991 19975
rect 16991 19941 17000 19975
rect 16948 19932 17000 19941
rect 17868 19932 17920 19984
rect 20076 19932 20128 19984
rect 15844 19796 15896 19848
rect 16580 19796 16632 19848
rect 19340 19839 19392 19848
rect 19340 19805 19349 19839
rect 19349 19805 19383 19839
rect 19383 19805 19392 19839
rect 19340 19796 19392 19805
rect 4739 19558 4791 19610
rect 4803 19558 4855 19610
rect 4867 19558 4919 19610
rect 4931 19558 4983 19610
rect 12255 19558 12307 19610
rect 12319 19558 12371 19610
rect 12383 19558 12435 19610
rect 12447 19558 12499 19610
rect 19770 19558 19822 19610
rect 19834 19558 19886 19610
rect 19898 19558 19950 19610
rect 19962 19558 20014 19610
rect 15476 19456 15528 19508
rect 15844 19499 15896 19508
rect 15844 19465 15853 19499
rect 15853 19465 15887 19499
rect 15887 19465 15896 19499
rect 15844 19456 15896 19465
rect 16948 19499 17000 19508
rect 16948 19465 16957 19499
rect 16957 19465 16991 19499
rect 16991 19465 17000 19499
rect 16948 19456 17000 19465
rect 17868 19499 17920 19508
rect 17868 19465 17877 19499
rect 17877 19465 17911 19499
rect 17911 19465 17920 19499
rect 17868 19456 17920 19465
rect 15016 19295 15068 19304
rect 15016 19261 15034 19295
rect 15034 19261 15068 19295
rect 15660 19320 15712 19372
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 19524 19320 19576 19372
rect 15016 19252 15068 19261
rect 19432 19184 19484 19236
rect 19340 19159 19392 19168
rect 19340 19125 19349 19159
rect 19349 19125 19383 19159
rect 19383 19125 19392 19159
rect 19340 19116 19392 19125
rect 8497 19014 8549 19066
rect 8561 19014 8613 19066
rect 8625 19014 8677 19066
rect 8689 19014 8741 19066
rect 16012 19014 16064 19066
rect 16076 19014 16128 19066
rect 16140 19014 16192 19066
rect 16204 19014 16256 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 19340 18912 19392 18964
rect 19524 18844 19576 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 6644 18776 6696 18828
rect 20352 18776 20404 18828
rect 6092 18572 6144 18624
rect 4739 18470 4791 18522
rect 4803 18470 4855 18522
rect 4867 18470 4919 18522
rect 4931 18470 4983 18522
rect 12255 18470 12307 18522
rect 12319 18470 12371 18522
rect 12383 18470 12435 18522
rect 12447 18470 12499 18522
rect 19770 18470 19822 18522
rect 19834 18470 19886 18522
rect 19898 18470 19950 18522
rect 19962 18470 20014 18522
rect 1400 18368 1452 18420
rect 7472 18411 7524 18420
rect 7472 18377 7481 18411
rect 7481 18377 7515 18411
rect 7515 18377 7524 18411
rect 7472 18368 7524 18377
rect 20352 18368 20404 18420
rect 6644 18275 6696 18284
rect 6644 18241 6653 18275
rect 6653 18241 6687 18275
rect 6687 18241 6696 18275
rect 6644 18232 6696 18241
rect 11704 18232 11756 18284
rect 7104 18164 7156 18216
rect 8852 18028 8904 18080
rect 9496 18028 9548 18080
rect 8497 17926 8549 17978
rect 8561 17926 8613 17978
rect 8625 17926 8677 17978
rect 8689 17926 8741 17978
rect 16012 17926 16064 17978
rect 16076 17926 16128 17978
rect 16140 17926 16192 17978
rect 16204 17926 16256 17978
rect 1400 17824 1452 17876
rect 6276 17867 6328 17876
rect 6276 17833 6285 17867
rect 6285 17833 6319 17867
rect 6319 17833 6328 17867
rect 6276 17824 6328 17833
rect 1768 17688 1820 17740
rect 6092 17731 6144 17740
rect 6092 17697 6101 17731
rect 6101 17697 6135 17731
rect 6135 17697 6144 17731
rect 6092 17688 6144 17697
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 4739 17382 4791 17434
rect 4803 17382 4855 17434
rect 4867 17382 4919 17434
rect 4931 17382 4983 17434
rect 12255 17382 12307 17434
rect 12319 17382 12371 17434
rect 12383 17382 12435 17434
rect 12447 17382 12499 17434
rect 19770 17382 19822 17434
rect 19834 17382 19886 17434
rect 19898 17382 19950 17434
rect 19962 17382 20014 17434
rect 2872 17280 2924 17332
rect 6092 17323 6144 17332
rect 6092 17289 6101 17323
rect 6101 17289 6135 17323
rect 6135 17289 6144 17323
rect 6092 17280 6144 17289
rect 7104 17323 7156 17332
rect 7104 17289 7113 17323
rect 7113 17289 7147 17323
rect 7147 17289 7156 17323
rect 7104 17280 7156 17289
rect 7656 17323 7708 17332
rect 7656 17289 7665 17323
rect 7665 17289 7699 17323
rect 7699 17289 7708 17323
rect 7656 17280 7708 17289
rect 7748 17144 7800 17196
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 1768 16983 1820 16992
rect 1768 16949 1777 16983
rect 1777 16949 1811 16983
rect 1811 16949 1820 16983
rect 1768 16940 1820 16949
rect 2688 16940 2740 16992
rect 8392 16940 8444 16992
rect 8497 16838 8549 16890
rect 8561 16838 8613 16890
rect 8625 16838 8677 16890
rect 8689 16838 8741 16890
rect 16012 16838 16064 16890
rect 16076 16838 16128 16890
rect 16140 16838 16192 16890
rect 16204 16838 16256 16890
rect 19248 16736 19300 16788
rect 19800 16779 19852 16788
rect 19800 16745 19809 16779
rect 19809 16745 19843 16779
rect 19843 16745 19852 16779
rect 19800 16736 19852 16745
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 19432 16600 19484 16652
rect 8116 16575 8168 16584
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 8392 16575 8444 16584
rect 8392 16541 8401 16575
rect 8401 16541 8435 16575
rect 8435 16541 8444 16575
rect 8392 16532 8444 16541
rect 4739 16294 4791 16346
rect 4803 16294 4855 16346
rect 4867 16294 4919 16346
rect 4931 16294 4983 16346
rect 12255 16294 12307 16346
rect 12319 16294 12371 16346
rect 12383 16294 12435 16346
rect 12447 16294 12499 16346
rect 19770 16294 19822 16346
rect 19834 16294 19886 16346
rect 19898 16294 19950 16346
rect 19962 16294 20014 16346
rect 19524 16056 19576 16108
rect 8024 15963 8076 15972
rect 8024 15929 8033 15963
rect 8033 15929 8067 15963
rect 8067 15929 8076 15963
rect 8024 15920 8076 15929
rect 8116 15852 8168 15904
rect 9128 15920 9180 15972
rect 19524 15920 19576 15972
rect 9680 15895 9732 15904
rect 9680 15861 9689 15895
rect 9689 15861 9723 15895
rect 9723 15861 9732 15895
rect 9680 15852 9732 15861
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 8497 15750 8549 15802
rect 8561 15750 8613 15802
rect 8625 15750 8677 15802
rect 8689 15750 8741 15802
rect 16012 15750 16064 15802
rect 16076 15750 16128 15802
rect 16140 15750 16192 15802
rect 16204 15750 16256 15802
rect 8024 15648 8076 15700
rect 19524 15580 19576 15632
rect 7380 15512 7432 15564
rect 9680 15512 9732 15564
rect 20076 15512 20128 15564
rect 4739 15206 4791 15258
rect 4803 15206 4855 15258
rect 4867 15206 4919 15258
rect 4931 15206 4983 15258
rect 12255 15206 12307 15258
rect 12319 15206 12371 15258
rect 12383 15206 12435 15258
rect 12447 15206 12499 15258
rect 19770 15206 19822 15258
rect 19834 15206 19886 15258
rect 19898 15206 19950 15258
rect 19962 15206 20014 15258
rect 14556 15147 14608 15156
rect 14556 15113 14565 15147
rect 14565 15113 14599 15147
rect 14599 15113 14608 15147
rect 14556 15104 14608 15113
rect 15016 15147 15068 15156
rect 15016 15113 15025 15147
rect 15025 15113 15059 15147
rect 15059 15113 15068 15147
rect 15016 15104 15068 15113
rect 9128 15011 9180 15020
rect 9128 14977 9137 15011
rect 9137 14977 9171 15011
rect 9171 14977 9180 15011
rect 9128 14968 9180 14977
rect 19432 15104 19484 15156
rect 20260 14943 20312 14952
rect 20260 14909 20269 14943
rect 20269 14909 20303 14943
rect 20303 14909 20312 14943
rect 20260 14900 20312 14909
rect 8852 14875 8904 14884
rect 8852 14841 8861 14875
rect 8861 14841 8895 14875
rect 8895 14841 8904 14875
rect 8852 14832 8904 14841
rect 20076 14832 20128 14884
rect 20720 14832 20772 14884
rect 7380 14764 7432 14816
rect 15844 14764 15896 14816
rect 8497 14662 8549 14714
rect 8561 14662 8613 14714
rect 8625 14662 8677 14714
rect 8689 14662 8741 14714
rect 16012 14662 16064 14714
rect 16076 14662 16128 14714
rect 16140 14662 16192 14714
rect 16204 14662 16256 14714
rect 8852 14560 8904 14612
rect 13452 14560 13504 14612
rect 15844 14492 15896 14544
rect 9772 14424 9824 14476
rect 13636 14467 13688 14476
rect 13636 14433 13645 14467
rect 13645 14433 13679 14467
rect 13679 14433 13688 14467
rect 13636 14424 13688 14433
rect 16672 14331 16724 14340
rect 16672 14297 16681 14331
rect 16681 14297 16715 14331
rect 16715 14297 16724 14331
rect 16672 14288 16724 14297
rect 4739 14118 4791 14170
rect 4803 14118 4855 14170
rect 4867 14118 4919 14170
rect 4931 14118 4983 14170
rect 12255 14118 12307 14170
rect 12319 14118 12371 14170
rect 12383 14118 12435 14170
rect 12447 14118 12499 14170
rect 19770 14118 19822 14170
rect 19834 14118 19886 14170
rect 19898 14118 19950 14170
rect 19962 14118 20014 14170
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 10876 14016 10928 14068
rect 13636 14059 13688 14068
rect 13636 14025 13645 14059
rect 13645 14025 13679 14059
rect 13679 14025 13688 14059
rect 13636 14016 13688 14025
rect 15844 14016 15896 14068
rect 18236 13948 18288 14000
rect 16672 13923 16724 13932
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 16672 13880 16724 13889
rect 19156 13880 19208 13932
rect 20260 13948 20312 14000
rect 16304 13744 16356 13796
rect 19156 13744 19208 13796
rect 19432 13744 19484 13796
rect 10048 13676 10100 13728
rect 8497 13574 8549 13626
rect 8561 13574 8613 13626
rect 8625 13574 8677 13626
rect 8689 13574 8741 13626
rect 16012 13574 16064 13626
rect 16076 13574 16128 13626
rect 16140 13574 16192 13626
rect 16204 13574 16256 13626
rect 16304 13472 16356 13524
rect 13636 13336 13688 13388
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 10048 13311 10100 13320
rect 10048 13277 10057 13311
rect 10057 13277 10091 13311
rect 10091 13277 10100 13311
rect 10048 13268 10100 13277
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 4739 13030 4791 13082
rect 4803 13030 4855 13082
rect 4867 13030 4919 13082
rect 4931 13030 4983 13082
rect 12255 13030 12307 13082
rect 12319 13030 12371 13082
rect 12383 13030 12435 13082
rect 12447 13030 12499 13082
rect 19770 13030 19822 13082
rect 19834 13030 19886 13082
rect 19898 13030 19950 13082
rect 19962 13030 20014 13082
rect 10048 12928 10100 12980
rect 10416 12903 10468 12912
rect 10416 12869 10425 12903
rect 10425 12869 10459 12903
rect 10459 12869 10468 12903
rect 10416 12860 10468 12869
rect 19432 12792 19484 12844
rect 9864 12699 9916 12708
rect 9864 12665 9873 12699
rect 9873 12665 9907 12699
rect 9907 12665 9916 12699
rect 9864 12656 9916 12665
rect 19432 12699 19484 12708
rect 19432 12665 19441 12699
rect 19441 12665 19475 12699
rect 19475 12665 19484 12699
rect 19432 12656 19484 12665
rect 15660 12631 15712 12640
rect 15660 12597 15669 12631
rect 15669 12597 15703 12631
rect 15703 12597 15712 12631
rect 15660 12588 15712 12597
rect 8497 12486 8549 12538
rect 8561 12486 8613 12538
rect 8625 12486 8677 12538
rect 8689 12486 8741 12538
rect 16012 12486 16064 12538
rect 16076 12486 16128 12538
rect 16140 12486 16192 12538
rect 16204 12486 16256 12538
rect 19432 12384 19484 12436
rect 9772 12359 9824 12368
rect 9772 12325 9781 12359
rect 9781 12325 9815 12359
rect 9815 12325 9824 12359
rect 9772 12316 9824 12325
rect 10416 12316 10468 12368
rect 19616 12291 19668 12300
rect 19616 12257 19625 12291
rect 19625 12257 19659 12291
rect 19659 12257 19668 12291
rect 19616 12248 19668 12257
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 9404 12180 9456 12232
rect 4739 11942 4791 11994
rect 4803 11942 4855 11994
rect 4867 11942 4919 11994
rect 4931 11942 4983 11994
rect 12255 11942 12307 11994
rect 12319 11942 12371 11994
rect 12383 11942 12435 11994
rect 12447 11942 12499 11994
rect 19770 11942 19822 11994
rect 19834 11942 19886 11994
rect 19898 11942 19950 11994
rect 19962 11942 20014 11994
rect 8484 11883 8536 11892
rect 8484 11849 8493 11883
rect 8493 11849 8527 11883
rect 8527 11849 8536 11883
rect 8484 11840 8536 11849
rect 9772 11883 9824 11892
rect 9772 11849 9781 11883
rect 9781 11849 9815 11883
rect 9815 11849 9824 11883
rect 9772 11840 9824 11849
rect 9864 11840 9916 11892
rect 12624 11883 12676 11892
rect 12624 11849 12633 11883
rect 12633 11849 12667 11883
rect 12667 11849 12676 11883
rect 12624 11840 12676 11849
rect 9404 11747 9456 11756
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 12624 11636 12676 11688
rect 15292 11636 15344 11688
rect 15660 11636 15712 11688
rect 16304 11636 16356 11688
rect 10876 11568 10928 11620
rect 7932 11500 7984 11552
rect 16396 11500 16448 11552
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 18696 11500 18748 11552
rect 19524 11500 19576 11552
rect 19616 11500 19668 11552
rect 20628 11500 20680 11552
rect 8497 11398 8549 11450
rect 8561 11398 8613 11450
rect 8625 11398 8677 11450
rect 8689 11398 8741 11450
rect 16012 11398 16064 11450
rect 16076 11398 16128 11450
rect 16140 11398 16192 11450
rect 16204 11398 16256 11450
rect 12624 11339 12676 11348
rect 12624 11305 12633 11339
rect 12633 11305 12667 11339
rect 12667 11305 12676 11339
rect 12624 11296 12676 11305
rect 19800 11339 19852 11348
rect 19800 11305 19809 11339
rect 19809 11305 19843 11339
rect 19843 11305 19852 11339
rect 19800 11296 19852 11305
rect 16396 11271 16448 11280
rect 16396 11237 16405 11271
rect 16405 11237 16439 11271
rect 16439 11237 16448 11271
rect 16396 11228 16448 11237
rect 7932 11203 7984 11212
rect 7932 11169 7941 11203
rect 7941 11169 7975 11203
rect 7975 11169 7984 11203
rect 7932 11160 7984 11169
rect 12900 11160 12952 11212
rect 19524 11160 19576 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 18788 11092 18840 11144
rect 8116 11067 8168 11076
rect 8116 11033 8125 11067
rect 8125 11033 8159 11067
rect 8159 11033 8168 11067
rect 8116 11024 8168 11033
rect 16948 11067 17000 11076
rect 16948 11033 16957 11067
rect 16957 11033 16991 11067
rect 16991 11033 17000 11067
rect 16948 11024 17000 11033
rect 4739 10854 4791 10906
rect 4803 10854 4855 10906
rect 4867 10854 4919 10906
rect 4931 10854 4983 10906
rect 12255 10854 12307 10906
rect 12319 10854 12371 10906
rect 12383 10854 12435 10906
rect 12447 10854 12499 10906
rect 19770 10854 19822 10906
rect 19834 10854 19886 10906
rect 19898 10854 19950 10906
rect 19962 10854 20014 10906
rect 7932 10752 7984 10804
rect 12900 10795 12952 10804
rect 12900 10761 12909 10795
rect 12909 10761 12943 10795
rect 12943 10761 12952 10795
rect 12900 10752 12952 10761
rect 16304 10795 16356 10804
rect 16304 10761 16313 10795
rect 16313 10761 16347 10795
rect 16347 10761 16356 10795
rect 16304 10752 16356 10761
rect 16396 10684 16448 10736
rect 7288 10616 7340 10668
rect 18052 10752 18104 10804
rect 16948 10659 17000 10668
rect 16948 10625 16957 10659
rect 16957 10625 16991 10659
rect 16991 10625 17000 10659
rect 19524 10752 19576 10804
rect 22100 10684 22152 10736
rect 16948 10616 17000 10625
rect 18788 10659 18840 10668
rect 18788 10625 18797 10659
rect 18797 10625 18831 10659
rect 18831 10625 18840 10659
rect 18788 10616 18840 10625
rect 112 10548 164 10600
rect 20076 10548 20128 10600
rect 1952 10480 2004 10532
rect 7472 10523 7524 10532
rect 7472 10489 7481 10523
rect 7481 10489 7515 10523
rect 7515 10489 7524 10523
rect 7472 10480 7524 10489
rect 1860 10412 1912 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 8497 10310 8549 10362
rect 8561 10310 8613 10362
rect 8625 10310 8677 10362
rect 8689 10310 8741 10362
rect 16012 10310 16064 10362
rect 16076 10310 16128 10362
rect 16140 10310 16192 10362
rect 16204 10310 16256 10362
rect 6184 10208 6236 10260
rect 7472 10208 7524 10260
rect 7288 10183 7340 10192
rect 7288 10149 7297 10183
rect 7297 10149 7331 10183
rect 7331 10149 7340 10183
rect 7288 10140 7340 10149
rect 12440 10140 12492 10192
rect 12808 10183 12860 10192
rect 12808 10149 12817 10183
rect 12817 10149 12851 10183
rect 12851 10149 12860 10183
rect 12808 10140 12860 10149
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 8116 10115 8168 10124
rect 8116 10081 8125 10115
rect 8125 10081 8159 10115
rect 8159 10081 8168 10115
rect 8116 10072 8168 10081
rect 10876 10072 10928 10124
rect 1952 10004 2004 10056
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 12900 10004 12952 10056
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 18696 10047 18748 10056
rect 18696 10013 18705 10047
rect 18705 10013 18739 10047
rect 18739 10013 18748 10047
rect 18696 10004 18748 10013
rect 2136 9979 2188 9988
rect 2136 9945 2145 9979
rect 2145 9945 2179 9979
rect 2179 9945 2188 9979
rect 2136 9936 2188 9945
rect 4739 9766 4791 9818
rect 4803 9766 4855 9818
rect 4867 9766 4919 9818
rect 4931 9766 4983 9818
rect 12255 9766 12307 9818
rect 12319 9766 12371 9818
rect 12383 9766 12435 9818
rect 12447 9766 12499 9818
rect 19770 9766 19822 9818
rect 19834 9766 19886 9818
rect 19898 9766 19950 9818
rect 19962 9766 20014 9818
rect 1400 9664 1452 9716
rect 3148 9664 3200 9716
rect 6644 9707 6696 9716
rect 6644 9673 6653 9707
rect 6653 9673 6687 9707
rect 6687 9673 6696 9707
rect 6644 9664 6696 9673
rect 8116 9707 8168 9716
rect 8116 9673 8125 9707
rect 8125 9673 8159 9707
rect 8159 9673 8168 9707
rect 8116 9664 8168 9673
rect 12808 9707 12860 9716
rect 12808 9673 12817 9707
rect 12817 9673 12851 9707
rect 12851 9673 12860 9707
rect 12808 9664 12860 9673
rect 18420 9664 18472 9716
rect 19156 9664 19208 9716
rect 2136 9639 2188 9648
rect 2136 9605 2145 9639
rect 2145 9605 2179 9639
rect 2179 9605 2188 9639
rect 2136 9596 2188 9605
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 5448 9596 5500 9648
rect 18696 9639 18748 9648
rect 18696 9605 18705 9639
rect 18705 9605 18739 9639
rect 18739 9605 18748 9639
rect 18696 9596 18748 9605
rect 7288 9528 7340 9580
rect 1676 9392 1728 9444
rect 7932 9392 7984 9444
rect 12900 9528 12952 9580
rect 9496 9460 9548 9512
rect 14556 9460 14608 9512
rect 14096 9392 14148 9444
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 9128 9324 9180 9376
rect 16672 9324 16724 9376
rect 17132 9324 17184 9376
rect 8497 9222 8549 9274
rect 8561 9222 8613 9274
rect 8625 9222 8677 9274
rect 8689 9222 8741 9274
rect 16012 9222 16064 9274
rect 16076 9222 16128 9274
rect 16140 9222 16192 9274
rect 16204 9222 16256 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 2136 9120 2188 9172
rect 7288 9120 7340 9172
rect 20076 9120 20128 9172
rect 7472 9052 7524 9104
rect 9128 9052 9180 9104
rect 16672 9052 16724 9104
rect 3976 8984 4028 9036
rect 9496 8984 9548 9036
rect 12072 8984 12124 9036
rect 18788 8984 18840 9036
rect 19432 8984 19484 9036
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2688 8916 2740 8925
rect 7748 8959 7800 8968
rect 5724 8848 5776 8900
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 14096 8959 14148 8968
rect 14096 8925 14105 8959
rect 14105 8925 14139 8959
rect 14139 8925 14148 8959
rect 14096 8916 14148 8925
rect 18144 8959 18196 8968
rect 18144 8925 18153 8959
rect 18153 8925 18187 8959
rect 18187 8925 18196 8959
rect 18144 8916 18196 8925
rect 7932 8848 7984 8900
rect 11704 8848 11756 8900
rect 17132 8891 17184 8900
rect 1676 8823 1728 8832
rect 1676 8789 1685 8823
rect 1685 8789 1719 8823
rect 1719 8789 1728 8823
rect 1676 8780 1728 8789
rect 2228 8780 2280 8832
rect 9404 8780 9456 8832
rect 17132 8857 17141 8891
rect 17141 8857 17175 8891
rect 17175 8857 17184 8891
rect 17132 8848 17184 8857
rect 4739 8678 4791 8730
rect 4803 8678 4855 8730
rect 4867 8678 4919 8730
rect 4931 8678 4983 8730
rect 12255 8678 12307 8730
rect 12319 8678 12371 8730
rect 12383 8678 12435 8730
rect 12447 8678 12499 8730
rect 19770 8678 19822 8730
rect 19834 8678 19886 8730
rect 19898 8678 19950 8730
rect 19962 8678 20014 8730
rect 2136 8576 2188 8628
rect 7472 8576 7524 8628
rect 9496 8619 9548 8628
rect 9496 8585 9505 8619
rect 9505 8585 9539 8619
rect 9539 8585 9548 8619
rect 9496 8576 9548 8585
rect 12072 8576 12124 8628
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 16672 8576 16724 8628
rect 19432 8619 19484 8628
rect 19432 8585 19441 8619
rect 19441 8585 19475 8619
rect 19475 8585 19484 8619
rect 19432 8576 19484 8585
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 2688 8440 2740 8492
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 14096 8440 14148 8492
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 18144 8440 18196 8492
rect 19156 8440 19208 8492
rect 2504 8347 2556 8356
rect 2504 8313 2513 8347
rect 2513 8313 2547 8347
rect 2547 8313 2556 8347
rect 2504 8304 2556 8313
rect 5448 8304 5500 8356
rect 9680 8347 9732 8356
rect 1860 8236 1912 8288
rect 3976 8279 4028 8288
rect 3976 8245 3985 8279
rect 3985 8245 4019 8279
rect 4019 8245 4028 8279
rect 3976 8236 4028 8245
rect 5724 8279 5776 8288
rect 5724 8245 5733 8279
rect 5733 8245 5767 8279
rect 5767 8245 5776 8279
rect 5724 8236 5776 8245
rect 9680 8313 9689 8347
rect 9689 8313 9723 8347
rect 9723 8313 9732 8347
rect 9680 8304 9732 8313
rect 14096 8347 14148 8356
rect 14096 8313 14105 8347
rect 14105 8313 14139 8347
rect 14139 8313 14148 8347
rect 14096 8304 14148 8313
rect 9036 8236 9088 8288
rect 10048 8236 10100 8288
rect 16396 8236 16448 8288
rect 17776 8279 17828 8288
rect 17776 8245 17785 8279
rect 17785 8245 17819 8279
rect 17819 8245 17828 8279
rect 17776 8236 17828 8245
rect 19064 8279 19116 8288
rect 19064 8245 19073 8279
rect 19073 8245 19107 8279
rect 19107 8245 19116 8279
rect 19064 8236 19116 8245
rect 8497 8134 8549 8186
rect 8561 8134 8613 8186
rect 8625 8134 8677 8186
rect 8689 8134 8741 8186
rect 16012 8134 16064 8186
rect 16076 8134 16128 8186
rect 16140 8134 16192 8186
rect 16204 8134 16256 8186
rect 5724 8032 5776 8084
rect 9680 8032 9732 8084
rect 14096 8032 14148 8084
rect 17776 8032 17828 8084
rect 1952 7964 2004 8016
rect 2228 7964 2280 8016
rect 2504 8007 2556 8016
rect 2504 7973 2513 8007
rect 2513 7973 2547 8007
rect 2547 7973 2556 8007
rect 2504 7964 2556 7973
rect 4620 7939 4672 7948
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 10692 7896 10744 7948
rect 11704 7896 11756 7948
rect 12624 7896 12676 7948
rect 15568 7896 15620 7948
rect 17868 7896 17920 7948
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 7748 7828 7800 7880
rect 8392 7828 8444 7880
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 19156 7871 19208 7880
rect 19156 7837 19165 7871
rect 19165 7837 19199 7871
rect 19199 7837 19208 7871
rect 19156 7828 19208 7837
rect 12992 7692 13044 7744
rect 16396 7735 16448 7744
rect 16396 7701 16405 7735
rect 16405 7701 16439 7735
rect 16439 7701 16448 7735
rect 16396 7692 16448 7701
rect 19248 7692 19300 7744
rect 4739 7590 4791 7642
rect 4803 7590 4855 7642
rect 4867 7590 4919 7642
rect 4931 7590 4983 7642
rect 12255 7590 12307 7642
rect 12319 7590 12371 7642
rect 12383 7590 12435 7642
rect 12447 7590 12499 7642
rect 19770 7590 19822 7642
rect 19834 7590 19886 7642
rect 19898 7590 19950 7642
rect 19962 7590 20014 7642
rect 1676 7488 1728 7540
rect 4620 7531 4672 7540
rect 4620 7497 4629 7531
rect 4629 7497 4663 7531
rect 4663 7497 4672 7531
rect 4620 7488 4672 7497
rect 9772 7488 9824 7540
rect 11704 7531 11756 7540
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 12624 7488 12676 7540
rect 16488 7531 16540 7540
rect 16488 7497 16497 7531
rect 16497 7497 16531 7531
rect 16531 7497 16540 7531
rect 16488 7488 16540 7497
rect 17868 7531 17920 7540
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 18696 7531 18748 7540
rect 17868 7488 17920 7497
rect 8392 7463 8444 7472
rect 8392 7429 8401 7463
rect 8401 7429 8435 7463
rect 8435 7429 8444 7463
rect 8392 7420 8444 7429
rect 9956 7463 10008 7472
rect 2504 7352 2556 7404
rect 4160 7352 4212 7404
rect 4344 7352 4396 7404
rect 5448 7395 5500 7404
rect 5448 7361 5457 7395
rect 5457 7361 5491 7395
rect 5491 7361 5500 7395
rect 9956 7429 9965 7463
rect 9965 7429 9999 7463
rect 9999 7429 10008 7463
rect 9956 7420 10008 7429
rect 5448 7352 5500 7361
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 1860 7327 1912 7336
rect 1860 7293 1869 7327
rect 1869 7293 1903 7327
rect 1903 7293 1912 7327
rect 1860 7284 1912 7293
rect 16580 7420 16632 7472
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 2596 7148 2648 7200
rect 4620 7216 4672 7268
rect 7564 7216 7616 7268
rect 7932 7216 7984 7268
rect 16488 7284 16540 7336
rect 18696 7497 18705 7531
rect 18705 7497 18739 7531
rect 18739 7497 18748 7531
rect 18696 7488 18748 7497
rect 18328 7352 18380 7404
rect 13636 7259 13688 7268
rect 13636 7225 13645 7259
rect 13645 7225 13679 7259
rect 13679 7225 13688 7259
rect 13636 7216 13688 7225
rect 18880 7216 18932 7268
rect 7748 7148 7800 7200
rect 11152 7148 11204 7200
rect 15568 7148 15620 7200
rect 18788 7148 18840 7200
rect 8497 7046 8549 7098
rect 8561 7046 8613 7098
rect 8625 7046 8677 7098
rect 8689 7046 8741 7098
rect 16012 7046 16064 7098
rect 16076 7046 16128 7098
rect 16140 7046 16192 7098
rect 16204 7046 16256 7098
rect 2228 6944 2280 6996
rect 7564 6987 7616 6996
rect 7564 6953 7573 6987
rect 7573 6953 7607 6987
rect 7607 6953 7616 6987
rect 7564 6944 7616 6953
rect 7748 6944 7800 6996
rect 16396 6944 16448 6996
rect 18880 6987 18932 6996
rect 18880 6953 18889 6987
rect 18889 6953 18923 6987
rect 18923 6953 18932 6987
rect 18880 6944 18932 6953
rect 1952 6919 2004 6928
rect 1952 6885 1961 6919
rect 1961 6885 1995 6919
rect 1995 6885 2004 6919
rect 1952 6876 2004 6885
rect 4160 6919 4212 6928
rect 4160 6885 4169 6919
rect 4169 6885 4203 6919
rect 4203 6885 4212 6919
rect 4160 6876 4212 6885
rect 11152 6876 11204 6928
rect 19248 6919 19300 6928
rect 19248 6885 19257 6919
rect 19257 6885 19291 6919
rect 19291 6885 19300 6919
rect 19248 6876 19300 6885
rect 2504 6808 2556 6860
rect 8852 6808 8904 6860
rect 13084 6808 13136 6860
rect 14556 6808 14608 6860
rect 16488 6808 16540 6860
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 12716 6740 12768 6792
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 6276 6715 6328 6724
rect 6276 6681 6285 6715
rect 6285 6681 6319 6715
rect 6319 6681 6328 6715
rect 6276 6672 6328 6681
rect 18236 6715 18288 6724
rect 18236 6681 18245 6715
rect 18245 6681 18279 6715
rect 18279 6681 18288 6715
rect 18236 6672 18288 6681
rect 19432 6672 19484 6724
rect 2780 6604 2832 6656
rect 11704 6604 11756 6656
rect 13452 6604 13504 6656
rect 4739 6502 4791 6554
rect 4803 6502 4855 6554
rect 4867 6502 4919 6554
rect 4931 6502 4983 6554
rect 12255 6502 12307 6554
rect 12319 6502 12371 6554
rect 12383 6502 12435 6554
rect 12447 6502 12499 6554
rect 19770 6502 19822 6554
rect 19834 6502 19886 6554
rect 19898 6502 19950 6554
rect 19962 6502 20014 6554
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 11152 6400 11204 6452
rect 13084 6400 13136 6452
rect 17684 6443 17736 6452
rect 17684 6409 17693 6443
rect 17693 6409 17727 6443
rect 17727 6409 17736 6443
rect 17684 6400 17736 6409
rect 19064 6400 19116 6452
rect 19248 6400 19300 6452
rect 2688 6332 2740 6384
rect 5724 6375 5776 6384
rect 5724 6341 5733 6375
rect 5733 6341 5767 6375
rect 5767 6341 5776 6375
rect 5724 6332 5776 6341
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 2780 6264 2832 6273
rect 4344 6264 4396 6316
rect 8392 6264 8444 6316
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 13636 6264 13688 6316
rect 19432 6307 19484 6316
rect 19432 6273 19441 6307
rect 19441 6273 19475 6307
rect 19475 6273 19484 6307
rect 19432 6264 19484 6273
rect 3240 6128 3292 6180
rect 3424 6171 3476 6180
rect 3424 6137 3433 6171
rect 3433 6137 3467 6171
rect 3467 6137 3476 6171
rect 3424 6128 3476 6137
rect 5080 6060 5132 6112
rect 8024 6103 8076 6112
rect 8024 6069 8033 6103
rect 8033 6069 8067 6103
rect 8067 6069 8076 6103
rect 11060 6128 11112 6180
rect 19156 6171 19208 6180
rect 19156 6137 19165 6171
rect 19165 6137 19199 6171
rect 19199 6137 19208 6171
rect 19156 6128 19208 6137
rect 8024 6060 8076 6069
rect 8852 6060 8904 6112
rect 9864 6103 9916 6112
rect 9864 6069 9873 6103
rect 9873 6069 9907 6103
rect 9907 6069 9916 6103
rect 9864 6060 9916 6069
rect 14556 6060 14608 6112
rect 16488 6060 16540 6112
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 8497 5958 8549 6010
rect 8561 5958 8613 6010
rect 8625 5958 8677 6010
rect 8689 5958 8741 6010
rect 16012 5958 16064 6010
rect 16076 5958 16128 6010
rect 16140 5958 16192 6010
rect 16204 5958 16256 6010
rect 8024 5856 8076 5908
rect 9864 5856 9916 5908
rect 3424 5788 3476 5840
rect 5724 5788 5776 5840
rect 9772 5788 9824 5840
rect 11704 5831 11756 5840
rect 11704 5797 11713 5831
rect 11713 5797 11747 5831
rect 11747 5797 11756 5831
rect 11704 5788 11756 5797
rect 5356 5720 5408 5772
rect 6552 5763 6604 5772
rect 6552 5729 6596 5763
rect 6596 5729 6604 5763
rect 6552 5720 6604 5729
rect 7840 5720 7892 5772
rect 7932 5720 7984 5772
rect 9128 5720 9180 5772
rect 13084 5720 13136 5772
rect 16672 5720 16724 5772
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 11060 5652 11112 5704
rect 18972 5695 19024 5704
rect 18972 5661 18981 5695
rect 18981 5661 19015 5695
rect 19015 5661 19024 5695
rect 18972 5652 19024 5661
rect 19432 5695 19484 5704
rect 19432 5661 19441 5695
rect 19441 5661 19475 5695
rect 19475 5661 19484 5695
rect 19432 5652 19484 5661
rect 7656 5516 7708 5568
rect 12624 5516 12676 5568
rect 15660 5516 15712 5568
rect 4739 5414 4791 5466
rect 4803 5414 4855 5466
rect 4867 5414 4919 5466
rect 4931 5414 4983 5466
rect 12255 5414 12307 5466
rect 12319 5414 12371 5466
rect 12383 5414 12435 5466
rect 12447 5414 12499 5466
rect 19770 5414 19822 5466
rect 19834 5414 19886 5466
rect 19898 5414 19950 5466
rect 19962 5414 20014 5466
rect 2136 5312 2188 5364
rect 3240 5312 3292 5364
rect 3884 5312 3936 5364
rect 6552 5355 6604 5364
rect 6552 5321 6561 5355
rect 6561 5321 6595 5355
rect 6595 5321 6604 5355
rect 6552 5312 6604 5321
rect 9128 5355 9180 5364
rect 9128 5321 9137 5355
rect 9137 5321 9171 5355
rect 9171 5321 9180 5355
rect 9128 5312 9180 5321
rect 9772 5312 9824 5364
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 11704 5355 11756 5364
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 13084 5312 13136 5364
rect 16672 5355 16724 5364
rect 16672 5321 16681 5355
rect 16681 5321 16715 5355
rect 16715 5321 16724 5355
rect 16672 5312 16724 5321
rect 18972 5312 19024 5364
rect 1216 5176 1268 5228
rect 3332 5244 3384 5296
rect 10416 5219 10468 5228
rect 10416 5185 10425 5219
rect 10425 5185 10459 5219
rect 10459 5185 10468 5219
rect 10416 5176 10468 5185
rect 12624 5176 12676 5228
rect 12716 5176 12768 5228
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 19156 5176 19208 5228
rect 5080 5108 5132 5160
rect 3884 5083 3936 5092
rect 3884 5049 3893 5083
rect 3893 5049 3927 5083
rect 3927 5049 3936 5083
rect 3884 5040 3936 5049
rect 4528 5083 4580 5092
rect 4528 5049 4537 5083
rect 4537 5049 4571 5083
rect 4571 5049 4580 5083
rect 4528 5040 4580 5049
rect 7932 5040 7984 5092
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 5724 4972 5776 5024
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 7840 5015 7892 5024
rect 5816 4972 5868 4981
rect 7840 4981 7849 5015
rect 7849 4981 7883 5015
rect 7883 4981 7892 5015
rect 7840 4972 7892 4981
rect 8944 4972 8996 5024
rect 9404 4972 9456 5024
rect 10692 4972 10744 5024
rect 18604 5108 18656 5160
rect 20168 5244 20220 5296
rect 16304 5083 16356 5092
rect 16304 5049 16313 5083
rect 16313 5049 16347 5083
rect 16347 5049 16356 5083
rect 16304 5040 16356 5049
rect 15384 4972 15436 5024
rect 8497 4870 8549 4922
rect 8561 4870 8613 4922
rect 8625 4870 8677 4922
rect 8689 4870 8741 4922
rect 16012 4870 16064 4922
rect 16076 4870 16128 4922
rect 16140 4870 16192 4922
rect 16204 4870 16256 4922
rect 4804 4768 4856 4820
rect 6552 4768 6604 4820
rect 10692 4768 10744 4820
rect 5724 4700 5776 4752
rect 6184 4700 6236 4752
rect 7656 4743 7708 4752
rect 7656 4709 7665 4743
rect 7665 4709 7699 4743
rect 7699 4709 7708 4743
rect 7656 4700 7708 4709
rect 10416 4743 10468 4752
rect 10416 4709 10425 4743
rect 10425 4709 10459 4743
rect 10459 4709 10468 4743
rect 10416 4700 10468 4709
rect 12716 4700 12768 4752
rect 15384 4743 15436 4752
rect 15384 4709 15393 4743
rect 15393 4709 15427 4743
rect 15427 4709 15436 4743
rect 15384 4700 15436 4709
rect 15752 4700 15804 4752
rect 16304 4700 16356 4752
rect 18788 4700 18840 4752
rect 3056 4564 3108 4616
rect 4620 4564 4672 4616
rect 7932 4607 7984 4616
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 19340 4607 19392 4616
rect 19340 4573 19349 4607
rect 19349 4573 19383 4607
rect 19383 4573 19392 4607
rect 19340 4564 19392 4573
rect 5080 4539 5132 4548
rect 5080 4505 5089 4539
rect 5089 4505 5123 4539
rect 5123 4505 5132 4539
rect 5080 4496 5132 4505
rect 16856 4496 16908 4548
rect 16304 4428 16356 4480
rect 4739 4326 4791 4378
rect 4803 4326 4855 4378
rect 4867 4326 4919 4378
rect 4931 4326 4983 4378
rect 12255 4326 12307 4378
rect 12319 4326 12371 4378
rect 12383 4326 12435 4378
rect 12447 4326 12499 4378
rect 19770 4326 19822 4378
rect 19834 4326 19886 4378
rect 19898 4326 19950 4378
rect 19962 4326 20014 4378
rect 4620 4224 4672 4276
rect 6184 4267 6236 4276
rect 6184 4233 6193 4267
rect 6193 4233 6227 4267
rect 6227 4233 6236 4267
rect 6184 4224 6236 4233
rect 7656 4224 7708 4276
rect 7932 4156 7984 4208
rect 9772 4224 9824 4276
rect 11980 4267 12032 4276
rect 11980 4233 11989 4267
rect 11989 4233 12023 4267
rect 12023 4233 12032 4267
rect 11980 4224 12032 4233
rect 15384 4267 15436 4276
rect 15384 4233 15393 4267
rect 15393 4233 15427 4267
rect 15427 4233 15436 4267
rect 15384 4224 15436 4233
rect 19340 4224 19392 4276
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 11704 4156 11756 4208
rect 12716 4088 12768 4140
rect 14464 4131 14516 4140
rect 7288 4063 7340 4072
rect 7288 4029 7306 4063
rect 7306 4029 7340 4063
rect 10692 4063 10744 4072
rect 7288 4020 7340 4029
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 20260 4088 20312 4140
rect 10692 4020 10744 4029
rect 8944 3952 8996 4004
rect 13176 3995 13228 4004
rect 13176 3961 13185 3995
rect 13185 3961 13219 3995
rect 13219 3961 13228 3995
rect 13176 3952 13228 3961
rect 15752 3995 15804 4004
rect 15752 3961 15761 3995
rect 15761 3961 15795 3995
rect 15795 3961 15804 3995
rect 15752 3952 15804 3961
rect 16856 3995 16908 4004
rect 16856 3961 16865 3995
rect 16865 3961 16899 3995
rect 16899 3961 16908 3995
rect 16856 3952 16908 3961
rect 2136 3884 2188 3936
rect 3056 3927 3108 3936
rect 3056 3893 3065 3927
rect 3065 3893 3099 3927
rect 3099 3893 3108 3927
rect 3056 3884 3108 3893
rect 3608 3927 3660 3936
rect 3608 3893 3617 3927
rect 3617 3893 3651 3927
rect 3651 3893 3660 3927
rect 3608 3884 3660 3893
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 7564 3884 7616 3936
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 11244 3884 11296 3936
rect 18512 3884 18564 3936
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 8497 3782 8549 3834
rect 8561 3782 8613 3834
rect 8625 3782 8677 3834
rect 8689 3782 8741 3834
rect 16012 3782 16064 3834
rect 16076 3782 16128 3834
rect 16140 3782 16192 3834
rect 16204 3782 16256 3834
rect 2136 3655 2188 3664
rect 2136 3621 2145 3655
rect 2145 3621 2179 3655
rect 2179 3621 2188 3655
rect 2136 3612 2188 3621
rect 7564 3655 7616 3664
rect 7564 3621 7573 3655
rect 7573 3621 7607 3655
rect 7607 3621 7616 3655
rect 7564 3612 7616 3621
rect 10416 3655 10468 3664
rect 10416 3621 10425 3655
rect 10425 3621 10459 3655
rect 10459 3621 10468 3655
rect 10416 3612 10468 3621
rect 4528 3544 4580 3596
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 11980 3544 12032 3596
rect 13452 3587 13504 3596
rect 13452 3553 13496 3587
rect 13496 3553 13504 3587
rect 13452 3544 13504 3553
rect 19524 3544 19576 3596
rect 5448 3476 5500 3528
rect 6000 3476 6052 3528
rect 10048 3476 10100 3528
rect 15384 3519 15436 3528
rect 12624 3408 12676 3460
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 16948 3519 17000 3528
rect 16948 3485 16957 3519
rect 16957 3485 16991 3519
rect 16991 3485 17000 3519
rect 16948 3476 17000 3485
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 17224 3476 17276 3485
rect 18420 3519 18472 3528
rect 18420 3485 18429 3519
rect 18429 3485 18463 3519
rect 18463 3485 18472 3519
rect 18420 3476 18472 3485
rect 4620 3340 4672 3392
rect 7012 3340 7064 3392
rect 12072 3340 12124 3392
rect 12808 3340 12860 3392
rect 12992 3340 13044 3392
rect 19616 3340 19668 3392
rect 4739 3238 4791 3290
rect 4803 3238 4855 3290
rect 4867 3238 4919 3290
rect 4931 3238 4983 3290
rect 12255 3238 12307 3290
rect 12319 3238 12371 3290
rect 12383 3238 12435 3290
rect 12447 3238 12499 3290
rect 19770 3238 19822 3290
rect 19834 3238 19886 3290
rect 19898 3238 19950 3290
rect 19962 3238 20014 3290
rect 2136 3179 2188 3188
rect 2136 3145 2145 3179
rect 2145 3145 2179 3179
rect 2179 3145 2188 3179
rect 2136 3136 2188 3145
rect 3608 3136 3660 3188
rect 5724 3136 5776 3188
rect 6368 3068 6420 3120
rect 4620 3000 4672 3052
rect 7564 3136 7616 3188
rect 10048 3179 10100 3188
rect 10048 3145 10057 3179
rect 10057 3145 10091 3179
rect 10091 3145 10100 3179
rect 10048 3136 10100 3145
rect 6644 3068 6696 3120
rect 5448 2975 5500 2984
rect 5448 2941 5457 2975
rect 5457 2941 5491 2975
rect 5491 2941 5500 2975
rect 5448 2932 5500 2941
rect 6644 2932 6696 2984
rect 12992 3136 13044 3188
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 15384 3136 15436 3188
rect 16948 3136 17000 3188
rect 11336 3068 11388 3120
rect 14924 3111 14976 3120
rect 14924 3077 14933 3111
rect 14933 3077 14967 3111
rect 14967 3077 14976 3111
rect 14924 3068 14976 3077
rect 12624 3000 12676 3052
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 17224 3068 17276 3120
rect 19616 3068 19668 3120
rect 16856 3043 16908 3052
rect 13176 3000 13228 3009
rect 14924 2932 14976 2984
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 18420 3000 18472 3052
rect 3884 2839 3936 2848
rect 3884 2805 3893 2839
rect 3893 2805 3927 2839
rect 3927 2805 3936 2839
rect 3884 2796 3936 2805
rect 4620 2796 4672 2848
rect 8208 2796 8260 2848
rect 8392 2796 8444 2848
rect 10140 2864 10192 2916
rect 10232 2864 10284 2916
rect 11980 2864 12032 2916
rect 13452 2864 13504 2916
rect 18788 2907 18840 2916
rect 18788 2873 18797 2907
rect 18797 2873 18831 2907
rect 18831 2873 18840 2907
rect 18788 2864 18840 2873
rect 10968 2796 11020 2848
rect 17316 2796 17368 2848
rect 19524 2839 19576 2848
rect 19524 2805 19533 2839
rect 19533 2805 19567 2839
rect 19567 2805 19576 2839
rect 19524 2796 19576 2805
rect 21732 2796 21784 2848
rect 8497 2694 8549 2746
rect 8561 2694 8613 2746
rect 8625 2694 8677 2746
rect 8689 2694 8741 2746
rect 16012 2694 16064 2746
rect 16076 2694 16128 2746
rect 16140 2694 16192 2746
rect 16204 2694 16256 2746
rect 8392 2592 8444 2644
rect 9404 2635 9456 2644
rect 9404 2601 9413 2635
rect 9413 2601 9447 2635
rect 9447 2601 9456 2635
rect 9404 2592 9456 2601
rect 2504 2456 2556 2508
rect 4620 2456 4672 2508
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 10140 2524 10192 2576
rect 8208 2499 8260 2508
rect 8208 2465 8217 2499
rect 8217 2465 8251 2499
rect 8251 2465 8260 2499
rect 12624 2592 12676 2644
rect 13452 2524 13504 2576
rect 8208 2456 8260 2465
rect 16304 2592 16356 2644
rect 17316 2592 17368 2644
rect 19616 2635 19668 2644
rect 18512 2524 18564 2576
rect 16488 2456 16540 2508
rect 19616 2601 19625 2635
rect 19625 2601 19659 2635
rect 19659 2601 19668 2635
rect 19616 2592 19668 2601
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 13176 2320 13228 2372
rect 17316 2320 17368 2372
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 4620 2252 4672 2304
rect 13820 2252 13872 2304
rect 14280 2252 14332 2304
rect 19432 2252 19484 2304
rect 4739 2150 4791 2202
rect 4803 2150 4855 2202
rect 4867 2150 4919 2202
rect 4931 2150 4983 2202
rect 12255 2150 12307 2202
rect 12319 2150 12371 2202
rect 12383 2150 12435 2202
rect 12447 2150 12499 2202
rect 19770 2150 19822 2202
rect 19834 2150 19886 2202
rect 19898 2150 19950 2202
rect 19962 2150 20014 2202
rect 12808 76 12860 128
rect 18420 76 18472 128
rect 20720 76 20772 128
rect 21364 76 21416 128
<< metal2 >>
rect 570 24210 626 24690
rect 1674 24210 1730 24690
rect 2870 24290 2926 24690
rect 2780 24268 2832 24274
rect 2780 24210 2832 24216
rect 2870 24262 3372 24290
rect 2870 24210 2926 24262
rect 18 24032 74 24041
rect 18 23967 74 23976
rect 32 22098 60 23967
rect 110 22672 166 22681
rect 110 22607 166 22616
rect 20 22092 72 22098
rect 20 22034 72 22040
rect 124 22030 152 22607
rect 112 22024 164 22030
rect 112 21966 164 21972
rect 1584 21004 1636 21010
rect 1584 20946 1636 20952
rect 1596 20777 1624 20946
rect 1952 20800 2004 20806
rect 1582 20768 1638 20777
rect 1952 20742 2004 20748
rect 1582 20703 1638 20712
rect 1596 20602 1624 20703
rect 1964 20602 1992 20742
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 1596 18970 1624 19343
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 18426 1440 18770
rect 1400 18420 1452 18426
rect 1400 18362 1452 18368
rect 1412 17882 1440 18362
rect 1400 17876 1452 17882
rect 1400 17818 1452 17824
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1780 16998 1808 17682
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 112 10600 164 10606
rect 112 10542 164 10548
rect 124 10305 152 10542
rect 110 10296 166 10305
rect 110 10231 166 10240
rect 1412 9722 1440 11086
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1688 8838 1716 9386
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 7546 1716 8774
rect 1872 8498 1900 10406
rect 1964 10062 1992 10474
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1964 9178 1992 9998
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 2148 9654 2176 9930
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2148 9178 2176 9590
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2148 8634 2176 9114
rect 2700 8974 2728 16934
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1858 8392 1914 8401
rect 1858 8327 1914 8336
rect 1872 8294 1900 8327
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1872 7342 1900 8230
rect 2240 8022 2268 8774
rect 2700 8498 2728 8910
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2516 8022 2544 8298
rect 1952 8016 2004 8022
rect 1952 7958 2004 7964
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1964 6934 1992 7958
rect 2516 7410 2544 7958
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2228 7200 2280 7206
rect 2596 7200 2648 7206
rect 2228 7142 2280 7148
rect 2516 7160 2596 7188
rect 2240 7002 2268 7142
rect 2516 7041 2544 7160
rect 2596 7142 2648 7148
rect 2502 7032 2558 7041
rect 2228 6996 2280 7002
rect 2502 6967 2558 6976
rect 2228 6938 2280 6944
rect 1952 6928 2004 6934
rect 1952 6870 2004 6876
rect 2516 6866 2544 6967
rect 2792 6882 2820 24210
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2884 17338 2912 20266
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3160 9586 3188 9658
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2700 6854 2820 6882
rect 2516 6458 2544 6802
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2700 6390 2728 6854
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2792 6322 2820 6598
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 2136 5704 2188 5710
rect 1214 5672 1270 5681
rect 2136 5646 2188 5652
rect 1214 5607 1270 5616
rect 1228 5234 1256 5607
rect 2148 5370 2176 5646
rect 3252 5370 3280 6122
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3344 5302 3372 24262
rect 4066 24268 4122 24690
rect 4066 24216 4068 24268
rect 4120 24216 4122 24268
rect 4066 24210 4122 24216
rect 5262 24268 5318 24690
rect 6458 24290 6514 24690
rect 7654 24290 7710 24690
rect 5262 24216 5264 24268
rect 5316 24216 5318 24268
rect 5262 24210 5318 24216
rect 6196 24262 6514 24290
rect 4080 24179 4108 24210
rect 5276 24179 5304 24210
rect 4713 21788 5009 21808
rect 4769 21786 4793 21788
rect 4849 21786 4873 21788
rect 4929 21786 4953 21788
rect 4791 21734 4793 21786
rect 4855 21734 4867 21786
rect 4929 21734 4931 21786
rect 4769 21732 4793 21734
rect 4849 21732 4873 21734
rect 4929 21732 4953 21734
rect 4713 21712 5009 21732
rect 4713 20700 5009 20720
rect 4769 20698 4793 20700
rect 4849 20698 4873 20700
rect 4929 20698 4953 20700
rect 4791 20646 4793 20698
rect 4855 20646 4867 20698
rect 4929 20646 4931 20698
rect 4769 20644 4793 20646
rect 4849 20644 4873 20646
rect 4929 20644 4953 20646
rect 4713 20624 5009 20644
rect 4713 19612 5009 19632
rect 4769 19610 4793 19612
rect 4849 19610 4873 19612
rect 4929 19610 4953 19612
rect 4791 19558 4793 19610
rect 4855 19558 4867 19610
rect 4929 19558 4931 19610
rect 4769 19556 4793 19558
rect 4849 19556 4873 19558
rect 4929 19556 4953 19558
rect 4713 19536 5009 19556
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 4713 18524 5009 18544
rect 4769 18522 4793 18524
rect 4849 18522 4873 18524
rect 4929 18522 4953 18524
rect 4791 18470 4793 18522
rect 4855 18470 4867 18522
rect 4929 18470 4931 18522
rect 4769 18468 4793 18470
rect 4849 18468 4873 18470
rect 4929 18468 4953 18470
rect 4713 18448 5009 18468
rect 6104 17746 6132 18566
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 4713 17436 5009 17456
rect 4769 17434 4793 17436
rect 4849 17434 4873 17436
rect 4929 17434 4953 17436
rect 4791 17382 4793 17434
rect 4855 17382 4867 17434
rect 4929 17382 4931 17434
rect 4769 17380 4793 17382
rect 4849 17380 4873 17382
rect 4929 17380 4953 17382
rect 4713 17360 5009 17380
rect 6104 17338 6132 17682
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 5354 16688 5410 16697
rect 5354 16623 5410 16632
rect 4713 16348 5009 16368
rect 4769 16346 4793 16348
rect 4849 16346 4873 16348
rect 4929 16346 4953 16348
rect 4791 16294 4793 16346
rect 4855 16294 4867 16346
rect 4929 16294 4931 16346
rect 4769 16292 4793 16294
rect 4849 16292 4873 16294
rect 4929 16292 4953 16294
rect 4713 16272 5009 16292
rect 4713 15260 5009 15280
rect 4769 15258 4793 15260
rect 4849 15258 4873 15260
rect 4929 15258 4953 15260
rect 4791 15206 4793 15258
rect 4855 15206 4867 15258
rect 4929 15206 4931 15258
rect 4769 15204 4793 15206
rect 4849 15204 4873 15206
rect 4929 15204 4953 15206
rect 4713 15184 5009 15204
rect 4713 14172 5009 14192
rect 4769 14170 4793 14172
rect 4849 14170 4873 14172
rect 4929 14170 4953 14172
rect 4791 14118 4793 14170
rect 4855 14118 4867 14170
rect 4929 14118 4931 14170
rect 4769 14116 4793 14118
rect 4849 14116 4873 14118
rect 4929 14116 4953 14118
rect 4713 14096 5009 14116
rect 4713 13084 5009 13104
rect 4769 13082 4793 13084
rect 4849 13082 4873 13084
rect 4929 13082 4953 13084
rect 4791 13030 4793 13082
rect 4855 13030 4867 13082
rect 4929 13030 4931 13082
rect 4769 13028 4793 13030
rect 4849 13028 4873 13030
rect 4929 13028 4953 13030
rect 4713 13008 5009 13028
rect 4713 11996 5009 12016
rect 4769 11994 4793 11996
rect 4849 11994 4873 11996
rect 4929 11994 4953 11996
rect 4791 11942 4793 11994
rect 4855 11942 4867 11994
rect 4929 11942 4931 11994
rect 4769 11940 4793 11942
rect 4849 11940 4873 11942
rect 4929 11940 4953 11942
rect 4713 11920 5009 11940
rect 4713 10908 5009 10928
rect 4769 10906 4793 10908
rect 4849 10906 4873 10908
rect 4929 10906 4953 10908
rect 4791 10854 4793 10906
rect 4855 10854 4867 10906
rect 4929 10854 4931 10906
rect 4769 10852 4793 10854
rect 4849 10852 4873 10854
rect 4929 10852 4953 10854
rect 4713 10832 5009 10852
rect 4713 9820 5009 9840
rect 4769 9818 4793 9820
rect 4849 9818 4873 9820
rect 4929 9818 4953 9820
rect 4791 9766 4793 9818
rect 4855 9766 4867 9818
rect 4929 9766 4931 9818
rect 4769 9764 4793 9766
rect 4849 9764 4873 9766
rect 4929 9764 4953 9766
rect 4713 9744 5009 9764
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3988 8294 4016 8978
rect 4713 8732 5009 8752
rect 4769 8730 4793 8732
rect 4849 8730 4873 8732
rect 4929 8730 4953 8732
rect 4791 8678 4793 8730
rect 4855 8678 4867 8730
rect 4929 8678 4931 8730
rect 4769 8676 4793 8678
rect 4849 8676 4873 8678
rect 4929 8676 4953 8678
rect 4713 8656 5009 8676
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4632 7546 4660 7890
rect 4713 7644 5009 7664
rect 4769 7642 4793 7644
rect 4849 7642 4873 7644
rect 4929 7642 4953 7644
rect 4791 7590 4793 7642
rect 4855 7590 4867 7642
rect 4929 7590 4931 7642
rect 4769 7588 4793 7590
rect 4849 7588 4873 7590
rect 4929 7588 4953 7590
rect 4713 7568 5009 7588
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4172 6934 4200 7346
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4172 6458 4200 6870
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4356 6322 4384 7346
rect 4632 7274 4660 7482
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4713 6556 5009 6576
rect 4769 6554 4793 6556
rect 4849 6554 4873 6556
rect 4929 6554 4953 6556
rect 4791 6502 4793 6554
rect 4855 6502 4867 6554
rect 4929 6502 4931 6554
rect 4769 6500 4793 6502
rect 4849 6500 4873 6502
rect 4929 6500 4953 6502
rect 4713 6480 5009 6500
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3436 5846 3464 6122
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 3424 5840 3476 5846
rect 3424 5782 3476 5788
rect 3436 5681 3464 5782
rect 4620 5704 4672 5710
rect 3422 5672 3478 5681
rect 4620 5646 4672 5652
rect 3422 5607 3478 5616
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 1216 5228 1268 5234
rect 1216 5170 1268 5176
rect 3896 5098 3924 5306
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 3056 4616 3108 4622
rect 4540 4604 4568 5034
rect 4632 5012 4660 5646
rect 4713 5468 5009 5488
rect 4769 5466 4793 5468
rect 4849 5466 4873 5468
rect 4929 5466 4953 5468
rect 4791 5414 4793 5466
rect 4855 5414 4867 5466
rect 4929 5414 4931 5466
rect 4769 5412 4793 5414
rect 4849 5412 4873 5414
rect 4929 5412 4953 5414
rect 4713 5392 5009 5412
rect 5092 5166 5120 6054
rect 5368 5778 5396 16623
rect 6196 10266 6224 24262
rect 6458 24210 6514 24262
rect 7484 24262 7710 24290
rect 8850 24290 8906 24690
rect 10046 24290 10102 24690
rect 11242 24290 11298 24690
rect 12346 24290 12402 24690
rect 13542 24290 13598 24690
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6656 18290 6684 18770
rect 7484 18426 7512 24262
rect 7654 24210 7710 24262
rect 7840 24268 7892 24274
rect 7840 24210 7892 24216
rect 8850 24262 8984 24290
rect 8850 24210 8906 24262
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 6274 18048 6330 18057
rect 6274 17983 6330 17992
rect 6288 17882 6316 17983
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 7116 17338 7144 18158
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7668 17338 7696 17614
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7760 17105 7788 17138
rect 7746 17096 7802 17105
rect 7746 17031 7802 17040
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7392 14822 7420 15506
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 7300 10198 7328 10610
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5460 9654 5488 10066
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 9722 6684 9998
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 7300 9586 7328 10134
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7300 9178 7328 9522
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5460 7410 5488 8298
rect 5736 8294 5764 8842
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5736 8090 5764 8230
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6390 5764 6734
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5736 5846 5764 6326
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4804 5024 4856 5030
rect 4632 4984 4804 5012
rect 4804 4966 4856 4972
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 4816 4826 4844 4966
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 5736 4758 5764 4966
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 4620 4616 4672 4622
rect 4540 4576 4620 4604
rect 3056 4558 3108 4564
rect 4620 4558 4672 4564
rect 1858 4448 1914 4457
rect 1858 4383 1914 4392
rect 1872 4146 1900 4383
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 3068 3942 3096 4558
rect 4632 4282 4660 4558
rect 5080 4548 5132 4554
rect 5080 4490 5132 4496
rect 4713 4380 5009 4400
rect 4769 4378 4793 4380
rect 4849 4378 4873 4380
rect 4929 4378 4953 4380
rect 4791 4326 4793 4378
rect 4855 4326 4867 4378
rect 4929 4326 4931 4378
rect 4769 4324 4793 4326
rect 4849 4324 4873 4326
rect 4929 4324 4953 4326
rect 4713 4304 5009 4324
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 5092 4185 5120 4490
rect 5078 4176 5134 4185
rect 5078 4111 5134 4120
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 2148 3670 2176 3878
rect 2136 3664 2188 3670
rect 2136 3606 2188 3612
rect 2148 3194 2176 3606
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2516 2310 2544 2450
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 2009 2544 2246
rect 2502 2000 2558 2009
rect 2502 1935 2558 1944
rect 386 0 442 480
rect 1122 0 1178 480
rect 1858 0 1914 480
rect 2594 0 2650 480
rect 3068 82 3096 3878
rect 3620 3194 3648 3878
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3884 2848 3936 2854
rect 4540 2836 4568 3538
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 3058 4660 3334
rect 4713 3292 5009 3312
rect 4769 3290 4793 3292
rect 4849 3290 4873 3292
rect 4929 3290 4953 3292
rect 4791 3238 4793 3290
rect 4855 3238 4867 3290
rect 4929 3238 4931 3290
rect 4769 3236 4793 3238
rect 4849 3236 4873 3238
rect 4929 3236 4953 3238
rect 4713 3216 5009 3236
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 5460 2990 5488 3470
rect 5736 3194 5764 3878
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 4620 2848 4672 2854
rect 4540 2808 4620 2836
rect 3884 2790 3936 2796
rect 4620 2790 4672 2796
rect 3330 82 3386 480
rect 3068 54 3386 82
rect 3896 82 3924 2790
rect 4632 2514 4660 2790
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4632 2310 4660 2450
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 4066 82 4122 480
rect 3896 54 4122 82
rect 4632 82 4660 2246
rect 4713 2204 5009 2224
rect 4769 2202 4793 2204
rect 4849 2202 4873 2204
rect 4929 2202 4953 2204
rect 4791 2150 4793 2202
rect 4855 2150 4867 2202
rect 4929 2150 4931 2202
rect 4769 2148 4793 2150
rect 4849 2148 4873 2150
rect 4929 2148 4953 2150
rect 4713 2128 5009 2148
rect 4894 82 4950 480
rect 4632 54 4950 82
rect 3330 0 3386 54
rect 4066 0 4122 54
rect 4894 0 4950 54
rect 5630 82 5686 480
rect 5828 82 5856 4966
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 6196 4282 6224 4694
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6288 4185 6316 6666
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6564 5370 6592 5714
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6564 4826 6592 5306
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6274 4176 6330 4185
rect 7392 4154 7420 14758
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7484 10266 7512 10474
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7484 8634 7512 9046
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7760 8498 7788 8910
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7760 7886 7788 8434
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7576 7002 7604 7210
rect 7668 7188 7696 7822
rect 7852 7256 7880 24210
rect 8471 22332 8767 22352
rect 8527 22330 8551 22332
rect 8607 22330 8631 22332
rect 8687 22330 8711 22332
rect 8549 22278 8551 22330
rect 8613 22278 8625 22330
rect 8687 22278 8689 22330
rect 8527 22276 8551 22278
rect 8607 22276 8631 22278
rect 8687 22276 8711 22278
rect 8471 22256 8767 22276
rect 8471 21244 8767 21264
rect 8527 21242 8551 21244
rect 8607 21242 8631 21244
rect 8687 21242 8711 21244
rect 8549 21190 8551 21242
rect 8613 21190 8625 21242
rect 8687 21190 8689 21242
rect 8527 21188 8551 21190
rect 8607 21188 8631 21190
rect 8687 21188 8711 21190
rect 8471 21168 8767 21188
rect 8956 21146 8984 24262
rect 10046 24262 10364 24290
rect 10046 24210 10102 24262
rect 10336 21554 10364 24262
rect 10888 24262 11298 24290
rect 10324 21548 10376 21554
rect 10324 21490 10376 21496
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 8576 20936 8628 20942
rect 8576 20878 8628 20884
rect 8588 20602 8616 20878
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 9600 20330 9628 20946
rect 9588 20324 9640 20330
rect 9588 20266 9640 20272
rect 8471 20156 8767 20176
rect 8527 20154 8551 20156
rect 8607 20154 8631 20156
rect 8687 20154 8711 20156
rect 8549 20102 8551 20154
rect 8613 20102 8625 20154
rect 8687 20102 8689 20154
rect 8527 20100 8551 20102
rect 8607 20100 8631 20102
rect 8687 20100 8711 20102
rect 8471 20080 8767 20100
rect 8471 19068 8767 19088
rect 8527 19066 8551 19068
rect 8607 19066 8631 19068
rect 8687 19066 8711 19068
rect 8549 19014 8551 19066
rect 8613 19014 8625 19066
rect 8687 19014 8689 19066
rect 8527 19012 8551 19014
rect 8607 19012 8631 19014
rect 8687 19012 8711 19014
rect 8471 18992 8767 19012
rect 8850 18184 8906 18193
rect 8850 18119 8906 18128
rect 8864 18086 8892 18119
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 8471 17980 8767 18000
rect 8527 17978 8551 17980
rect 8607 17978 8631 17980
rect 8687 17978 8711 17980
rect 8549 17926 8551 17978
rect 8613 17926 8625 17978
rect 8687 17926 8689 17978
rect 8527 17924 8551 17926
rect 8607 17924 8631 17926
rect 8687 17924 8711 17926
rect 8471 17904 8767 17924
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8404 16998 8432 17138
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16590 8432 16934
rect 8471 16892 8767 16912
rect 8527 16890 8551 16892
rect 8607 16890 8631 16892
rect 8687 16890 8711 16892
rect 8549 16838 8551 16890
rect 8613 16838 8625 16890
rect 8687 16838 8689 16890
rect 8527 16836 8551 16838
rect 8607 16836 8631 16838
rect 8687 16836 8711 16838
rect 8471 16816 8767 16836
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 8036 15706 8064 15914
rect 8128 15910 8156 16526
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8471 15804 8767 15824
rect 8527 15802 8551 15804
rect 8607 15802 8631 15804
rect 8687 15802 8711 15804
rect 8549 15750 8551 15802
rect 8613 15750 8625 15802
rect 8687 15750 8689 15802
rect 8527 15748 8551 15750
rect 8607 15748 8631 15750
rect 8687 15748 8711 15750
rect 8471 15728 8767 15748
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 9140 15026 9168 15914
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9508 14929 9536 18022
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9692 15910 9720 16594
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9692 15570 9720 15846
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9494 14920 9550 14929
rect 8852 14884 8904 14890
rect 9494 14855 9550 14864
rect 8852 14826 8904 14832
rect 8471 14716 8767 14736
rect 8527 14714 8551 14716
rect 8607 14714 8631 14716
rect 8687 14714 8711 14716
rect 8549 14662 8551 14714
rect 8613 14662 8625 14714
rect 8687 14662 8689 14714
rect 8527 14660 8551 14662
rect 8607 14660 8631 14662
rect 8687 14660 8711 14662
rect 8471 14640 8767 14660
rect 8864 14618 8892 14826
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8471 13628 8767 13648
rect 8527 13626 8551 13628
rect 8607 13626 8631 13628
rect 8687 13626 8711 13628
rect 8549 13574 8551 13626
rect 8613 13574 8625 13626
rect 8687 13574 8689 13626
rect 8527 13572 8551 13574
rect 8607 13572 8631 13574
rect 8687 13572 8711 13574
rect 8471 13552 8767 13572
rect 8471 12540 8767 12560
rect 8527 12538 8551 12540
rect 8607 12538 8631 12540
rect 8687 12538 8711 12540
rect 8549 12486 8551 12538
rect 8613 12486 8625 12538
rect 8687 12486 8689 12538
rect 8527 12484 8551 12486
rect 8607 12484 8631 12486
rect 8687 12484 8711 12486
rect 8471 12464 8767 12484
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 8496 11898 8524 12174
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 9416 11762 9444 12174
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7944 11218 7972 11494
rect 8471 11452 8767 11472
rect 8527 11450 8551 11452
rect 8607 11450 8631 11452
rect 8687 11450 8711 11452
rect 8549 11398 8551 11450
rect 8613 11398 8625 11450
rect 8687 11398 8689 11450
rect 8527 11396 8551 11398
rect 8607 11396 8631 11398
rect 8687 11396 8711 11398
rect 8114 11384 8170 11393
rect 8471 11376 8767 11396
rect 8114 11319 8170 11328
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7944 10810 7972 11154
rect 8128 11082 8156 11319
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8471 10364 8767 10384
rect 8527 10362 8551 10364
rect 8607 10362 8631 10364
rect 8687 10362 8711 10364
rect 8549 10310 8551 10362
rect 8613 10310 8625 10362
rect 8687 10310 8689 10362
rect 8527 10308 8551 10310
rect 8607 10308 8631 10310
rect 8687 10308 8711 10310
rect 8471 10288 8767 10308
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8128 9722 8156 10066
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 9508 9518 9536 14855
rect 9770 14512 9826 14521
rect 9770 14447 9772 14456
rect 9824 14447 9826 14456
rect 9772 14418 9824 14424
rect 9784 14074 9812 14418
rect 10888 14074 10916 24262
rect 11242 24210 11298 24262
rect 12084 24262 12402 24290
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10980 13814 11008 21490
rect 12084 21146 12112 24262
rect 12346 24210 12402 24262
rect 13464 24262 13598 24290
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 12229 21788 12525 21808
rect 12285 21786 12309 21788
rect 12365 21786 12389 21788
rect 12445 21786 12469 21788
rect 12307 21734 12309 21786
rect 12371 21734 12383 21786
rect 12445 21734 12447 21786
rect 12285 21732 12309 21734
rect 12365 21732 12389 21734
rect 12445 21732 12469 21734
rect 12229 21712 12525 21732
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 13004 21010 13032 21966
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 12992 21004 13044 21010
rect 12992 20946 13044 20952
rect 12084 20262 12112 20946
rect 12229 20700 12525 20720
rect 12285 20698 12309 20700
rect 12365 20698 12389 20700
rect 12445 20698 12469 20700
rect 12307 20646 12309 20698
rect 12371 20646 12383 20698
rect 12445 20646 12447 20698
rect 12285 20644 12309 20646
rect 12365 20644 12389 20646
rect 12445 20644 12469 20646
rect 12229 20624 12525 20644
rect 13004 20602 13032 20946
rect 12992 20596 13044 20602
rect 12992 20538 13044 20544
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11716 17785 11744 18226
rect 11702 17776 11758 17785
rect 11702 17711 11758 17720
rect 10888 13786 11008 13814
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10060 13326 10088 13670
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10060 12986 10088 13262
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10428 12918 10456 13262
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9784 11898 9812 12310
rect 9876 11898 9904 12650
rect 10428 12374 10456 12854
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7944 8906 7972 9386
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 8471 9276 8767 9296
rect 8527 9274 8551 9276
rect 8607 9274 8631 9276
rect 8687 9274 8711 9276
rect 8549 9222 8551 9274
rect 8613 9222 8625 9274
rect 8687 9222 8689 9274
rect 8527 9220 8551 9222
rect 8607 9220 8631 9222
rect 8687 9220 8711 9222
rect 8471 9200 8767 9220
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 9048 8294 9076 9318
rect 9140 9110 9168 9318
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8471 8188 8767 8208
rect 8527 8186 8551 8188
rect 8607 8186 8631 8188
rect 8687 8186 8711 8188
rect 8549 8134 8551 8186
rect 8613 8134 8625 8186
rect 8687 8134 8689 8186
rect 8527 8132 8551 8134
rect 8607 8132 8631 8134
rect 8687 8132 8711 8134
rect 8471 8112 8767 8132
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8404 7478 8432 7822
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 7932 7268 7984 7274
rect 7852 7228 7932 7256
rect 7748 7200 7800 7206
rect 7668 7160 7748 7188
rect 7748 7142 7800 7148
rect 7760 7002 7788 7142
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7852 5896 7880 7228
rect 7932 7210 7984 7216
rect 8404 6322 8432 7414
rect 9416 7410 9444 8774
rect 9508 8634 9536 8978
rect 9496 8628 9548 8634
rect 9548 8588 9628 8616
rect 9496 8570 9548 8576
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 8471 7100 8767 7120
rect 8527 7098 8551 7100
rect 8607 7098 8631 7100
rect 8687 7098 8711 7100
rect 8549 7046 8551 7098
rect 8613 7046 8625 7098
rect 8687 7046 8689 7098
rect 8527 7044 8551 7046
rect 8607 7044 8631 7046
rect 8687 7044 8711 7046
rect 8471 7024 8767 7044
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8864 6118 8892 6802
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8036 5914 8064 6054
rect 8471 6012 8767 6032
rect 8527 6010 8551 6012
rect 8607 6010 8631 6012
rect 8687 6010 8711 6012
rect 8549 5958 8551 6010
rect 8613 5958 8625 6010
rect 8687 5958 8689 6010
rect 8527 5956 8551 5958
rect 8607 5956 8631 5958
rect 8687 5956 8711 5958
rect 8471 5936 8767 5956
rect 8024 5908 8076 5914
rect 7852 5868 7972 5896
rect 7944 5778 7972 5868
rect 8024 5850 8076 5856
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7668 4758 7696 5510
rect 7852 5030 7880 5714
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7668 4282 7696 4694
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 6274 4111 6330 4120
rect 7300 4126 7420 4154
rect 7300 4078 7328 4126
rect 7288 4072 7340 4078
rect 7852 4049 7880 4966
rect 7944 4622 7972 5034
rect 8471 4924 8767 4944
rect 8527 4922 8551 4924
rect 8607 4922 8631 4924
rect 8687 4922 8711 4924
rect 8549 4870 8551 4922
rect 8613 4870 8625 4922
rect 8687 4870 8689 4922
rect 8527 4868 8551 4870
rect 8607 4868 8631 4870
rect 8687 4868 8711 4870
rect 8471 4848 8767 4868
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7944 4214 7972 4558
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7288 4014 7340 4020
rect 7838 4040 7894 4049
rect 7838 3975 7894 3984
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7576 3670 7604 3878
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6012 2514 6040 3470
rect 6380 3126 6408 3538
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6656 2990 6684 3062
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 5630 54 5856 82
rect 6366 96 6422 480
rect 5630 0 5686 54
rect 7024 82 7052 3334
rect 7576 3194 7604 3606
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7102 82 7158 480
rect 7024 54 7158 82
rect 7760 82 7788 3878
rect 8471 3836 8767 3856
rect 8527 3834 8551 3836
rect 8607 3834 8631 3836
rect 8687 3834 8711 3836
rect 8549 3782 8551 3834
rect 8613 3782 8625 3834
rect 8687 3782 8689 3834
rect 8527 3780 8551 3782
rect 8607 3780 8631 3782
rect 8687 3780 8711 3782
rect 8471 3760 8767 3780
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8220 2514 8248 2790
rect 8404 2650 8432 2790
rect 8471 2748 8767 2768
rect 8527 2746 8551 2748
rect 8607 2746 8631 2748
rect 8687 2746 8711 2748
rect 8549 2694 8551 2746
rect 8613 2694 8625 2746
rect 8687 2694 8689 2746
rect 8527 2692 8551 2694
rect 8607 2692 8631 2694
rect 8687 2692 8711 2694
rect 8471 2672 8767 2692
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 7838 82 7894 480
rect 7760 54 7894 82
rect 6366 0 6422 40
rect 7102 0 7158 54
rect 7838 0 7894 54
rect 8574 82 8630 480
rect 8864 82 8892 6054
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9140 5370 9168 5714
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 8956 4010 8984 4966
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 9416 2650 9444 4966
rect 9600 4154 9628 8588
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9692 8090 9720 8298
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9784 7546 9812 7822
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9968 7478 9996 8434
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 7886 10088 8230
rect 10704 7954 10732 11630
rect 10888 11626 10916 13786
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10888 10130 10916 11562
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 11716 8906 11744 17711
rect 12084 9042 12112 20198
rect 12229 19612 12525 19632
rect 12285 19610 12309 19612
rect 12365 19610 12389 19612
rect 12445 19610 12469 19612
rect 12307 19558 12309 19610
rect 12371 19558 12383 19610
rect 12445 19558 12447 19610
rect 12285 19556 12309 19558
rect 12365 19556 12389 19558
rect 12445 19556 12469 19558
rect 12229 19536 12525 19556
rect 12229 18524 12525 18544
rect 12285 18522 12309 18524
rect 12365 18522 12389 18524
rect 12445 18522 12469 18524
rect 12307 18470 12309 18522
rect 12371 18470 12383 18522
rect 12445 18470 12447 18522
rect 12285 18468 12309 18470
rect 12365 18468 12389 18470
rect 12445 18468 12469 18470
rect 12229 18448 12525 18468
rect 12229 17436 12525 17456
rect 12285 17434 12309 17436
rect 12365 17434 12389 17436
rect 12445 17434 12469 17436
rect 12307 17382 12309 17434
rect 12371 17382 12383 17434
rect 12445 17382 12447 17434
rect 12285 17380 12309 17382
rect 12365 17380 12389 17382
rect 12445 17380 12469 17382
rect 12229 17360 12525 17380
rect 12229 16348 12525 16368
rect 12285 16346 12309 16348
rect 12365 16346 12389 16348
rect 12445 16346 12469 16348
rect 12307 16294 12309 16346
rect 12371 16294 12383 16346
rect 12445 16294 12447 16346
rect 12285 16292 12309 16294
rect 12365 16292 12389 16294
rect 12445 16292 12469 16294
rect 12229 16272 12525 16292
rect 12229 15260 12525 15280
rect 12285 15258 12309 15260
rect 12365 15258 12389 15260
rect 12445 15258 12469 15260
rect 12307 15206 12309 15258
rect 12371 15206 12383 15258
rect 12445 15206 12447 15258
rect 12285 15204 12309 15206
rect 12365 15204 12389 15206
rect 12445 15204 12469 15206
rect 12229 15184 12525 15204
rect 13464 14618 13492 24262
rect 13542 24210 13598 24262
rect 14738 24290 14794 24690
rect 15934 24290 15990 24690
rect 17130 24290 17186 24690
rect 14738 24262 14872 24290
rect 14738 24210 14794 24262
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13924 20602 13952 20742
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 14108 20058 14136 21286
rect 14844 21078 14872 24262
rect 15672 24262 15990 24290
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15580 21486 15608 22034
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15016 21412 15068 21418
rect 15016 21354 15068 21360
rect 14832 21072 14884 21078
rect 14832 21014 14884 21020
rect 15028 20262 15056 21354
rect 15016 20256 15068 20262
rect 15016 20198 15068 20204
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 15028 19990 15056 20198
rect 15016 19984 15068 19990
rect 15016 19926 15068 19932
rect 15488 19514 15516 20198
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15672 19378 15700 24262
rect 15934 24210 15990 24262
rect 16776 24262 17186 24290
rect 15986 22332 16282 22352
rect 16042 22330 16066 22332
rect 16122 22330 16146 22332
rect 16202 22330 16226 22332
rect 16064 22278 16066 22330
rect 16128 22278 16140 22330
rect 16202 22278 16204 22330
rect 16042 22276 16066 22278
rect 16122 22276 16146 22278
rect 16202 22276 16226 22278
rect 15986 22256 16282 22276
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 15986 21244 16282 21264
rect 16042 21242 16066 21244
rect 16122 21242 16146 21244
rect 16202 21242 16226 21244
rect 16064 21190 16066 21242
rect 16128 21190 16140 21242
rect 16202 21190 16204 21242
rect 16042 21188 16066 21190
rect 16122 21188 16146 21190
rect 16202 21188 16226 21190
rect 15986 21168 16282 21188
rect 15986 20156 16282 20176
rect 16042 20154 16066 20156
rect 16122 20154 16146 20156
rect 16202 20154 16226 20156
rect 16064 20102 16066 20154
rect 16128 20102 16140 20154
rect 16202 20102 16204 20154
rect 16042 20100 16066 20102
rect 16122 20100 16146 20102
rect 16202 20100 16226 20102
rect 15986 20080 16282 20100
rect 16316 19990 16344 21286
rect 16408 21078 16436 21286
rect 16396 21072 16448 21078
rect 16396 21014 16448 21020
rect 16408 20602 16436 21014
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16592 20466 16620 20878
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16592 19854 16620 20402
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 15856 19514 15884 19790
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 14554 15464 14610 15473
rect 14554 15399 14610 15408
rect 14568 15162 14596 15399
rect 15028 15162 15056 19246
rect 15986 19068 16282 19088
rect 16042 19066 16066 19068
rect 16122 19066 16146 19068
rect 16202 19066 16226 19068
rect 16064 19014 16066 19066
rect 16128 19014 16140 19066
rect 16202 19014 16204 19066
rect 16042 19012 16066 19014
rect 16122 19012 16146 19014
rect 16202 19012 16226 19014
rect 15986 18992 16282 19012
rect 15986 17980 16282 18000
rect 16042 17978 16066 17980
rect 16122 17978 16146 17980
rect 16202 17978 16226 17980
rect 16064 17926 16066 17978
rect 16128 17926 16140 17978
rect 16202 17926 16204 17978
rect 16042 17924 16066 17926
rect 16122 17924 16146 17926
rect 16202 17924 16226 17926
rect 15986 17904 16282 17924
rect 15986 16892 16282 16912
rect 16042 16890 16066 16892
rect 16122 16890 16146 16892
rect 16202 16890 16226 16892
rect 16064 16838 16066 16890
rect 16128 16838 16140 16890
rect 16202 16838 16204 16890
rect 16042 16836 16066 16838
rect 16122 16836 16146 16838
rect 16202 16836 16226 16838
rect 15986 16816 16282 16836
rect 15986 15804 16282 15824
rect 16042 15802 16066 15804
rect 16122 15802 16146 15804
rect 16202 15802 16226 15804
rect 16064 15750 16066 15802
rect 16128 15750 16140 15802
rect 16202 15750 16204 15802
rect 16042 15748 16066 15750
rect 16122 15748 16146 15750
rect 16202 15748 16226 15750
rect 15986 15728 16282 15748
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 15856 14550 15884 14758
rect 15986 14716 16282 14736
rect 16042 14714 16066 14716
rect 16122 14714 16146 14716
rect 16202 14714 16226 14716
rect 16064 14662 16066 14714
rect 16128 14662 16140 14714
rect 16202 14662 16204 14714
rect 16042 14660 16066 14662
rect 16122 14660 16146 14662
rect 16202 14660 16226 14662
rect 15986 14640 16282 14660
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 12229 14172 12525 14192
rect 12285 14170 12309 14172
rect 12365 14170 12389 14172
rect 12445 14170 12469 14172
rect 12307 14118 12309 14170
rect 12371 14118 12383 14170
rect 12445 14118 12447 14170
rect 12285 14116 12309 14118
rect 12365 14116 12389 14118
rect 12445 14116 12469 14118
rect 12229 14096 12525 14116
rect 13648 14074 13676 14418
rect 15856 14074 15884 14486
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 13648 13394 13676 14010
rect 16684 13938 16712 14282
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16776 13814 16804 24262
rect 17130 24210 17186 24262
rect 18326 24290 18382 24690
rect 19522 24290 19578 24690
rect 20718 24290 20774 24690
rect 21914 24290 21970 24690
rect 18326 24262 18460 24290
rect 18326 24210 18382 24262
rect 18432 21690 18460 24262
rect 19260 24262 19578 24290
rect 18510 21992 18566 22001
rect 18510 21927 18566 21936
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18524 21010 18552 21927
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18524 20602 18552 20946
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 17040 20528 17092 20534
rect 17040 20470 17092 20476
rect 16948 19984 17000 19990
rect 16948 19926 17000 19932
rect 16960 19514 16988 19926
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16592 13786 16804 13814
rect 15986 13628 16282 13648
rect 16042 13626 16066 13628
rect 16122 13626 16146 13628
rect 16202 13626 16226 13628
rect 16064 13574 16066 13626
rect 16128 13574 16140 13626
rect 16202 13574 16204 13626
rect 16042 13572 16066 13574
rect 16122 13572 16146 13574
rect 16202 13572 16226 13574
rect 15986 13552 16282 13572
rect 16316 13530 16344 13738
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 12229 13084 12525 13104
rect 12285 13082 12309 13084
rect 12365 13082 12389 13084
rect 12445 13082 12469 13084
rect 12307 13030 12309 13082
rect 12371 13030 12383 13082
rect 12445 13030 12447 13082
rect 12285 13028 12309 13030
rect 12365 13028 12389 13030
rect 12445 13028 12469 13030
rect 12229 13008 12525 13028
rect 12622 12744 12678 12753
rect 12622 12679 12678 12688
rect 12229 11996 12525 12016
rect 12285 11994 12309 11996
rect 12365 11994 12389 11996
rect 12445 11994 12469 11996
rect 12307 11942 12309 11994
rect 12371 11942 12383 11994
rect 12445 11942 12447 11994
rect 12285 11940 12309 11942
rect 12365 11940 12389 11942
rect 12445 11940 12469 11942
rect 12229 11920 12525 11940
rect 12636 11898 12664 12679
rect 15672 12646 15700 13330
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 16486 12608 16542 12617
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 15672 11694 15700 12582
rect 15986 12540 16282 12560
rect 16486 12543 16542 12552
rect 16042 12538 16066 12540
rect 16122 12538 16146 12540
rect 16202 12538 16226 12540
rect 16064 12486 16066 12538
rect 16128 12486 16140 12538
rect 16202 12486 16204 12538
rect 16042 12484 16066 12486
rect 16122 12484 16146 12486
rect 16202 12484 16226 12486
rect 15986 12464 16282 12484
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 12636 11354 12664 11630
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12229 10908 12525 10928
rect 12285 10906 12309 10908
rect 12365 10906 12389 10908
rect 12445 10906 12469 10908
rect 12307 10854 12309 10906
rect 12371 10854 12383 10906
rect 12445 10854 12447 10906
rect 12285 10852 12309 10854
rect 12365 10852 12389 10854
rect 12445 10852 12469 10854
rect 12229 10832 12525 10852
rect 12912 10810 12940 11154
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10198 12480 10406
rect 12440 10192 12492 10198
rect 12440 10134 12492 10140
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12229 9820 12525 9840
rect 12285 9818 12309 9820
rect 12365 9818 12389 9820
rect 12445 9818 12469 9820
rect 12307 9766 12309 9818
rect 12371 9766 12383 9818
rect 12445 9766 12447 9818
rect 12285 9764 12309 9766
rect 12365 9764 12389 9766
rect 12445 9764 12469 9766
rect 12229 9744 12525 9764
rect 12820 9722 12848 10134
rect 12912 10062 12940 10746
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12912 9586 12940 9998
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14096 9444 14148 9450
rect 14096 9386 14148 9392
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 12084 8634 12112 8978
rect 14108 8974 14136 9386
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 12229 8732 12525 8752
rect 12285 8730 12309 8732
rect 12365 8730 12389 8732
rect 12445 8730 12469 8732
rect 12307 8678 12309 8730
rect 12371 8678 12383 8730
rect 12445 8678 12447 8730
rect 12285 8676 12309 8678
rect 12365 8676 12389 8678
rect 12445 8676 12469 8678
rect 12229 8656 12525 8676
rect 13464 8634 13492 8910
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 12636 7954 12664 8570
rect 14108 8498 14136 8910
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14108 8090 14136 8298
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 11716 7546 11744 7890
rect 12229 7644 12525 7664
rect 12285 7642 12309 7644
rect 12365 7642 12389 7644
rect 12445 7642 12469 7644
rect 12307 7590 12309 7642
rect 12371 7590 12383 7642
rect 12445 7590 12447 7642
rect 12285 7588 12309 7590
rect 12365 7588 12389 7590
rect 12445 7588 12469 7590
rect 12229 7568 12525 7588
rect 12636 7546 12664 7890
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 13004 7410 13032 7686
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 6934 11192 7142
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9784 5846 9812 6734
rect 11164 6458 11192 6870
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 12716 6792 12768 6798
rect 13096 6769 13124 6802
rect 12716 6734 12768 6740
rect 13082 6760 13138 6769
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9876 5914 9904 6054
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9784 5370 9812 5782
rect 11072 5710 11100 6122
rect 11716 5846 11744 6598
rect 12229 6556 12525 6576
rect 12285 6554 12309 6556
rect 12365 6554 12389 6556
rect 12445 6554 12469 6556
rect 12307 6502 12309 6554
rect 12371 6502 12383 6554
rect 12445 6502 12447 6554
rect 12285 6500 12309 6502
rect 12365 6500 12389 6502
rect 12445 6500 12469 6502
rect 12229 6480 12525 6500
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 5370 11100 5646
rect 11716 5370 11744 5782
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12229 5468 12525 5488
rect 12285 5466 12309 5468
rect 12365 5466 12389 5468
rect 12445 5466 12469 5468
rect 12307 5414 12309 5466
rect 12371 5414 12383 5466
rect 12445 5414 12447 5466
rect 12285 5412 12309 5414
rect 12365 5412 12389 5414
rect 12445 5412 12469 5414
rect 12229 5392 12525 5412
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 12636 5234 12664 5510
rect 12728 5234 12756 6734
rect 13082 6695 13138 6704
rect 13096 6458 13124 6695
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13096 5778 13124 6394
rect 13464 6322 13492 6598
rect 13648 6322 13676 7210
rect 14568 6866 14596 9454
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 14568 6118 14596 6802
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 13096 5370 13124 5714
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 10428 4758 10456 5170
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10704 4826 10732 4966
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9784 4282 9812 4558
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9600 4126 9720 4154
rect 9692 4060 9720 4126
rect 9600 4032 9720 4060
rect 9600 3505 9628 4032
rect 10428 3670 10456 4694
rect 10704 4078 10732 4762
rect 12728 4758 12756 5170
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11992 4282 12020 4558
rect 12229 4380 12525 4400
rect 12285 4378 12309 4380
rect 12365 4378 12389 4380
rect 12445 4378 12469 4380
rect 12307 4326 12309 4378
rect 12371 4326 12383 4378
rect 12445 4326 12447 4378
rect 12285 4324 12309 4326
rect 12365 4324 12389 4326
rect 12445 4324 12469 4326
rect 12229 4304 12525 4324
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 11256 3602 11284 3878
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10048 3528 10100 3534
rect 9586 3496 9642 3505
rect 10048 3470 10100 3476
rect 9586 3431 9642 3440
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 8574 54 8892 82
rect 9402 82 9458 480
rect 9600 82 9628 3431
rect 10060 3194 10088 3470
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 11256 3108 11284 3538
rect 11336 3120 11388 3126
rect 11256 3080 11336 3108
rect 11336 3062 11388 3068
rect 10140 2916 10192 2922
rect 10140 2858 10192 2864
rect 10232 2916 10284 2922
rect 10232 2858 10284 2864
rect 10152 2582 10180 2858
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 10152 2446 10180 2518
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10244 2009 10272 2858
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10230 2000 10286 2009
rect 10230 1935 10286 1944
rect 9402 54 9628 82
rect 10138 82 10194 480
rect 10244 82 10272 1935
rect 10138 54 10272 82
rect 10874 82 10930 480
rect 10980 82 11008 2790
rect 10874 54 11008 82
rect 11610 82 11666 480
rect 11716 82 11744 4150
rect 12728 4146 12756 4694
rect 14462 4176 14518 4185
rect 12716 4140 12768 4146
rect 14462 4111 14464 4120
rect 12716 4082 12768 4088
rect 14516 4111 14518 4120
rect 14464 4082 14516 4088
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11992 2922 12020 3538
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 11610 54 11744 82
rect 12084 82 12112 3334
rect 12229 3292 12525 3312
rect 12285 3290 12309 3292
rect 12365 3290 12389 3292
rect 12445 3290 12469 3292
rect 12307 3238 12309 3290
rect 12371 3238 12383 3290
rect 12445 3238 12447 3290
rect 12285 3236 12309 3238
rect 12365 3236 12389 3238
rect 12445 3236 12469 3238
rect 12229 3216 12525 3236
rect 12636 3058 12664 3402
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12636 2650 12664 2994
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12229 2204 12525 2224
rect 12285 2202 12309 2204
rect 12365 2202 12389 2204
rect 12445 2202 12469 2204
rect 12307 2150 12309 2202
rect 12371 2150 12383 2202
rect 12445 2150 12447 2202
rect 12285 2148 12309 2150
rect 12365 2148 12389 2150
rect 12445 2148 12469 2150
rect 12229 2128 12525 2148
rect 12346 82 12402 480
rect 12820 134 12848 3334
rect 13004 3194 13032 3334
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13188 3058 13216 3946
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 13464 3194 13492 3538
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 13464 2582 13492 2858
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13176 2372 13228 2378
rect 13176 2314 13228 2320
rect 12084 54 12402 82
rect 12808 128 12860 134
rect 12808 70 12860 76
rect 13082 82 13138 480
rect 13188 82 13216 2314
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 8574 0 8630 54
rect 9402 0 9458 54
rect 10138 0 10194 54
rect 10874 0 10930 54
rect 11610 0 11666 54
rect 12346 0 12402 54
rect 13082 54 13216 82
rect 13832 82 13860 2246
rect 13910 82 13966 480
rect 14292 105 14320 2246
rect 13832 54 13966 82
rect 13082 0 13138 54
rect 13910 0 13966 54
rect 14278 96 14334 105
rect 14568 82 14596 6054
rect 14922 3496 14978 3505
rect 14922 3431 14978 3440
rect 14936 3126 14964 3431
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 14936 2990 14964 3062
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14646 82 14702 480
rect 14568 54 14702 82
rect 15304 82 15332 11630
rect 15986 11452 16282 11472
rect 16042 11450 16066 11452
rect 16122 11450 16146 11452
rect 16202 11450 16226 11452
rect 16064 11398 16066 11450
rect 16128 11398 16140 11450
rect 16202 11398 16204 11450
rect 16042 11396 16066 11398
rect 16122 11396 16146 11398
rect 16202 11396 16226 11398
rect 15986 11376 16282 11396
rect 16316 10810 16344 11630
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16408 11286 16436 11494
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16408 10742 16436 11222
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 15986 10364 16282 10384
rect 16042 10362 16066 10364
rect 16122 10362 16146 10364
rect 16202 10362 16226 10364
rect 16064 10310 16066 10362
rect 16128 10310 16140 10362
rect 16202 10310 16204 10362
rect 16042 10308 16066 10310
rect 16122 10308 16146 10310
rect 16202 10308 16226 10310
rect 15986 10288 16282 10308
rect 15986 9276 16282 9296
rect 16042 9274 16066 9276
rect 16122 9274 16146 9276
rect 16202 9274 16226 9276
rect 16064 9222 16066 9274
rect 16128 9222 16140 9274
rect 16202 9222 16204 9274
rect 16042 9220 16066 9222
rect 16122 9220 16146 9222
rect 16202 9220 16226 9222
rect 15986 9200 16282 9220
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 15986 8188 16282 8208
rect 16042 8186 16066 8188
rect 16122 8186 16146 8188
rect 16202 8186 16226 8188
rect 16064 8134 16066 8186
rect 16128 8134 16140 8186
rect 16202 8134 16204 8186
rect 16042 8132 16066 8134
rect 16122 8132 16146 8134
rect 16202 8132 16226 8134
rect 15986 8112 16282 8132
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15580 7206 15608 7890
rect 16408 7750 16436 8230
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15396 4758 15424 4966
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15396 4282 15424 4694
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15580 4154 15608 7142
rect 15986 7100 16282 7120
rect 16042 7098 16066 7100
rect 16122 7098 16146 7100
rect 16202 7098 16226 7100
rect 16064 7046 16066 7098
rect 16128 7046 16140 7098
rect 16202 7046 16204 7098
rect 16042 7044 16066 7046
rect 16122 7044 16146 7046
rect 16202 7044 16226 7046
rect 15986 7024 16282 7044
rect 16408 7002 16436 7686
rect 16500 7546 16528 12543
rect 16592 8242 16620 13786
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16960 10674 16988 11018
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 9110 16712 9318
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16684 8634 16712 9046
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16592 8214 16712 8242
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16500 7342 16528 7482
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16500 6118 16528 6802
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 15986 6012 16282 6032
rect 16042 6010 16066 6012
rect 16122 6010 16146 6012
rect 16202 6010 16226 6012
rect 16064 5958 16066 6010
rect 16128 5958 16140 6010
rect 16202 5958 16204 6010
rect 16042 5956 16066 5958
rect 16122 5956 16146 5958
rect 16202 5956 16226 5958
rect 15986 5936 16282 5956
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15672 5234 15700 5510
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 15986 4924 16282 4944
rect 16042 4922 16066 4924
rect 16122 4922 16146 4924
rect 16202 4922 16226 4924
rect 16064 4870 16066 4922
rect 16128 4870 16140 4922
rect 16202 4870 16204 4922
rect 16042 4868 16066 4870
rect 16122 4868 16146 4870
rect 16202 4868 16226 4870
rect 15986 4848 16282 4868
rect 16316 4758 16344 5034
rect 15752 4752 15804 4758
rect 15752 4694 15804 4700
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 15580 4126 15700 4154
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15396 3194 15424 3470
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15382 82 15438 480
rect 15304 54 15438 82
rect 15672 82 15700 4126
rect 15764 4010 15792 4694
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 15752 4004 15804 4010
rect 15752 3946 15804 3952
rect 15986 3836 16282 3856
rect 16042 3834 16066 3836
rect 16122 3834 16146 3836
rect 16202 3834 16226 3836
rect 16064 3782 16066 3834
rect 16128 3782 16140 3834
rect 16202 3782 16204 3834
rect 16042 3780 16066 3782
rect 16122 3780 16146 3782
rect 16202 3780 16226 3782
rect 15986 3760 16282 3780
rect 15986 2748 16282 2768
rect 16042 2746 16066 2748
rect 16122 2746 16146 2748
rect 16202 2746 16226 2748
rect 16064 2694 16066 2746
rect 16128 2694 16140 2746
rect 16202 2694 16204 2746
rect 16042 2692 16066 2694
rect 16122 2692 16146 2694
rect 16202 2692 16226 2694
rect 15986 2672 16282 2692
rect 16316 2650 16344 4422
rect 16500 3641 16528 6054
rect 16486 3632 16542 3641
rect 16486 3567 16542 3576
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 16500 2514 16528 3567
rect 16488 2508 16540 2514
rect 16488 2450 16540 2456
rect 16118 82 16174 480
rect 15672 54 16174 82
rect 16592 82 16620 7414
rect 16684 5778 16712 8214
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16684 5370 16712 5714
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16868 4010 16896 4490
rect 17052 4154 17080 20470
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 17880 19514 17908 19926
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18432 17785 18460 19314
rect 18418 17776 18474 17785
rect 18418 17711 18474 17720
rect 19260 16794 19288 24262
rect 19522 24210 19578 24262
rect 20272 24262 20774 24290
rect 20166 23352 20222 23361
rect 20166 23287 20222 23296
rect 20180 22098 20208 23287
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 19352 20602 19380 21014
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19352 19174 19380 19790
rect 19536 19378 19564 20742
rect 19628 20466 19656 21830
rect 19744 21788 20040 21808
rect 19800 21786 19824 21788
rect 19880 21786 19904 21788
rect 19960 21786 19984 21788
rect 19822 21734 19824 21786
rect 19886 21734 19898 21786
rect 19960 21734 19962 21786
rect 19800 21732 19824 21734
rect 19880 21732 19904 21734
rect 19960 21732 19984 21734
rect 19744 21712 20040 21732
rect 20180 21690 20208 22034
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20272 21622 20300 24262
rect 20718 24210 20774 24262
rect 21560 24262 21970 24290
rect 21560 21690 21588 24262
rect 21914 24210 21970 24262
rect 21548 21684 21600 21690
rect 21548 21626 21600 21632
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19720 21078 19748 21286
rect 19708 21072 19760 21078
rect 19708 21014 19760 21020
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 19744 20700 20040 20720
rect 19800 20698 19824 20700
rect 19880 20698 19904 20700
rect 19960 20698 19984 20700
rect 19822 20646 19824 20698
rect 19886 20646 19898 20698
rect 19960 20646 19962 20698
rect 19800 20644 19824 20646
rect 19880 20644 19904 20646
rect 19960 20644 19984 20646
rect 19744 20624 20040 20644
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 20088 19990 20116 20878
rect 20350 20224 20406 20233
rect 20350 20159 20406 20168
rect 20076 19984 20128 19990
rect 20076 19926 20128 19932
rect 19744 19612 20040 19632
rect 19800 19610 19824 19612
rect 19880 19610 19904 19612
rect 19960 19610 19984 19612
rect 19822 19558 19824 19610
rect 19886 19558 19898 19610
rect 19960 19558 19962 19610
rect 19800 19556 19824 19558
rect 19880 19556 19904 19558
rect 19960 19556 19984 19558
rect 19744 19536 20040 19556
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19432 19236 19484 19242
rect 19432 19178 19484 19184
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19352 18970 19380 19110
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19444 17082 19472 19178
rect 19536 18902 19564 19314
rect 19524 18896 19576 18902
rect 19524 18838 19576 18844
rect 20364 18834 20392 20159
rect 22098 19272 22154 19281
rect 22098 19207 22154 19216
rect 20352 18828 20404 18834
rect 20352 18770 20404 18776
rect 19744 18524 20040 18544
rect 19800 18522 19824 18524
rect 19880 18522 19904 18524
rect 19960 18522 19984 18524
rect 19822 18470 19824 18522
rect 19886 18470 19898 18522
rect 19960 18470 19962 18522
rect 19800 18468 19824 18470
rect 19880 18468 19904 18470
rect 19960 18468 19984 18470
rect 19744 18448 20040 18468
rect 20364 18426 20392 18770
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 22112 18193 22140 19207
rect 22098 18184 22154 18193
rect 22098 18119 22154 18128
rect 19744 17436 20040 17456
rect 19800 17434 19824 17436
rect 19880 17434 19904 17436
rect 19960 17434 19984 17436
rect 19822 17382 19824 17434
rect 19886 17382 19898 17434
rect 19960 17382 19962 17434
rect 19800 17380 19824 17382
rect 19880 17380 19904 17382
rect 19960 17380 19984 17382
rect 19744 17360 20040 17380
rect 19798 17232 19854 17241
rect 19798 17167 19854 17176
rect 19522 17096 19578 17105
rect 19444 17054 19522 17082
rect 19522 17031 19578 17040
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19444 15910 19472 16594
rect 19536 16114 19564 17031
rect 19812 16794 19840 17167
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19744 16348 20040 16368
rect 19800 16346 19824 16348
rect 19880 16346 19904 16348
rect 19960 16346 19984 16348
rect 19822 16294 19824 16346
rect 19886 16294 19898 16346
rect 19960 16294 19962 16346
rect 19800 16292 19824 16294
rect 19880 16292 19904 16294
rect 19960 16292 19984 16294
rect 19744 16272 20040 16292
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19524 15972 19576 15978
rect 19524 15914 19576 15920
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19062 15600 19118 15609
rect 19062 15535 19118 15544
rect 18236 14000 18288 14006
rect 18236 13942 18288 13948
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 10810 18092 11494
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17144 8906 17172 9318
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17144 8498 17172 8842
rect 18156 8498 18184 8910
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17788 8090 17816 8230
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17880 7546 17908 7890
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18248 7392 18276 13942
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 10062 18736 11494
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18800 10674 18828 11086
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18432 9722 18460 9998
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18708 9654 18736 9998
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18800 9042 18828 10610
rect 19076 9704 19104 15535
rect 19444 15162 19472 15846
rect 19536 15638 19564 15914
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 19744 15260 20040 15280
rect 19800 15258 19824 15260
rect 19880 15258 19904 15260
rect 19960 15258 19984 15260
rect 19822 15206 19824 15258
rect 19886 15206 19898 15258
rect 19960 15206 19962 15258
rect 19800 15204 19824 15206
rect 19880 15204 19904 15206
rect 19960 15204 19984 15206
rect 19744 15184 20040 15204
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 20088 14890 20116 15506
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19744 14172 20040 14192
rect 19800 14170 19824 14172
rect 19880 14170 19904 14172
rect 19960 14170 19984 14172
rect 19822 14118 19824 14170
rect 19886 14118 19898 14170
rect 19960 14118 19962 14170
rect 19800 14116 19824 14118
rect 19880 14116 19904 14118
rect 19960 14116 19984 14118
rect 19744 14096 20040 14116
rect 20272 14006 20300 14894
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20260 14000 20312 14006
rect 20260 13942 20312 13948
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19168 13802 19196 13874
rect 19156 13796 19208 13802
rect 19156 13738 19208 13744
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19444 12850 19472 13738
rect 19744 13084 20040 13104
rect 19800 13082 19824 13084
rect 19880 13082 19904 13084
rect 19960 13082 19984 13084
rect 19822 13030 19824 13082
rect 19886 13030 19898 13082
rect 19960 13030 19962 13082
rect 19800 13028 19824 13030
rect 19880 13028 19904 13030
rect 19960 13028 19984 13030
rect 19744 13008 20040 13028
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19444 12442 19472 12650
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19616 12300 19668 12306
rect 19616 12242 19668 12248
rect 19628 11558 19656 12242
rect 19744 11996 20040 12016
rect 19800 11994 19824 11996
rect 19880 11994 19904 11996
rect 19960 11994 19984 11996
rect 19822 11942 19824 11994
rect 19886 11942 19898 11994
rect 19960 11942 19962 11994
rect 19800 11940 19824 11942
rect 19880 11940 19904 11942
rect 19960 11940 19984 11942
rect 19744 11920 20040 11940
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19616 11552 19668 11558
rect 20628 11552 20680 11558
rect 19616 11494 19668 11500
rect 19798 11520 19854 11529
rect 19536 11218 19564 11494
rect 20628 11494 20680 11500
rect 19798 11455 19854 11464
rect 19812 11354 19840 11455
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19536 10810 19564 11154
rect 19744 10908 20040 10928
rect 19800 10906 19824 10908
rect 19880 10906 19904 10908
rect 19960 10906 19984 10908
rect 19822 10854 19824 10906
rect 19886 10854 19898 10906
rect 19960 10854 19962 10906
rect 19800 10852 19824 10854
rect 19880 10852 19904 10854
rect 19960 10852 19984 10854
rect 19744 10832 20040 10852
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19744 9820 20040 9840
rect 19800 9818 19824 9820
rect 19880 9818 19904 9820
rect 19960 9818 19984 9820
rect 19822 9766 19824 9818
rect 19886 9766 19898 9818
rect 19960 9766 19962 9818
rect 19800 9764 19824 9766
rect 19880 9764 19904 9766
rect 19960 9764 19984 9766
rect 19744 9744 20040 9764
rect 19156 9716 19208 9722
rect 19076 9676 19156 9704
rect 19156 9658 19208 9664
rect 20088 9178 20116 10542
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19444 8634 19472 8978
rect 19744 8732 20040 8752
rect 19800 8730 19824 8732
rect 19880 8730 19904 8732
rect 19960 8730 19984 8732
rect 19822 8678 19824 8730
rect 19886 8678 19898 8730
rect 19960 8678 19962 8730
rect 19800 8676 19824 8678
rect 19880 8676 19904 8678
rect 19960 8676 19984 8678
rect 19744 8656 20040 8676
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 18880 7880 18932 7886
rect 18694 7848 18750 7857
rect 18880 7822 18932 7828
rect 18694 7783 18750 7792
rect 18708 7546 18736 7783
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18328 7404 18380 7410
rect 18248 7364 18328 7392
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17696 6458 17724 6734
rect 18248 6730 18276 7364
rect 18328 7346 18380 7352
rect 18892 7274 18920 7822
rect 18880 7268 18932 7274
rect 18880 7210 18932 7216
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18616 5166 18644 6054
rect 18800 5681 18828 7142
rect 18892 7002 18920 7210
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 19076 6458 19104 8230
rect 19168 7886 19196 8434
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 6934 19288 7686
rect 19744 7644 20040 7664
rect 19800 7642 19824 7644
rect 19880 7642 19904 7644
rect 19960 7642 19984 7644
rect 19822 7590 19824 7642
rect 19886 7590 19898 7642
rect 19960 7590 19962 7642
rect 19800 7588 19824 7590
rect 19880 7588 19904 7590
rect 19960 7588 19984 7590
rect 19744 7568 20040 7588
rect 19248 6928 19300 6934
rect 19248 6870 19300 6876
rect 19260 6458 19288 6870
rect 19432 6724 19484 6730
rect 19432 6666 19484 6672
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19444 6322 19472 6666
rect 19744 6556 20040 6576
rect 19800 6554 19824 6556
rect 19880 6554 19904 6556
rect 19960 6554 19984 6556
rect 19822 6502 19824 6554
rect 19886 6502 19898 6554
rect 19960 6502 19962 6554
rect 19800 6500 19824 6502
rect 19880 6500 19904 6502
rect 19960 6500 19984 6502
rect 19744 6480 20040 6500
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19156 6180 19208 6186
rect 19156 6122 19208 6128
rect 18972 5704 19024 5710
rect 18786 5672 18842 5681
rect 18972 5646 19024 5652
rect 18786 5607 18842 5616
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18800 4758 18828 5607
rect 18984 5370 19012 5646
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 19168 5234 19196 6122
rect 19444 5710 19472 6258
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19744 5468 20040 5488
rect 19800 5466 19824 5468
rect 19880 5466 19904 5468
rect 19960 5466 19984 5468
rect 19822 5414 19824 5466
rect 19886 5414 19898 5466
rect 19960 5414 19962 5466
rect 19800 5412 19824 5414
rect 19880 5412 19904 5414
rect 19960 5412 19984 5414
rect 19744 5392 20040 5412
rect 20166 5400 20222 5409
rect 20166 5335 20222 5344
rect 20180 5302 20208 5335
rect 20168 5296 20220 5302
rect 20168 5238 20220 5244
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 18788 4752 18840 4758
rect 18788 4694 18840 4700
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19352 4282 19380 4558
rect 19744 4380 20040 4400
rect 19800 4378 19824 4380
rect 19880 4378 19904 4380
rect 19960 4378 19984 4380
rect 19822 4326 19824 4378
rect 19886 4326 19898 4378
rect 19960 4326 19962 4378
rect 19800 4324 19824 4326
rect 19880 4324 19904 4326
rect 19960 4324 19984 4326
rect 19744 4304 20040 4324
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 16960 4126 17080 4154
rect 20260 4140 20312 4146
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16868 3058 16896 3946
rect 16960 3534 16988 4126
rect 20260 4082 20312 4088
rect 20074 4040 20130 4049
rect 20074 3975 20130 3984
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 16960 3194 16988 3470
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17236 3126 17264 3470
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 18432 3058 18460 3470
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17328 2650 17356 2790
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 18524 2582 18552 3878
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 18512 2576 18564 2582
rect 18512 2518 18564 2524
rect 18800 2446 18828 2858
rect 19536 2854 19564 3538
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19628 3126 19656 3334
rect 19744 3292 20040 3312
rect 19800 3290 19824 3292
rect 19880 3290 19904 3292
rect 19960 3290 19984 3292
rect 19822 3238 19824 3290
rect 19886 3238 19898 3290
rect 19960 3238 19962 3290
rect 19800 3236 19824 3238
rect 19880 3236 19904 3238
rect 19960 3236 19984 3238
rect 19744 3216 20040 3236
rect 19616 3120 19668 3126
rect 19616 3062 19668 3068
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 19628 2650 19656 3062
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 17316 2372 17368 2378
rect 17316 2314 17368 2320
rect 16854 82 16910 480
rect 16592 54 16910 82
rect 17328 82 17356 2314
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 17590 82 17646 480
rect 17328 54 17646 82
rect 14278 31 14334 40
rect 14646 0 14702 54
rect 15382 0 15438 54
rect 16118 0 16174 54
rect 16854 0 16910 54
rect 17590 0 17646 54
rect 18418 128 18474 480
rect 18418 76 18420 128
rect 18472 76 18474 128
rect 18418 0 18474 76
rect 19154 82 19210 480
rect 19444 82 19472 2246
rect 19744 2204 20040 2224
rect 19800 2202 19824 2204
rect 19880 2202 19904 2204
rect 19960 2202 19984 2204
rect 19822 2150 19824 2202
rect 19886 2150 19898 2202
rect 19960 2150 19962 2202
rect 19800 2148 19824 2150
rect 19880 2148 19904 2150
rect 19960 2148 19984 2150
rect 19744 2128 20040 2148
rect 19154 54 19472 82
rect 19890 82 19946 480
rect 20088 82 20116 3975
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20180 1329 20208 3878
rect 20166 1320 20222 1329
rect 20166 1255 20222 1264
rect 19890 54 20116 82
rect 20272 82 20300 4082
rect 20640 2825 20668 11494
rect 20626 2816 20682 2825
rect 20626 2751 20682 2760
rect 20626 82 20682 480
rect 20732 134 20760 14826
rect 22100 10736 22152 10742
rect 22100 10678 22152 10684
rect 22112 10033 22140 10678
rect 22098 10024 22154 10033
rect 22098 9959 22154 9968
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 20272 54 20682 82
rect 20720 128 20772 134
rect 20720 70 20772 76
rect 21362 128 21418 480
rect 21362 76 21364 128
rect 21416 76 21418 128
rect 19154 0 19210 54
rect 19890 0 19946 54
rect 20626 0 20682 54
rect 21362 0 21418 76
rect 21744 82 21772 2790
rect 22098 82 22154 480
rect 21744 54 22154 82
rect 22098 0 22154 54
<< via2 >>
rect 18 23976 74 24032
rect 110 22616 166 22672
rect 1582 20712 1638 20768
rect 1582 19352 1638 19408
rect 110 10240 166 10296
rect 1858 8336 1914 8392
rect 2502 6976 2558 7032
rect 1214 5616 1270 5672
rect 4713 21786 4769 21788
rect 4793 21786 4849 21788
rect 4873 21786 4929 21788
rect 4953 21786 5009 21788
rect 4713 21734 4739 21786
rect 4739 21734 4769 21786
rect 4793 21734 4803 21786
rect 4803 21734 4849 21786
rect 4873 21734 4919 21786
rect 4919 21734 4929 21786
rect 4953 21734 4983 21786
rect 4983 21734 5009 21786
rect 4713 21732 4769 21734
rect 4793 21732 4849 21734
rect 4873 21732 4929 21734
rect 4953 21732 5009 21734
rect 4713 20698 4769 20700
rect 4793 20698 4849 20700
rect 4873 20698 4929 20700
rect 4953 20698 5009 20700
rect 4713 20646 4739 20698
rect 4739 20646 4769 20698
rect 4793 20646 4803 20698
rect 4803 20646 4849 20698
rect 4873 20646 4919 20698
rect 4919 20646 4929 20698
rect 4953 20646 4983 20698
rect 4983 20646 5009 20698
rect 4713 20644 4769 20646
rect 4793 20644 4849 20646
rect 4873 20644 4929 20646
rect 4953 20644 5009 20646
rect 4713 19610 4769 19612
rect 4793 19610 4849 19612
rect 4873 19610 4929 19612
rect 4953 19610 5009 19612
rect 4713 19558 4739 19610
rect 4739 19558 4769 19610
rect 4793 19558 4803 19610
rect 4803 19558 4849 19610
rect 4873 19558 4919 19610
rect 4919 19558 4929 19610
rect 4953 19558 4983 19610
rect 4983 19558 5009 19610
rect 4713 19556 4769 19558
rect 4793 19556 4849 19558
rect 4873 19556 4929 19558
rect 4953 19556 5009 19558
rect 4713 18522 4769 18524
rect 4793 18522 4849 18524
rect 4873 18522 4929 18524
rect 4953 18522 5009 18524
rect 4713 18470 4739 18522
rect 4739 18470 4769 18522
rect 4793 18470 4803 18522
rect 4803 18470 4849 18522
rect 4873 18470 4919 18522
rect 4919 18470 4929 18522
rect 4953 18470 4983 18522
rect 4983 18470 5009 18522
rect 4713 18468 4769 18470
rect 4793 18468 4849 18470
rect 4873 18468 4929 18470
rect 4953 18468 5009 18470
rect 4713 17434 4769 17436
rect 4793 17434 4849 17436
rect 4873 17434 4929 17436
rect 4953 17434 5009 17436
rect 4713 17382 4739 17434
rect 4739 17382 4769 17434
rect 4793 17382 4803 17434
rect 4803 17382 4849 17434
rect 4873 17382 4919 17434
rect 4919 17382 4929 17434
rect 4953 17382 4983 17434
rect 4983 17382 5009 17434
rect 4713 17380 4769 17382
rect 4793 17380 4849 17382
rect 4873 17380 4929 17382
rect 4953 17380 5009 17382
rect 5354 16632 5410 16688
rect 4713 16346 4769 16348
rect 4793 16346 4849 16348
rect 4873 16346 4929 16348
rect 4953 16346 5009 16348
rect 4713 16294 4739 16346
rect 4739 16294 4769 16346
rect 4793 16294 4803 16346
rect 4803 16294 4849 16346
rect 4873 16294 4919 16346
rect 4919 16294 4929 16346
rect 4953 16294 4983 16346
rect 4983 16294 5009 16346
rect 4713 16292 4769 16294
rect 4793 16292 4849 16294
rect 4873 16292 4929 16294
rect 4953 16292 5009 16294
rect 4713 15258 4769 15260
rect 4793 15258 4849 15260
rect 4873 15258 4929 15260
rect 4953 15258 5009 15260
rect 4713 15206 4739 15258
rect 4739 15206 4769 15258
rect 4793 15206 4803 15258
rect 4803 15206 4849 15258
rect 4873 15206 4919 15258
rect 4919 15206 4929 15258
rect 4953 15206 4983 15258
rect 4983 15206 5009 15258
rect 4713 15204 4769 15206
rect 4793 15204 4849 15206
rect 4873 15204 4929 15206
rect 4953 15204 5009 15206
rect 4713 14170 4769 14172
rect 4793 14170 4849 14172
rect 4873 14170 4929 14172
rect 4953 14170 5009 14172
rect 4713 14118 4739 14170
rect 4739 14118 4769 14170
rect 4793 14118 4803 14170
rect 4803 14118 4849 14170
rect 4873 14118 4919 14170
rect 4919 14118 4929 14170
rect 4953 14118 4983 14170
rect 4983 14118 5009 14170
rect 4713 14116 4769 14118
rect 4793 14116 4849 14118
rect 4873 14116 4929 14118
rect 4953 14116 5009 14118
rect 4713 13082 4769 13084
rect 4793 13082 4849 13084
rect 4873 13082 4929 13084
rect 4953 13082 5009 13084
rect 4713 13030 4739 13082
rect 4739 13030 4769 13082
rect 4793 13030 4803 13082
rect 4803 13030 4849 13082
rect 4873 13030 4919 13082
rect 4919 13030 4929 13082
rect 4953 13030 4983 13082
rect 4983 13030 5009 13082
rect 4713 13028 4769 13030
rect 4793 13028 4849 13030
rect 4873 13028 4929 13030
rect 4953 13028 5009 13030
rect 4713 11994 4769 11996
rect 4793 11994 4849 11996
rect 4873 11994 4929 11996
rect 4953 11994 5009 11996
rect 4713 11942 4739 11994
rect 4739 11942 4769 11994
rect 4793 11942 4803 11994
rect 4803 11942 4849 11994
rect 4873 11942 4919 11994
rect 4919 11942 4929 11994
rect 4953 11942 4983 11994
rect 4983 11942 5009 11994
rect 4713 11940 4769 11942
rect 4793 11940 4849 11942
rect 4873 11940 4929 11942
rect 4953 11940 5009 11942
rect 4713 10906 4769 10908
rect 4793 10906 4849 10908
rect 4873 10906 4929 10908
rect 4953 10906 5009 10908
rect 4713 10854 4739 10906
rect 4739 10854 4769 10906
rect 4793 10854 4803 10906
rect 4803 10854 4849 10906
rect 4873 10854 4919 10906
rect 4919 10854 4929 10906
rect 4953 10854 4983 10906
rect 4983 10854 5009 10906
rect 4713 10852 4769 10854
rect 4793 10852 4849 10854
rect 4873 10852 4929 10854
rect 4953 10852 5009 10854
rect 4713 9818 4769 9820
rect 4793 9818 4849 9820
rect 4873 9818 4929 9820
rect 4953 9818 5009 9820
rect 4713 9766 4739 9818
rect 4739 9766 4769 9818
rect 4793 9766 4803 9818
rect 4803 9766 4849 9818
rect 4873 9766 4919 9818
rect 4919 9766 4929 9818
rect 4953 9766 4983 9818
rect 4983 9766 5009 9818
rect 4713 9764 4769 9766
rect 4793 9764 4849 9766
rect 4873 9764 4929 9766
rect 4953 9764 5009 9766
rect 4713 8730 4769 8732
rect 4793 8730 4849 8732
rect 4873 8730 4929 8732
rect 4953 8730 5009 8732
rect 4713 8678 4739 8730
rect 4739 8678 4769 8730
rect 4793 8678 4803 8730
rect 4803 8678 4849 8730
rect 4873 8678 4919 8730
rect 4919 8678 4929 8730
rect 4953 8678 4983 8730
rect 4983 8678 5009 8730
rect 4713 8676 4769 8678
rect 4793 8676 4849 8678
rect 4873 8676 4929 8678
rect 4953 8676 5009 8678
rect 4713 7642 4769 7644
rect 4793 7642 4849 7644
rect 4873 7642 4929 7644
rect 4953 7642 5009 7644
rect 4713 7590 4739 7642
rect 4739 7590 4769 7642
rect 4793 7590 4803 7642
rect 4803 7590 4849 7642
rect 4873 7590 4919 7642
rect 4919 7590 4929 7642
rect 4953 7590 4983 7642
rect 4983 7590 5009 7642
rect 4713 7588 4769 7590
rect 4793 7588 4849 7590
rect 4873 7588 4929 7590
rect 4953 7588 5009 7590
rect 4713 6554 4769 6556
rect 4793 6554 4849 6556
rect 4873 6554 4929 6556
rect 4953 6554 5009 6556
rect 4713 6502 4739 6554
rect 4739 6502 4769 6554
rect 4793 6502 4803 6554
rect 4803 6502 4849 6554
rect 4873 6502 4919 6554
rect 4919 6502 4929 6554
rect 4953 6502 4983 6554
rect 4983 6502 5009 6554
rect 4713 6500 4769 6502
rect 4793 6500 4849 6502
rect 4873 6500 4929 6502
rect 4953 6500 5009 6502
rect 3422 5616 3478 5672
rect 4713 5466 4769 5468
rect 4793 5466 4849 5468
rect 4873 5466 4929 5468
rect 4953 5466 5009 5468
rect 4713 5414 4739 5466
rect 4739 5414 4769 5466
rect 4793 5414 4803 5466
rect 4803 5414 4849 5466
rect 4873 5414 4919 5466
rect 4919 5414 4929 5466
rect 4953 5414 4983 5466
rect 4983 5414 5009 5466
rect 4713 5412 4769 5414
rect 4793 5412 4849 5414
rect 4873 5412 4929 5414
rect 4953 5412 5009 5414
rect 6274 17992 6330 18048
rect 7746 17040 7802 17096
rect 1858 4392 1914 4448
rect 4713 4378 4769 4380
rect 4793 4378 4849 4380
rect 4873 4378 4929 4380
rect 4953 4378 5009 4380
rect 4713 4326 4739 4378
rect 4739 4326 4769 4378
rect 4793 4326 4803 4378
rect 4803 4326 4849 4378
rect 4873 4326 4919 4378
rect 4919 4326 4929 4378
rect 4953 4326 4983 4378
rect 4983 4326 5009 4378
rect 4713 4324 4769 4326
rect 4793 4324 4849 4326
rect 4873 4324 4929 4326
rect 4953 4324 5009 4326
rect 5078 4120 5134 4176
rect 2502 1944 2558 2000
rect 4713 3290 4769 3292
rect 4793 3290 4849 3292
rect 4873 3290 4929 3292
rect 4953 3290 5009 3292
rect 4713 3238 4739 3290
rect 4739 3238 4769 3290
rect 4793 3238 4803 3290
rect 4803 3238 4849 3290
rect 4873 3238 4919 3290
rect 4919 3238 4929 3290
rect 4953 3238 4983 3290
rect 4983 3238 5009 3290
rect 4713 3236 4769 3238
rect 4793 3236 4849 3238
rect 4873 3236 4929 3238
rect 4953 3236 5009 3238
rect 4713 2202 4769 2204
rect 4793 2202 4849 2204
rect 4873 2202 4929 2204
rect 4953 2202 5009 2204
rect 4713 2150 4739 2202
rect 4739 2150 4769 2202
rect 4793 2150 4803 2202
rect 4803 2150 4849 2202
rect 4873 2150 4919 2202
rect 4919 2150 4929 2202
rect 4953 2150 4983 2202
rect 4983 2150 5009 2202
rect 4713 2148 4769 2150
rect 4793 2148 4849 2150
rect 4873 2148 4929 2150
rect 4953 2148 5009 2150
rect 6274 4120 6330 4176
rect 8471 22330 8527 22332
rect 8551 22330 8607 22332
rect 8631 22330 8687 22332
rect 8711 22330 8767 22332
rect 8471 22278 8497 22330
rect 8497 22278 8527 22330
rect 8551 22278 8561 22330
rect 8561 22278 8607 22330
rect 8631 22278 8677 22330
rect 8677 22278 8687 22330
rect 8711 22278 8741 22330
rect 8741 22278 8767 22330
rect 8471 22276 8527 22278
rect 8551 22276 8607 22278
rect 8631 22276 8687 22278
rect 8711 22276 8767 22278
rect 8471 21242 8527 21244
rect 8551 21242 8607 21244
rect 8631 21242 8687 21244
rect 8711 21242 8767 21244
rect 8471 21190 8497 21242
rect 8497 21190 8527 21242
rect 8551 21190 8561 21242
rect 8561 21190 8607 21242
rect 8631 21190 8677 21242
rect 8677 21190 8687 21242
rect 8711 21190 8741 21242
rect 8741 21190 8767 21242
rect 8471 21188 8527 21190
rect 8551 21188 8607 21190
rect 8631 21188 8687 21190
rect 8711 21188 8767 21190
rect 8471 20154 8527 20156
rect 8551 20154 8607 20156
rect 8631 20154 8687 20156
rect 8711 20154 8767 20156
rect 8471 20102 8497 20154
rect 8497 20102 8527 20154
rect 8551 20102 8561 20154
rect 8561 20102 8607 20154
rect 8631 20102 8677 20154
rect 8677 20102 8687 20154
rect 8711 20102 8741 20154
rect 8741 20102 8767 20154
rect 8471 20100 8527 20102
rect 8551 20100 8607 20102
rect 8631 20100 8687 20102
rect 8711 20100 8767 20102
rect 8471 19066 8527 19068
rect 8551 19066 8607 19068
rect 8631 19066 8687 19068
rect 8711 19066 8767 19068
rect 8471 19014 8497 19066
rect 8497 19014 8527 19066
rect 8551 19014 8561 19066
rect 8561 19014 8607 19066
rect 8631 19014 8677 19066
rect 8677 19014 8687 19066
rect 8711 19014 8741 19066
rect 8741 19014 8767 19066
rect 8471 19012 8527 19014
rect 8551 19012 8607 19014
rect 8631 19012 8687 19014
rect 8711 19012 8767 19014
rect 8850 18128 8906 18184
rect 8471 17978 8527 17980
rect 8551 17978 8607 17980
rect 8631 17978 8687 17980
rect 8711 17978 8767 17980
rect 8471 17926 8497 17978
rect 8497 17926 8527 17978
rect 8551 17926 8561 17978
rect 8561 17926 8607 17978
rect 8631 17926 8677 17978
rect 8677 17926 8687 17978
rect 8711 17926 8741 17978
rect 8741 17926 8767 17978
rect 8471 17924 8527 17926
rect 8551 17924 8607 17926
rect 8631 17924 8687 17926
rect 8711 17924 8767 17926
rect 8471 16890 8527 16892
rect 8551 16890 8607 16892
rect 8631 16890 8687 16892
rect 8711 16890 8767 16892
rect 8471 16838 8497 16890
rect 8497 16838 8527 16890
rect 8551 16838 8561 16890
rect 8561 16838 8607 16890
rect 8631 16838 8677 16890
rect 8677 16838 8687 16890
rect 8711 16838 8741 16890
rect 8741 16838 8767 16890
rect 8471 16836 8527 16838
rect 8551 16836 8607 16838
rect 8631 16836 8687 16838
rect 8711 16836 8767 16838
rect 8471 15802 8527 15804
rect 8551 15802 8607 15804
rect 8631 15802 8687 15804
rect 8711 15802 8767 15804
rect 8471 15750 8497 15802
rect 8497 15750 8527 15802
rect 8551 15750 8561 15802
rect 8561 15750 8607 15802
rect 8631 15750 8677 15802
rect 8677 15750 8687 15802
rect 8711 15750 8741 15802
rect 8741 15750 8767 15802
rect 8471 15748 8527 15750
rect 8551 15748 8607 15750
rect 8631 15748 8687 15750
rect 8711 15748 8767 15750
rect 9494 14864 9550 14920
rect 8471 14714 8527 14716
rect 8551 14714 8607 14716
rect 8631 14714 8687 14716
rect 8711 14714 8767 14716
rect 8471 14662 8497 14714
rect 8497 14662 8527 14714
rect 8551 14662 8561 14714
rect 8561 14662 8607 14714
rect 8631 14662 8677 14714
rect 8677 14662 8687 14714
rect 8711 14662 8741 14714
rect 8741 14662 8767 14714
rect 8471 14660 8527 14662
rect 8551 14660 8607 14662
rect 8631 14660 8687 14662
rect 8711 14660 8767 14662
rect 8471 13626 8527 13628
rect 8551 13626 8607 13628
rect 8631 13626 8687 13628
rect 8711 13626 8767 13628
rect 8471 13574 8497 13626
rect 8497 13574 8527 13626
rect 8551 13574 8561 13626
rect 8561 13574 8607 13626
rect 8631 13574 8677 13626
rect 8677 13574 8687 13626
rect 8711 13574 8741 13626
rect 8741 13574 8767 13626
rect 8471 13572 8527 13574
rect 8551 13572 8607 13574
rect 8631 13572 8687 13574
rect 8711 13572 8767 13574
rect 8471 12538 8527 12540
rect 8551 12538 8607 12540
rect 8631 12538 8687 12540
rect 8711 12538 8767 12540
rect 8471 12486 8497 12538
rect 8497 12486 8527 12538
rect 8551 12486 8561 12538
rect 8561 12486 8607 12538
rect 8631 12486 8677 12538
rect 8677 12486 8687 12538
rect 8711 12486 8741 12538
rect 8741 12486 8767 12538
rect 8471 12484 8527 12486
rect 8551 12484 8607 12486
rect 8631 12484 8687 12486
rect 8711 12484 8767 12486
rect 8471 11450 8527 11452
rect 8551 11450 8607 11452
rect 8631 11450 8687 11452
rect 8711 11450 8767 11452
rect 8471 11398 8497 11450
rect 8497 11398 8527 11450
rect 8551 11398 8561 11450
rect 8561 11398 8607 11450
rect 8631 11398 8677 11450
rect 8677 11398 8687 11450
rect 8711 11398 8741 11450
rect 8741 11398 8767 11450
rect 8471 11396 8527 11398
rect 8551 11396 8607 11398
rect 8631 11396 8687 11398
rect 8711 11396 8767 11398
rect 8114 11328 8170 11384
rect 8471 10362 8527 10364
rect 8551 10362 8607 10364
rect 8631 10362 8687 10364
rect 8711 10362 8767 10364
rect 8471 10310 8497 10362
rect 8497 10310 8527 10362
rect 8551 10310 8561 10362
rect 8561 10310 8607 10362
rect 8631 10310 8677 10362
rect 8677 10310 8687 10362
rect 8711 10310 8741 10362
rect 8741 10310 8767 10362
rect 8471 10308 8527 10310
rect 8551 10308 8607 10310
rect 8631 10308 8687 10310
rect 8711 10308 8767 10310
rect 9770 14476 9826 14512
rect 9770 14456 9772 14476
rect 9772 14456 9824 14476
rect 9824 14456 9826 14476
rect 12229 21786 12285 21788
rect 12309 21786 12365 21788
rect 12389 21786 12445 21788
rect 12469 21786 12525 21788
rect 12229 21734 12255 21786
rect 12255 21734 12285 21786
rect 12309 21734 12319 21786
rect 12319 21734 12365 21786
rect 12389 21734 12435 21786
rect 12435 21734 12445 21786
rect 12469 21734 12499 21786
rect 12499 21734 12525 21786
rect 12229 21732 12285 21734
rect 12309 21732 12365 21734
rect 12389 21732 12445 21734
rect 12469 21732 12525 21734
rect 12229 20698 12285 20700
rect 12309 20698 12365 20700
rect 12389 20698 12445 20700
rect 12469 20698 12525 20700
rect 12229 20646 12255 20698
rect 12255 20646 12285 20698
rect 12309 20646 12319 20698
rect 12319 20646 12365 20698
rect 12389 20646 12435 20698
rect 12435 20646 12445 20698
rect 12469 20646 12499 20698
rect 12499 20646 12525 20698
rect 12229 20644 12285 20646
rect 12309 20644 12365 20646
rect 12389 20644 12445 20646
rect 12469 20644 12525 20646
rect 11702 17720 11758 17776
rect 8471 9274 8527 9276
rect 8551 9274 8607 9276
rect 8631 9274 8687 9276
rect 8711 9274 8767 9276
rect 8471 9222 8497 9274
rect 8497 9222 8527 9274
rect 8551 9222 8561 9274
rect 8561 9222 8607 9274
rect 8631 9222 8677 9274
rect 8677 9222 8687 9274
rect 8711 9222 8741 9274
rect 8741 9222 8767 9274
rect 8471 9220 8527 9222
rect 8551 9220 8607 9222
rect 8631 9220 8687 9222
rect 8711 9220 8767 9222
rect 8471 8186 8527 8188
rect 8551 8186 8607 8188
rect 8631 8186 8687 8188
rect 8711 8186 8767 8188
rect 8471 8134 8497 8186
rect 8497 8134 8527 8186
rect 8551 8134 8561 8186
rect 8561 8134 8607 8186
rect 8631 8134 8677 8186
rect 8677 8134 8687 8186
rect 8711 8134 8741 8186
rect 8741 8134 8767 8186
rect 8471 8132 8527 8134
rect 8551 8132 8607 8134
rect 8631 8132 8687 8134
rect 8711 8132 8767 8134
rect 8471 7098 8527 7100
rect 8551 7098 8607 7100
rect 8631 7098 8687 7100
rect 8711 7098 8767 7100
rect 8471 7046 8497 7098
rect 8497 7046 8527 7098
rect 8551 7046 8561 7098
rect 8561 7046 8607 7098
rect 8631 7046 8677 7098
rect 8677 7046 8687 7098
rect 8711 7046 8741 7098
rect 8741 7046 8767 7098
rect 8471 7044 8527 7046
rect 8551 7044 8607 7046
rect 8631 7044 8687 7046
rect 8711 7044 8767 7046
rect 8471 6010 8527 6012
rect 8551 6010 8607 6012
rect 8631 6010 8687 6012
rect 8711 6010 8767 6012
rect 8471 5958 8497 6010
rect 8497 5958 8527 6010
rect 8551 5958 8561 6010
rect 8561 5958 8607 6010
rect 8631 5958 8677 6010
rect 8677 5958 8687 6010
rect 8711 5958 8741 6010
rect 8741 5958 8767 6010
rect 8471 5956 8527 5958
rect 8551 5956 8607 5958
rect 8631 5956 8687 5958
rect 8711 5956 8767 5958
rect 8471 4922 8527 4924
rect 8551 4922 8607 4924
rect 8631 4922 8687 4924
rect 8711 4922 8767 4924
rect 8471 4870 8497 4922
rect 8497 4870 8527 4922
rect 8551 4870 8561 4922
rect 8561 4870 8607 4922
rect 8631 4870 8677 4922
rect 8677 4870 8687 4922
rect 8711 4870 8741 4922
rect 8741 4870 8767 4922
rect 8471 4868 8527 4870
rect 8551 4868 8607 4870
rect 8631 4868 8687 4870
rect 8711 4868 8767 4870
rect 7838 3984 7894 4040
rect 6366 40 6422 96
rect 8471 3834 8527 3836
rect 8551 3834 8607 3836
rect 8631 3834 8687 3836
rect 8711 3834 8767 3836
rect 8471 3782 8497 3834
rect 8497 3782 8527 3834
rect 8551 3782 8561 3834
rect 8561 3782 8607 3834
rect 8631 3782 8677 3834
rect 8677 3782 8687 3834
rect 8711 3782 8741 3834
rect 8741 3782 8767 3834
rect 8471 3780 8527 3782
rect 8551 3780 8607 3782
rect 8631 3780 8687 3782
rect 8711 3780 8767 3782
rect 8471 2746 8527 2748
rect 8551 2746 8607 2748
rect 8631 2746 8687 2748
rect 8711 2746 8767 2748
rect 8471 2694 8497 2746
rect 8497 2694 8527 2746
rect 8551 2694 8561 2746
rect 8561 2694 8607 2746
rect 8631 2694 8677 2746
rect 8677 2694 8687 2746
rect 8711 2694 8741 2746
rect 8741 2694 8767 2746
rect 8471 2692 8527 2694
rect 8551 2692 8607 2694
rect 8631 2692 8687 2694
rect 8711 2692 8767 2694
rect 12229 19610 12285 19612
rect 12309 19610 12365 19612
rect 12389 19610 12445 19612
rect 12469 19610 12525 19612
rect 12229 19558 12255 19610
rect 12255 19558 12285 19610
rect 12309 19558 12319 19610
rect 12319 19558 12365 19610
rect 12389 19558 12435 19610
rect 12435 19558 12445 19610
rect 12469 19558 12499 19610
rect 12499 19558 12525 19610
rect 12229 19556 12285 19558
rect 12309 19556 12365 19558
rect 12389 19556 12445 19558
rect 12469 19556 12525 19558
rect 12229 18522 12285 18524
rect 12309 18522 12365 18524
rect 12389 18522 12445 18524
rect 12469 18522 12525 18524
rect 12229 18470 12255 18522
rect 12255 18470 12285 18522
rect 12309 18470 12319 18522
rect 12319 18470 12365 18522
rect 12389 18470 12435 18522
rect 12435 18470 12445 18522
rect 12469 18470 12499 18522
rect 12499 18470 12525 18522
rect 12229 18468 12285 18470
rect 12309 18468 12365 18470
rect 12389 18468 12445 18470
rect 12469 18468 12525 18470
rect 12229 17434 12285 17436
rect 12309 17434 12365 17436
rect 12389 17434 12445 17436
rect 12469 17434 12525 17436
rect 12229 17382 12255 17434
rect 12255 17382 12285 17434
rect 12309 17382 12319 17434
rect 12319 17382 12365 17434
rect 12389 17382 12435 17434
rect 12435 17382 12445 17434
rect 12469 17382 12499 17434
rect 12499 17382 12525 17434
rect 12229 17380 12285 17382
rect 12309 17380 12365 17382
rect 12389 17380 12445 17382
rect 12469 17380 12525 17382
rect 12229 16346 12285 16348
rect 12309 16346 12365 16348
rect 12389 16346 12445 16348
rect 12469 16346 12525 16348
rect 12229 16294 12255 16346
rect 12255 16294 12285 16346
rect 12309 16294 12319 16346
rect 12319 16294 12365 16346
rect 12389 16294 12435 16346
rect 12435 16294 12445 16346
rect 12469 16294 12499 16346
rect 12499 16294 12525 16346
rect 12229 16292 12285 16294
rect 12309 16292 12365 16294
rect 12389 16292 12445 16294
rect 12469 16292 12525 16294
rect 12229 15258 12285 15260
rect 12309 15258 12365 15260
rect 12389 15258 12445 15260
rect 12469 15258 12525 15260
rect 12229 15206 12255 15258
rect 12255 15206 12285 15258
rect 12309 15206 12319 15258
rect 12319 15206 12365 15258
rect 12389 15206 12435 15258
rect 12435 15206 12445 15258
rect 12469 15206 12499 15258
rect 12499 15206 12525 15258
rect 12229 15204 12285 15206
rect 12309 15204 12365 15206
rect 12389 15204 12445 15206
rect 12469 15204 12525 15206
rect 15986 22330 16042 22332
rect 16066 22330 16122 22332
rect 16146 22330 16202 22332
rect 16226 22330 16282 22332
rect 15986 22278 16012 22330
rect 16012 22278 16042 22330
rect 16066 22278 16076 22330
rect 16076 22278 16122 22330
rect 16146 22278 16192 22330
rect 16192 22278 16202 22330
rect 16226 22278 16256 22330
rect 16256 22278 16282 22330
rect 15986 22276 16042 22278
rect 16066 22276 16122 22278
rect 16146 22276 16202 22278
rect 16226 22276 16282 22278
rect 15986 21242 16042 21244
rect 16066 21242 16122 21244
rect 16146 21242 16202 21244
rect 16226 21242 16282 21244
rect 15986 21190 16012 21242
rect 16012 21190 16042 21242
rect 16066 21190 16076 21242
rect 16076 21190 16122 21242
rect 16146 21190 16192 21242
rect 16192 21190 16202 21242
rect 16226 21190 16256 21242
rect 16256 21190 16282 21242
rect 15986 21188 16042 21190
rect 16066 21188 16122 21190
rect 16146 21188 16202 21190
rect 16226 21188 16282 21190
rect 15986 20154 16042 20156
rect 16066 20154 16122 20156
rect 16146 20154 16202 20156
rect 16226 20154 16282 20156
rect 15986 20102 16012 20154
rect 16012 20102 16042 20154
rect 16066 20102 16076 20154
rect 16076 20102 16122 20154
rect 16146 20102 16192 20154
rect 16192 20102 16202 20154
rect 16226 20102 16256 20154
rect 16256 20102 16282 20154
rect 15986 20100 16042 20102
rect 16066 20100 16122 20102
rect 16146 20100 16202 20102
rect 16226 20100 16282 20102
rect 14554 15408 14610 15464
rect 15986 19066 16042 19068
rect 16066 19066 16122 19068
rect 16146 19066 16202 19068
rect 16226 19066 16282 19068
rect 15986 19014 16012 19066
rect 16012 19014 16042 19066
rect 16066 19014 16076 19066
rect 16076 19014 16122 19066
rect 16146 19014 16192 19066
rect 16192 19014 16202 19066
rect 16226 19014 16256 19066
rect 16256 19014 16282 19066
rect 15986 19012 16042 19014
rect 16066 19012 16122 19014
rect 16146 19012 16202 19014
rect 16226 19012 16282 19014
rect 15986 17978 16042 17980
rect 16066 17978 16122 17980
rect 16146 17978 16202 17980
rect 16226 17978 16282 17980
rect 15986 17926 16012 17978
rect 16012 17926 16042 17978
rect 16066 17926 16076 17978
rect 16076 17926 16122 17978
rect 16146 17926 16192 17978
rect 16192 17926 16202 17978
rect 16226 17926 16256 17978
rect 16256 17926 16282 17978
rect 15986 17924 16042 17926
rect 16066 17924 16122 17926
rect 16146 17924 16202 17926
rect 16226 17924 16282 17926
rect 15986 16890 16042 16892
rect 16066 16890 16122 16892
rect 16146 16890 16202 16892
rect 16226 16890 16282 16892
rect 15986 16838 16012 16890
rect 16012 16838 16042 16890
rect 16066 16838 16076 16890
rect 16076 16838 16122 16890
rect 16146 16838 16192 16890
rect 16192 16838 16202 16890
rect 16226 16838 16256 16890
rect 16256 16838 16282 16890
rect 15986 16836 16042 16838
rect 16066 16836 16122 16838
rect 16146 16836 16202 16838
rect 16226 16836 16282 16838
rect 15986 15802 16042 15804
rect 16066 15802 16122 15804
rect 16146 15802 16202 15804
rect 16226 15802 16282 15804
rect 15986 15750 16012 15802
rect 16012 15750 16042 15802
rect 16066 15750 16076 15802
rect 16076 15750 16122 15802
rect 16146 15750 16192 15802
rect 16192 15750 16202 15802
rect 16226 15750 16256 15802
rect 16256 15750 16282 15802
rect 15986 15748 16042 15750
rect 16066 15748 16122 15750
rect 16146 15748 16202 15750
rect 16226 15748 16282 15750
rect 15986 14714 16042 14716
rect 16066 14714 16122 14716
rect 16146 14714 16202 14716
rect 16226 14714 16282 14716
rect 15986 14662 16012 14714
rect 16012 14662 16042 14714
rect 16066 14662 16076 14714
rect 16076 14662 16122 14714
rect 16146 14662 16192 14714
rect 16192 14662 16202 14714
rect 16226 14662 16256 14714
rect 16256 14662 16282 14714
rect 15986 14660 16042 14662
rect 16066 14660 16122 14662
rect 16146 14660 16202 14662
rect 16226 14660 16282 14662
rect 12229 14170 12285 14172
rect 12309 14170 12365 14172
rect 12389 14170 12445 14172
rect 12469 14170 12525 14172
rect 12229 14118 12255 14170
rect 12255 14118 12285 14170
rect 12309 14118 12319 14170
rect 12319 14118 12365 14170
rect 12389 14118 12435 14170
rect 12435 14118 12445 14170
rect 12469 14118 12499 14170
rect 12499 14118 12525 14170
rect 12229 14116 12285 14118
rect 12309 14116 12365 14118
rect 12389 14116 12445 14118
rect 12469 14116 12525 14118
rect 18510 21936 18566 21992
rect 15986 13626 16042 13628
rect 16066 13626 16122 13628
rect 16146 13626 16202 13628
rect 16226 13626 16282 13628
rect 15986 13574 16012 13626
rect 16012 13574 16042 13626
rect 16066 13574 16076 13626
rect 16076 13574 16122 13626
rect 16146 13574 16192 13626
rect 16192 13574 16202 13626
rect 16226 13574 16256 13626
rect 16256 13574 16282 13626
rect 15986 13572 16042 13574
rect 16066 13572 16122 13574
rect 16146 13572 16202 13574
rect 16226 13572 16282 13574
rect 12229 13082 12285 13084
rect 12309 13082 12365 13084
rect 12389 13082 12445 13084
rect 12469 13082 12525 13084
rect 12229 13030 12255 13082
rect 12255 13030 12285 13082
rect 12309 13030 12319 13082
rect 12319 13030 12365 13082
rect 12389 13030 12435 13082
rect 12435 13030 12445 13082
rect 12469 13030 12499 13082
rect 12499 13030 12525 13082
rect 12229 13028 12285 13030
rect 12309 13028 12365 13030
rect 12389 13028 12445 13030
rect 12469 13028 12525 13030
rect 12622 12688 12678 12744
rect 12229 11994 12285 11996
rect 12309 11994 12365 11996
rect 12389 11994 12445 11996
rect 12469 11994 12525 11996
rect 12229 11942 12255 11994
rect 12255 11942 12285 11994
rect 12309 11942 12319 11994
rect 12319 11942 12365 11994
rect 12389 11942 12435 11994
rect 12435 11942 12445 11994
rect 12469 11942 12499 11994
rect 12499 11942 12525 11994
rect 12229 11940 12285 11942
rect 12309 11940 12365 11942
rect 12389 11940 12445 11942
rect 12469 11940 12525 11942
rect 16486 12552 16542 12608
rect 15986 12538 16042 12540
rect 16066 12538 16122 12540
rect 16146 12538 16202 12540
rect 16226 12538 16282 12540
rect 15986 12486 16012 12538
rect 16012 12486 16042 12538
rect 16066 12486 16076 12538
rect 16076 12486 16122 12538
rect 16146 12486 16192 12538
rect 16192 12486 16202 12538
rect 16226 12486 16256 12538
rect 16256 12486 16282 12538
rect 15986 12484 16042 12486
rect 16066 12484 16122 12486
rect 16146 12484 16202 12486
rect 16226 12484 16282 12486
rect 12229 10906 12285 10908
rect 12309 10906 12365 10908
rect 12389 10906 12445 10908
rect 12469 10906 12525 10908
rect 12229 10854 12255 10906
rect 12255 10854 12285 10906
rect 12309 10854 12319 10906
rect 12319 10854 12365 10906
rect 12389 10854 12435 10906
rect 12435 10854 12445 10906
rect 12469 10854 12499 10906
rect 12499 10854 12525 10906
rect 12229 10852 12285 10854
rect 12309 10852 12365 10854
rect 12389 10852 12445 10854
rect 12469 10852 12525 10854
rect 12229 9818 12285 9820
rect 12309 9818 12365 9820
rect 12389 9818 12445 9820
rect 12469 9818 12525 9820
rect 12229 9766 12255 9818
rect 12255 9766 12285 9818
rect 12309 9766 12319 9818
rect 12319 9766 12365 9818
rect 12389 9766 12435 9818
rect 12435 9766 12445 9818
rect 12469 9766 12499 9818
rect 12499 9766 12525 9818
rect 12229 9764 12285 9766
rect 12309 9764 12365 9766
rect 12389 9764 12445 9766
rect 12469 9764 12525 9766
rect 12229 8730 12285 8732
rect 12309 8730 12365 8732
rect 12389 8730 12445 8732
rect 12469 8730 12525 8732
rect 12229 8678 12255 8730
rect 12255 8678 12285 8730
rect 12309 8678 12319 8730
rect 12319 8678 12365 8730
rect 12389 8678 12435 8730
rect 12435 8678 12445 8730
rect 12469 8678 12499 8730
rect 12499 8678 12525 8730
rect 12229 8676 12285 8678
rect 12309 8676 12365 8678
rect 12389 8676 12445 8678
rect 12469 8676 12525 8678
rect 12229 7642 12285 7644
rect 12309 7642 12365 7644
rect 12389 7642 12445 7644
rect 12469 7642 12525 7644
rect 12229 7590 12255 7642
rect 12255 7590 12285 7642
rect 12309 7590 12319 7642
rect 12319 7590 12365 7642
rect 12389 7590 12435 7642
rect 12435 7590 12445 7642
rect 12469 7590 12499 7642
rect 12499 7590 12525 7642
rect 12229 7588 12285 7590
rect 12309 7588 12365 7590
rect 12389 7588 12445 7590
rect 12469 7588 12525 7590
rect 12229 6554 12285 6556
rect 12309 6554 12365 6556
rect 12389 6554 12445 6556
rect 12469 6554 12525 6556
rect 12229 6502 12255 6554
rect 12255 6502 12285 6554
rect 12309 6502 12319 6554
rect 12319 6502 12365 6554
rect 12389 6502 12435 6554
rect 12435 6502 12445 6554
rect 12469 6502 12499 6554
rect 12499 6502 12525 6554
rect 12229 6500 12285 6502
rect 12309 6500 12365 6502
rect 12389 6500 12445 6502
rect 12469 6500 12525 6502
rect 12229 5466 12285 5468
rect 12309 5466 12365 5468
rect 12389 5466 12445 5468
rect 12469 5466 12525 5468
rect 12229 5414 12255 5466
rect 12255 5414 12285 5466
rect 12309 5414 12319 5466
rect 12319 5414 12365 5466
rect 12389 5414 12435 5466
rect 12435 5414 12445 5466
rect 12469 5414 12499 5466
rect 12499 5414 12525 5466
rect 12229 5412 12285 5414
rect 12309 5412 12365 5414
rect 12389 5412 12445 5414
rect 12469 5412 12525 5414
rect 13082 6704 13138 6760
rect 12229 4378 12285 4380
rect 12309 4378 12365 4380
rect 12389 4378 12445 4380
rect 12469 4378 12525 4380
rect 12229 4326 12255 4378
rect 12255 4326 12285 4378
rect 12309 4326 12319 4378
rect 12319 4326 12365 4378
rect 12389 4326 12435 4378
rect 12435 4326 12445 4378
rect 12469 4326 12499 4378
rect 12499 4326 12525 4378
rect 12229 4324 12285 4326
rect 12309 4324 12365 4326
rect 12389 4324 12445 4326
rect 12469 4324 12525 4326
rect 9586 3440 9642 3496
rect 10230 1944 10286 2000
rect 14462 4140 14518 4176
rect 14462 4120 14464 4140
rect 14464 4120 14516 4140
rect 14516 4120 14518 4140
rect 12229 3290 12285 3292
rect 12309 3290 12365 3292
rect 12389 3290 12445 3292
rect 12469 3290 12525 3292
rect 12229 3238 12255 3290
rect 12255 3238 12285 3290
rect 12309 3238 12319 3290
rect 12319 3238 12365 3290
rect 12389 3238 12435 3290
rect 12435 3238 12445 3290
rect 12469 3238 12499 3290
rect 12499 3238 12525 3290
rect 12229 3236 12285 3238
rect 12309 3236 12365 3238
rect 12389 3236 12445 3238
rect 12469 3236 12525 3238
rect 12229 2202 12285 2204
rect 12309 2202 12365 2204
rect 12389 2202 12445 2204
rect 12469 2202 12525 2204
rect 12229 2150 12255 2202
rect 12255 2150 12285 2202
rect 12309 2150 12319 2202
rect 12319 2150 12365 2202
rect 12389 2150 12435 2202
rect 12435 2150 12445 2202
rect 12469 2150 12499 2202
rect 12499 2150 12525 2202
rect 12229 2148 12285 2150
rect 12309 2148 12365 2150
rect 12389 2148 12445 2150
rect 12469 2148 12525 2150
rect 14278 40 14334 96
rect 14922 3440 14978 3496
rect 15986 11450 16042 11452
rect 16066 11450 16122 11452
rect 16146 11450 16202 11452
rect 16226 11450 16282 11452
rect 15986 11398 16012 11450
rect 16012 11398 16042 11450
rect 16066 11398 16076 11450
rect 16076 11398 16122 11450
rect 16146 11398 16192 11450
rect 16192 11398 16202 11450
rect 16226 11398 16256 11450
rect 16256 11398 16282 11450
rect 15986 11396 16042 11398
rect 16066 11396 16122 11398
rect 16146 11396 16202 11398
rect 16226 11396 16282 11398
rect 15986 10362 16042 10364
rect 16066 10362 16122 10364
rect 16146 10362 16202 10364
rect 16226 10362 16282 10364
rect 15986 10310 16012 10362
rect 16012 10310 16042 10362
rect 16066 10310 16076 10362
rect 16076 10310 16122 10362
rect 16146 10310 16192 10362
rect 16192 10310 16202 10362
rect 16226 10310 16256 10362
rect 16256 10310 16282 10362
rect 15986 10308 16042 10310
rect 16066 10308 16122 10310
rect 16146 10308 16202 10310
rect 16226 10308 16282 10310
rect 15986 9274 16042 9276
rect 16066 9274 16122 9276
rect 16146 9274 16202 9276
rect 16226 9274 16282 9276
rect 15986 9222 16012 9274
rect 16012 9222 16042 9274
rect 16066 9222 16076 9274
rect 16076 9222 16122 9274
rect 16146 9222 16192 9274
rect 16192 9222 16202 9274
rect 16226 9222 16256 9274
rect 16256 9222 16282 9274
rect 15986 9220 16042 9222
rect 16066 9220 16122 9222
rect 16146 9220 16202 9222
rect 16226 9220 16282 9222
rect 15986 8186 16042 8188
rect 16066 8186 16122 8188
rect 16146 8186 16202 8188
rect 16226 8186 16282 8188
rect 15986 8134 16012 8186
rect 16012 8134 16042 8186
rect 16066 8134 16076 8186
rect 16076 8134 16122 8186
rect 16146 8134 16192 8186
rect 16192 8134 16202 8186
rect 16226 8134 16256 8186
rect 16256 8134 16282 8186
rect 15986 8132 16042 8134
rect 16066 8132 16122 8134
rect 16146 8132 16202 8134
rect 16226 8132 16282 8134
rect 15986 7098 16042 7100
rect 16066 7098 16122 7100
rect 16146 7098 16202 7100
rect 16226 7098 16282 7100
rect 15986 7046 16012 7098
rect 16012 7046 16042 7098
rect 16066 7046 16076 7098
rect 16076 7046 16122 7098
rect 16146 7046 16192 7098
rect 16192 7046 16202 7098
rect 16226 7046 16256 7098
rect 16256 7046 16282 7098
rect 15986 7044 16042 7046
rect 16066 7044 16122 7046
rect 16146 7044 16202 7046
rect 16226 7044 16282 7046
rect 15986 6010 16042 6012
rect 16066 6010 16122 6012
rect 16146 6010 16202 6012
rect 16226 6010 16282 6012
rect 15986 5958 16012 6010
rect 16012 5958 16042 6010
rect 16066 5958 16076 6010
rect 16076 5958 16122 6010
rect 16146 5958 16192 6010
rect 16192 5958 16202 6010
rect 16226 5958 16256 6010
rect 16256 5958 16282 6010
rect 15986 5956 16042 5958
rect 16066 5956 16122 5958
rect 16146 5956 16202 5958
rect 16226 5956 16282 5958
rect 15986 4922 16042 4924
rect 16066 4922 16122 4924
rect 16146 4922 16202 4924
rect 16226 4922 16282 4924
rect 15986 4870 16012 4922
rect 16012 4870 16042 4922
rect 16066 4870 16076 4922
rect 16076 4870 16122 4922
rect 16146 4870 16192 4922
rect 16192 4870 16202 4922
rect 16226 4870 16256 4922
rect 16256 4870 16282 4922
rect 15986 4868 16042 4870
rect 16066 4868 16122 4870
rect 16146 4868 16202 4870
rect 16226 4868 16282 4870
rect 15986 3834 16042 3836
rect 16066 3834 16122 3836
rect 16146 3834 16202 3836
rect 16226 3834 16282 3836
rect 15986 3782 16012 3834
rect 16012 3782 16042 3834
rect 16066 3782 16076 3834
rect 16076 3782 16122 3834
rect 16146 3782 16192 3834
rect 16192 3782 16202 3834
rect 16226 3782 16256 3834
rect 16256 3782 16282 3834
rect 15986 3780 16042 3782
rect 16066 3780 16122 3782
rect 16146 3780 16202 3782
rect 16226 3780 16282 3782
rect 15986 2746 16042 2748
rect 16066 2746 16122 2748
rect 16146 2746 16202 2748
rect 16226 2746 16282 2748
rect 15986 2694 16012 2746
rect 16012 2694 16042 2746
rect 16066 2694 16076 2746
rect 16076 2694 16122 2746
rect 16146 2694 16192 2746
rect 16192 2694 16202 2746
rect 16226 2694 16256 2746
rect 16256 2694 16282 2746
rect 15986 2692 16042 2694
rect 16066 2692 16122 2694
rect 16146 2692 16202 2694
rect 16226 2692 16282 2694
rect 16486 3576 16542 3632
rect 18418 17720 18474 17776
rect 20166 23296 20222 23352
rect 19744 21786 19800 21788
rect 19824 21786 19880 21788
rect 19904 21786 19960 21788
rect 19984 21786 20040 21788
rect 19744 21734 19770 21786
rect 19770 21734 19800 21786
rect 19824 21734 19834 21786
rect 19834 21734 19880 21786
rect 19904 21734 19950 21786
rect 19950 21734 19960 21786
rect 19984 21734 20014 21786
rect 20014 21734 20040 21786
rect 19744 21732 19800 21734
rect 19824 21732 19880 21734
rect 19904 21732 19960 21734
rect 19984 21732 20040 21734
rect 19744 20698 19800 20700
rect 19824 20698 19880 20700
rect 19904 20698 19960 20700
rect 19984 20698 20040 20700
rect 19744 20646 19770 20698
rect 19770 20646 19800 20698
rect 19824 20646 19834 20698
rect 19834 20646 19880 20698
rect 19904 20646 19950 20698
rect 19950 20646 19960 20698
rect 19984 20646 20014 20698
rect 20014 20646 20040 20698
rect 19744 20644 19800 20646
rect 19824 20644 19880 20646
rect 19904 20644 19960 20646
rect 19984 20644 20040 20646
rect 20350 20168 20406 20224
rect 19744 19610 19800 19612
rect 19824 19610 19880 19612
rect 19904 19610 19960 19612
rect 19984 19610 20040 19612
rect 19744 19558 19770 19610
rect 19770 19558 19800 19610
rect 19824 19558 19834 19610
rect 19834 19558 19880 19610
rect 19904 19558 19950 19610
rect 19950 19558 19960 19610
rect 19984 19558 20014 19610
rect 20014 19558 20040 19610
rect 19744 19556 19800 19558
rect 19824 19556 19880 19558
rect 19904 19556 19960 19558
rect 19984 19556 20040 19558
rect 22098 19216 22154 19272
rect 19744 18522 19800 18524
rect 19824 18522 19880 18524
rect 19904 18522 19960 18524
rect 19984 18522 20040 18524
rect 19744 18470 19770 18522
rect 19770 18470 19800 18522
rect 19824 18470 19834 18522
rect 19834 18470 19880 18522
rect 19904 18470 19950 18522
rect 19950 18470 19960 18522
rect 19984 18470 20014 18522
rect 20014 18470 20040 18522
rect 19744 18468 19800 18470
rect 19824 18468 19880 18470
rect 19904 18468 19960 18470
rect 19984 18468 20040 18470
rect 22098 18128 22154 18184
rect 19744 17434 19800 17436
rect 19824 17434 19880 17436
rect 19904 17434 19960 17436
rect 19984 17434 20040 17436
rect 19744 17382 19770 17434
rect 19770 17382 19800 17434
rect 19824 17382 19834 17434
rect 19834 17382 19880 17434
rect 19904 17382 19950 17434
rect 19950 17382 19960 17434
rect 19984 17382 20014 17434
rect 20014 17382 20040 17434
rect 19744 17380 19800 17382
rect 19824 17380 19880 17382
rect 19904 17380 19960 17382
rect 19984 17380 20040 17382
rect 19798 17176 19854 17232
rect 19522 17040 19578 17096
rect 19744 16346 19800 16348
rect 19824 16346 19880 16348
rect 19904 16346 19960 16348
rect 19984 16346 20040 16348
rect 19744 16294 19770 16346
rect 19770 16294 19800 16346
rect 19824 16294 19834 16346
rect 19834 16294 19880 16346
rect 19904 16294 19950 16346
rect 19950 16294 19960 16346
rect 19984 16294 20014 16346
rect 20014 16294 20040 16346
rect 19744 16292 19800 16294
rect 19824 16292 19880 16294
rect 19904 16292 19960 16294
rect 19984 16292 20040 16294
rect 19062 15544 19118 15600
rect 19744 15258 19800 15260
rect 19824 15258 19880 15260
rect 19904 15258 19960 15260
rect 19984 15258 20040 15260
rect 19744 15206 19770 15258
rect 19770 15206 19800 15258
rect 19824 15206 19834 15258
rect 19834 15206 19880 15258
rect 19904 15206 19950 15258
rect 19950 15206 19960 15258
rect 19984 15206 20014 15258
rect 20014 15206 20040 15258
rect 19744 15204 19800 15206
rect 19824 15204 19880 15206
rect 19904 15204 19960 15206
rect 19984 15204 20040 15206
rect 19744 14170 19800 14172
rect 19824 14170 19880 14172
rect 19904 14170 19960 14172
rect 19984 14170 20040 14172
rect 19744 14118 19770 14170
rect 19770 14118 19800 14170
rect 19824 14118 19834 14170
rect 19834 14118 19880 14170
rect 19904 14118 19950 14170
rect 19950 14118 19960 14170
rect 19984 14118 20014 14170
rect 20014 14118 20040 14170
rect 19744 14116 19800 14118
rect 19824 14116 19880 14118
rect 19904 14116 19960 14118
rect 19984 14116 20040 14118
rect 19744 13082 19800 13084
rect 19824 13082 19880 13084
rect 19904 13082 19960 13084
rect 19984 13082 20040 13084
rect 19744 13030 19770 13082
rect 19770 13030 19800 13082
rect 19824 13030 19834 13082
rect 19834 13030 19880 13082
rect 19904 13030 19950 13082
rect 19950 13030 19960 13082
rect 19984 13030 20014 13082
rect 20014 13030 20040 13082
rect 19744 13028 19800 13030
rect 19824 13028 19880 13030
rect 19904 13028 19960 13030
rect 19984 13028 20040 13030
rect 19744 11994 19800 11996
rect 19824 11994 19880 11996
rect 19904 11994 19960 11996
rect 19984 11994 20040 11996
rect 19744 11942 19770 11994
rect 19770 11942 19800 11994
rect 19824 11942 19834 11994
rect 19834 11942 19880 11994
rect 19904 11942 19950 11994
rect 19950 11942 19960 11994
rect 19984 11942 20014 11994
rect 20014 11942 20040 11994
rect 19744 11940 19800 11942
rect 19824 11940 19880 11942
rect 19904 11940 19960 11942
rect 19984 11940 20040 11942
rect 19798 11464 19854 11520
rect 19744 10906 19800 10908
rect 19824 10906 19880 10908
rect 19904 10906 19960 10908
rect 19984 10906 20040 10908
rect 19744 10854 19770 10906
rect 19770 10854 19800 10906
rect 19824 10854 19834 10906
rect 19834 10854 19880 10906
rect 19904 10854 19950 10906
rect 19950 10854 19960 10906
rect 19984 10854 20014 10906
rect 20014 10854 20040 10906
rect 19744 10852 19800 10854
rect 19824 10852 19880 10854
rect 19904 10852 19960 10854
rect 19984 10852 20040 10854
rect 19744 9818 19800 9820
rect 19824 9818 19880 9820
rect 19904 9818 19960 9820
rect 19984 9818 20040 9820
rect 19744 9766 19770 9818
rect 19770 9766 19800 9818
rect 19824 9766 19834 9818
rect 19834 9766 19880 9818
rect 19904 9766 19950 9818
rect 19950 9766 19960 9818
rect 19984 9766 20014 9818
rect 20014 9766 20040 9818
rect 19744 9764 19800 9766
rect 19824 9764 19880 9766
rect 19904 9764 19960 9766
rect 19984 9764 20040 9766
rect 19744 8730 19800 8732
rect 19824 8730 19880 8732
rect 19904 8730 19960 8732
rect 19984 8730 20040 8732
rect 19744 8678 19770 8730
rect 19770 8678 19800 8730
rect 19824 8678 19834 8730
rect 19834 8678 19880 8730
rect 19904 8678 19950 8730
rect 19950 8678 19960 8730
rect 19984 8678 20014 8730
rect 20014 8678 20040 8730
rect 19744 8676 19800 8678
rect 19824 8676 19880 8678
rect 19904 8676 19960 8678
rect 19984 8676 20040 8678
rect 18694 7792 18750 7848
rect 19744 7642 19800 7644
rect 19824 7642 19880 7644
rect 19904 7642 19960 7644
rect 19984 7642 20040 7644
rect 19744 7590 19770 7642
rect 19770 7590 19800 7642
rect 19824 7590 19834 7642
rect 19834 7590 19880 7642
rect 19904 7590 19950 7642
rect 19950 7590 19960 7642
rect 19984 7590 20014 7642
rect 20014 7590 20040 7642
rect 19744 7588 19800 7590
rect 19824 7588 19880 7590
rect 19904 7588 19960 7590
rect 19984 7588 20040 7590
rect 19744 6554 19800 6556
rect 19824 6554 19880 6556
rect 19904 6554 19960 6556
rect 19984 6554 20040 6556
rect 19744 6502 19770 6554
rect 19770 6502 19800 6554
rect 19824 6502 19834 6554
rect 19834 6502 19880 6554
rect 19904 6502 19950 6554
rect 19950 6502 19960 6554
rect 19984 6502 20014 6554
rect 20014 6502 20040 6554
rect 19744 6500 19800 6502
rect 19824 6500 19880 6502
rect 19904 6500 19960 6502
rect 19984 6500 20040 6502
rect 18786 5616 18842 5672
rect 19744 5466 19800 5468
rect 19824 5466 19880 5468
rect 19904 5466 19960 5468
rect 19984 5466 20040 5468
rect 19744 5414 19770 5466
rect 19770 5414 19800 5466
rect 19824 5414 19834 5466
rect 19834 5414 19880 5466
rect 19904 5414 19950 5466
rect 19950 5414 19960 5466
rect 19984 5414 20014 5466
rect 20014 5414 20040 5466
rect 19744 5412 19800 5414
rect 19824 5412 19880 5414
rect 19904 5412 19960 5414
rect 19984 5412 20040 5414
rect 20166 5344 20222 5400
rect 19744 4378 19800 4380
rect 19824 4378 19880 4380
rect 19904 4378 19960 4380
rect 19984 4378 20040 4380
rect 19744 4326 19770 4378
rect 19770 4326 19800 4378
rect 19824 4326 19834 4378
rect 19834 4326 19880 4378
rect 19904 4326 19950 4378
rect 19950 4326 19960 4378
rect 19984 4326 20014 4378
rect 20014 4326 20040 4378
rect 19744 4324 19800 4326
rect 19824 4324 19880 4326
rect 19904 4324 19960 4326
rect 19984 4324 20040 4326
rect 20074 3984 20130 4040
rect 19744 3290 19800 3292
rect 19824 3290 19880 3292
rect 19904 3290 19960 3292
rect 19984 3290 20040 3292
rect 19744 3238 19770 3290
rect 19770 3238 19800 3290
rect 19824 3238 19834 3290
rect 19834 3238 19880 3290
rect 19904 3238 19950 3290
rect 19950 3238 19960 3290
rect 19984 3238 20014 3290
rect 20014 3238 20040 3290
rect 19744 3236 19800 3238
rect 19824 3236 19880 3238
rect 19904 3236 19960 3238
rect 19984 3236 20040 3238
rect 19744 2202 19800 2204
rect 19824 2202 19880 2204
rect 19904 2202 19960 2204
rect 19984 2202 20040 2204
rect 19744 2150 19770 2202
rect 19770 2150 19800 2202
rect 19824 2150 19834 2202
rect 19834 2150 19880 2202
rect 19904 2150 19950 2202
rect 19950 2150 19960 2202
rect 19984 2150 20014 2202
rect 20014 2150 20040 2202
rect 19744 2148 19800 2150
rect 19824 2148 19880 2150
rect 19904 2148 19960 2150
rect 19984 2148 20040 2150
rect 20166 1264 20222 1320
rect 20626 2760 20682 2816
rect 22098 9968 22154 10024
<< metal3 >>
rect 0 24032 480 24064
rect 0 23976 18 24032
rect 74 23976 480 24032
rect 0 23944 480 23976
rect 22066 23808 22546 23928
rect 20161 23354 20227 23357
rect 22142 23354 22202 23808
rect 20161 23352 22202 23354
rect 20161 23296 20166 23352
rect 20222 23296 22202 23352
rect 20161 23294 22202 23296
rect 20161 23291 20227 23294
rect 0 22672 480 22704
rect 0 22616 110 22672
rect 166 22616 480 22672
rect 0 22584 480 22616
rect 8459 22336 8779 22337
rect 8459 22272 8467 22336
rect 8531 22272 8547 22336
rect 8611 22272 8627 22336
rect 8691 22272 8707 22336
rect 8771 22272 8779 22336
rect 8459 22271 8779 22272
rect 15974 22336 16294 22337
rect 15974 22272 15982 22336
rect 16046 22272 16062 22336
rect 16126 22272 16142 22336
rect 16206 22272 16222 22336
rect 16286 22272 16294 22336
rect 22066 22312 22546 22432
rect 15974 22271 16294 22272
rect 18505 21994 18571 21997
rect 22142 21994 22202 22312
rect 18505 21992 22202 21994
rect 18505 21936 18510 21992
rect 18566 21936 22202 21992
rect 18505 21934 22202 21936
rect 18505 21931 18571 21934
rect 4701 21792 5021 21793
rect 4701 21728 4709 21792
rect 4773 21728 4789 21792
rect 4853 21728 4869 21792
rect 4933 21728 4949 21792
rect 5013 21728 5021 21792
rect 4701 21727 5021 21728
rect 12217 21792 12537 21793
rect 12217 21728 12225 21792
rect 12289 21728 12305 21792
rect 12369 21728 12385 21792
rect 12449 21728 12465 21792
rect 12529 21728 12537 21792
rect 12217 21727 12537 21728
rect 19732 21792 20052 21793
rect 19732 21728 19740 21792
rect 19804 21728 19820 21792
rect 19884 21728 19900 21792
rect 19964 21728 19980 21792
rect 20044 21728 20052 21792
rect 19732 21727 20052 21728
rect 0 21224 480 21344
rect 8459 21248 8779 21249
rect 62 20770 122 21224
rect 8459 21184 8467 21248
rect 8531 21184 8547 21248
rect 8611 21184 8627 21248
rect 8691 21184 8707 21248
rect 8771 21184 8779 21248
rect 8459 21183 8779 21184
rect 15974 21248 16294 21249
rect 15974 21184 15982 21248
rect 16046 21184 16062 21248
rect 16126 21184 16142 21248
rect 16206 21184 16222 21248
rect 16286 21184 16294 21248
rect 15974 21183 16294 21184
rect 1577 20770 1643 20773
rect 62 20768 1643 20770
rect 62 20712 1582 20768
rect 1638 20712 1643 20768
rect 62 20710 1643 20712
rect 1577 20707 1643 20710
rect 4701 20704 5021 20705
rect 4701 20640 4709 20704
rect 4773 20640 4789 20704
rect 4853 20640 4869 20704
rect 4933 20640 4949 20704
rect 5013 20640 5021 20704
rect 4701 20639 5021 20640
rect 12217 20704 12537 20705
rect 12217 20640 12225 20704
rect 12289 20640 12305 20704
rect 12369 20640 12385 20704
rect 12449 20640 12465 20704
rect 12529 20640 12537 20704
rect 12217 20639 12537 20640
rect 19732 20704 20052 20705
rect 19732 20640 19740 20704
rect 19804 20640 19820 20704
rect 19884 20640 19900 20704
rect 19964 20640 19980 20704
rect 20044 20640 20052 20704
rect 22066 20680 22546 20800
rect 19732 20639 20052 20640
rect 20345 20226 20411 20229
rect 22142 20226 22202 20680
rect 20345 20224 22202 20226
rect 20345 20168 20350 20224
rect 20406 20168 22202 20224
rect 20345 20166 22202 20168
rect 20345 20163 20411 20166
rect 8459 20160 8779 20161
rect 8459 20096 8467 20160
rect 8531 20096 8547 20160
rect 8611 20096 8627 20160
rect 8691 20096 8707 20160
rect 8771 20096 8779 20160
rect 8459 20095 8779 20096
rect 15974 20160 16294 20161
rect 15974 20096 15982 20160
rect 16046 20096 16062 20160
rect 16126 20096 16142 20160
rect 16206 20096 16222 20160
rect 16286 20096 16294 20160
rect 15974 20095 16294 20096
rect 0 19864 480 19984
rect 62 19410 122 19864
rect 4701 19616 5021 19617
rect 4701 19552 4709 19616
rect 4773 19552 4789 19616
rect 4853 19552 4869 19616
rect 4933 19552 4949 19616
rect 5013 19552 5021 19616
rect 4701 19551 5021 19552
rect 12217 19616 12537 19617
rect 12217 19552 12225 19616
rect 12289 19552 12305 19616
rect 12369 19552 12385 19616
rect 12449 19552 12465 19616
rect 12529 19552 12537 19616
rect 12217 19551 12537 19552
rect 19732 19616 20052 19617
rect 19732 19552 19740 19616
rect 19804 19552 19820 19616
rect 19884 19552 19900 19616
rect 19964 19552 19980 19616
rect 20044 19552 20052 19616
rect 19732 19551 20052 19552
rect 1577 19410 1643 19413
rect 62 19408 1643 19410
rect 62 19352 1582 19408
rect 1638 19352 1643 19408
rect 62 19350 1643 19352
rect 1577 19347 1643 19350
rect 22066 19274 22546 19304
rect 22012 19272 22546 19274
rect 22012 19216 22098 19272
rect 22154 19216 22546 19272
rect 22012 19214 22546 19216
rect 22066 19184 22546 19214
rect 8459 19072 8779 19073
rect 8459 19008 8467 19072
rect 8531 19008 8547 19072
rect 8611 19008 8627 19072
rect 8691 19008 8707 19072
rect 8771 19008 8779 19072
rect 8459 19007 8779 19008
rect 15974 19072 16294 19073
rect 15974 19008 15982 19072
rect 16046 19008 16062 19072
rect 16126 19008 16142 19072
rect 16206 19008 16222 19072
rect 16286 19008 16294 19072
rect 15974 19007 16294 19008
rect 0 18504 480 18624
rect 4701 18528 5021 18529
rect 62 18050 122 18504
rect 4701 18464 4709 18528
rect 4773 18464 4789 18528
rect 4853 18464 4869 18528
rect 4933 18464 4949 18528
rect 5013 18464 5021 18528
rect 4701 18463 5021 18464
rect 12217 18528 12537 18529
rect 12217 18464 12225 18528
rect 12289 18464 12305 18528
rect 12369 18464 12385 18528
rect 12449 18464 12465 18528
rect 12529 18464 12537 18528
rect 12217 18463 12537 18464
rect 19732 18528 20052 18529
rect 19732 18464 19740 18528
rect 19804 18464 19820 18528
rect 19884 18464 19900 18528
rect 19964 18464 19980 18528
rect 20044 18464 20052 18528
rect 19732 18463 20052 18464
rect 8845 18186 8911 18189
rect 22093 18186 22159 18189
rect 8845 18184 22159 18186
rect 8845 18128 8850 18184
rect 8906 18128 22098 18184
rect 22154 18128 22159 18184
rect 8845 18126 22159 18128
rect 8845 18123 8911 18126
rect 22093 18123 22159 18126
rect 6269 18050 6335 18053
rect 62 18048 6335 18050
rect 62 17992 6274 18048
rect 6330 17992 6335 18048
rect 62 17990 6335 17992
rect 6269 17987 6335 17990
rect 8459 17984 8779 17985
rect 8459 17920 8467 17984
rect 8531 17920 8547 17984
rect 8611 17920 8627 17984
rect 8691 17920 8707 17984
rect 8771 17920 8779 17984
rect 8459 17919 8779 17920
rect 15974 17984 16294 17985
rect 15974 17920 15982 17984
rect 16046 17920 16062 17984
rect 16126 17920 16142 17984
rect 16206 17920 16222 17984
rect 16286 17920 16294 17984
rect 15974 17919 16294 17920
rect 11697 17778 11763 17781
rect 18413 17778 18479 17781
rect 11697 17776 18479 17778
rect 11697 17720 11702 17776
rect 11758 17720 18418 17776
rect 18474 17720 18479 17776
rect 11697 17718 18479 17720
rect 11697 17715 11763 17718
rect 18413 17715 18479 17718
rect 22066 17688 22546 17808
rect 4701 17440 5021 17441
rect 4701 17376 4709 17440
rect 4773 17376 4789 17440
rect 4853 17376 4869 17440
rect 4933 17376 4949 17440
rect 5013 17376 5021 17440
rect 4701 17375 5021 17376
rect 12217 17440 12537 17441
rect 12217 17376 12225 17440
rect 12289 17376 12305 17440
rect 12369 17376 12385 17440
rect 12449 17376 12465 17440
rect 12529 17376 12537 17440
rect 12217 17375 12537 17376
rect 19732 17440 20052 17441
rect 19732 17376 19740 17440
rect 19804 17376 19820 17440
rect 19884 17376 19900 17440
rect 19964 17376 19980 17440
rect 20044 17376 20052 17440
rect 19732 17375 20052 17376
rect 0 17144 480 17264
rect 19793 17234 19859 17237
rect 22142 17234 22202 17688
rect 19793 17232 22202 17234
rect 19793 17176 19798 17232
rect 19854 17176 22202 17232
rect 19793 17174 22202 17176
rect 19793 17171 19859 17174
rect 62 16690 122 17144
rect 7741 17098 7807 17101
rect 19517 17098 19583 17101
rect 7741 17096 19583 17098
rect 7741 17040 7746 17096
rect 7802 17040 19522 17096
rect 19578 17040 19583 17096
rect 7741 17038 19583 17040
rect 7741 17035 7807 17038
rect 19517 17035 19583 17038
rect 8459 16896 8779 16897
rect 8459 16832 8467 16896
rect 8531 16832 8547 16896
rect 8611 16832 8627 16896
rect 8691 16832 8707 16896
rect 8771 16832 8779 16896
rect 8459 16831 8779 16832
rect 15974 16896 16294 16897
rect 15974 16832 15982 16896
rect 16046 16832 16062 16896
rect 16126 16832 16142 16896
rect 16206 16832 16222 16896
rect 16286 16832 16294 16896
rect 15974 16831 16294 16832
rect 5349 16690 5415 16693
rect 62 16688 5415 16690
rect 62 16632 5354 16688
rect 5410 16632 5415 16688
rect 62 16630 5415 16632
rect 5349 16627 5415 16630
rect 4701 16352 5021 16353
rect 4701 16288 4709 16352
rect 4773 16288 4789 16352
rect 4853 16288 4869 16352
rect 4933 16288 4949 16352
rect 5013 16288 5021 16352
rect 4701 16287 5021 16288
rect 12217 16352 12537 16353
rect 12217 16288 12225 16352
rect 12289 16288 12305 16352
rect 12369 16288 12385 16352
rect 12449 16288 12465 16352
rect 12529 16288 12537 16352
rect 12217 16287 12537 16288
rect 19732 16352 20052 16353
rect 19732 16288 19740 16352
rect 19804 16288 19820 16352
rect 19884 16288 19900 16352
rect 19964 16288 19980 16352
rect 20044 16288 20052 16352
rect 19732 16287 20052 16288
rect 22066 16056 22546 16176
rect 0 15784 480 15904
rect 8459 15808 8779 15809
rect 62 15466 122 15784
rect 8459 15744 8467 15808
rect 8531 15744 8547 15808
rect 8611 15744 8627 15808
rect 8691 15744 8707 15808
rect 8771 15744 8779 15808
rect 8459 15743 8779 15744
rect 15974 15808 16294 15809
rect 15974 15744 15982 15808
rect 16046 15744 16062 15808
rect 16126 15744 16142 15808
rect 16206 15744 16222 15808
rect 16286 15744 16294 15808
rect 15974 15743 16294 15744
rect 19057 15602 19123 15605
rect 22142 15602 22202 16056
rect 19057 15600 22202 15602
rect 19057 15544 19062 15600
rect 19118 15544 22202 15600
rect 19057 15542 22202 15544
rect 19057 15539 19123 15542
rect 14549 15466 14615 15469
rect 62 15464 14615 15466
rect 62 15408 14554 15464
rect 14610 15408 14615 15464
rect 62 15406 14615 15408
rect 14549 15403 14615 15406
rect 4701 15264 5021 15265
rect 4701 15200 4709 15264
rect 4773 15200 4789 15264
rect 4853 15200 4869 15264
rect 4933 15200 4949 15264
rect 5013 15200 5021 15264
rect 4701 15199 5021 15200
rect 12217 15264 12537 15265
rect 12217 15200 12225 15264
rect 12289 15200 12305 15264
rect 12369 15200 12385 15264
rect 12449 15200 12465 15264
rect 12529 15200 12537 15264
rect 12217 15199 12537 15200
rect 19732 15264 20052 15265
rect 19732 15200 19740 15264
rect 19804 15200 19820 15264
rect 19884 15200 19900 15264
rect 19964 15200 19980 15264
rect 20044 15200 20052 15264
rect 19732 15199 20052 15200
rect 54 14860 60 14924
rect 124 14922 130 14924
rect 9489 14922 9555 14925
rect 124 14920 9555 14922
rect 124 14864 9494 14920
rect 9550 14864 9555 14920
rect 124 14862 9555 14864
rect 124 14860 130 14862
rect 9489 14859 9555 14862
rect 8459 14720 8779 14721
rect 8459 14656 8467 14720
rect 8531 14656 8547 14720
rect 8611 14656 8627 14720
rect 8691 14656 8707 14720
rect 8771 14656 8779 14720
rect 8459 14655 8779 14656
rect 15974 14720 16294 14721
rect 15974 14656 15982 14720
rect 16046 14656 16062 14720
rect 16126 14656 16142 14720
rect 16206 14656 16222 14720
rect 16286 14656 16294 14720
rect 15974 14655 16294 14656
rect 22066 14652 22546 14680
rect 22066 14650 22140 14652
rect 22012 14590 22140 14650
rect 22066 14588 22140 14590
rect 22204 14588 22546 14652
rect 22066 14560 22546 14588
rect 0 14516 480 14544
rect 0 14452 60 14516
rect 124 14452 480 14516
rect 0 14424 480 14452
rect 9765 14514 9831 14517
rect 9765 14512 19350 14514
rect 9765 14456 9770 14512
rect 9826 14456 19350 14512
rect 9765 14454 19350 14456
rect 9765 14451 9831 14454
rect 19290 14378 19350 14454
rect 22134 14378 22140 14380
rect 19290 14318 22140 14378
rect 22134 14316 22140 14318
rect 22204 14316 22210 14380
rect 4701 14176 5021 14177
rect 4701 14112 4709 14176
rect 4773 14112 4789 14176
rect 4853 14112 4869 14176
rect 4933 14112 4949 14176
rect 5013 14112 5021 14176
rect 4701 14111 5021 14112
rect 12217 14176 12537 14177
rect 12217 14112 12225 14176
rect 12289 14112 12305 14176
rect 12369 14112 12385 14176
rect 12449 14112 12465 14176
rect 12529 14112 12537 14176
rect 12217 14111 12537 14112
rect 19732 14176 20052 14177
rect 19732 14112 19740 14176
rect 19804 14112 19820 14176
rect 19884 14112 19900 14176
rect 19964 14112 19980 14176
rect 20044 14112 20052 14176
rect 19732 14111 20052 14112
rect 8459 13632 8779 13633
rect 8459 13568 8467 13632
rect 8531 13568 8547 13632
rect 8611 13568 8627 13632
rect 8691 13568 8707 13632
rect 8771 13568 8779 13632
rect 8459 13567 8779 13568
rect 15974 13632 16294 13633
rect 15974 13568 15982 13632
rect 16046 13568 16062 13632
rect 16126 13568 16142 13632
rect 16206 13568 16222 13632
rect 16286 13568 16294 13632
rect 15974 13567 16294 13568
rect 0 13064 480 13184
rect 4701 13088 5021 13089
rect 62 12746 122 13064
rect 4701 13024 4709 13088
rect 4773 13024 4789 13088
rect 4853 13024 4869 13088
rect 4933 13024 4949 13088
rect 5013 13024 5021 13088
rect 4701 13023 5021 13024
rect 12217 13088 12537 13089
rect 12217 13024 12225 13088
rect 12289 13024 12305 13088
rect 12369 13024 12385 13088
rect 12449 13024 12465 13088
rect 12529 13024 12537 13088
rect 12217 13023 12537 13024
rect 19732 13088 20052 13089
rect 19732 13024 19740 13088
rect 19804 13024 19820 13088
rect 19884 13024 19900 13088
rect 19964 13024 19980 13088
rect 20044 13024 20052 13088
rect 22066 13064 22546 13184
rect 19732 13023 20052 13024
rect 12617 12746 12683 12749
rect 62 12744 12683 12746
rect 62 12688 12622 12744
rect 12678 12688 12683 12744
rect 62 12686 12683 12688
rect 12617 12683 12683 12686
rect 16481 12610 16547 12613
rect 22142 12610 22202 13064
rect 16481 12608 22202 12610
rect 16481 12552 16486 12608
rect 16542 12552 22202 12608
rect 16481 12550 22202 12552
rect 16481 12547 16547 12550
rect 8459 12544 8779 12545
rect 8459 12480 8467 12544
rect 8531 12480 8547 12544
rect 8611 12480 8627 12544
rect 8691 12480 8707 12544
rect 8771 12480 8779 12544
rect 8459 12479 8779 12480
rect 15974 12544 16294 12545
rect 15974 12480 15982 12544
rect 16046 12480 16062 12544
rect 16126 12480 16142 12544
rect 16206 12480 16222 12544
rect 16286 12480 16294 12544
rect 15974 12479 16294 12480
rect 4701 12000 5021 12001
rect 4701 11936 4709 12000
rect 4773 11936 4789 12000
rect 4853 11936 4869 12000
rect 4933 11936 4949 12000
rect 5013 11936 5021 12000
rect 4701 11935 5021 11936
rect 12217 12000 12537 12001
rect 12217 11936 12225 12000
rect 12289 11936 12305 12000
rect 12369 11936 12385 12000
rect 12449 11936 12465 12000
rect 12529 11936 12537 12000
rect 12217 11935 12537 11936
rect 19732 12000 20052 12001
rect 19732 11936 19740 12000
rect 19804 11936 19820 12000
rect 19884 11936 19900 12000
rect 19964 11936 19980 12000
rect 20044 11936 20052 12000
rect 19732 11935 20052 11936
rect 0 11568 480 11688
rect 62 11386 122 11568
rect 19793 11522 19859 11525
rect 22066 11522 22546 11552
rect 19793 11520 22546 11522
rect 19793 11464 19798 11520
rect 19854 11464 22546 11520
rect 19793 11462 22546 11464
rect 19793 11459 19859 11462
rect 8459 11456 8779 11457
rect 8459 11392 8467 11456
rect 8531 11392 8547 11456
rect 8611 11392 8627 11456
rect 8691 11392 8707 11456
rect 8771 11392 8779 11456
rect 8459 11391 8779 11392
rect 15974 11456 16294 11457
rect 15974 11392 15982 11456
rect 16046 11392 16062 11456
rect 16126 11392 16142 11456
rect 16206 11392 16222 11456
rect 16286 11392 16294 11456
rect 22066 11432 22546 11462
rect 15974 11391 16294 11392
rect 8109 11386 8175 11389
rect 62 11384 8175 11386
rect 62 11328 8114 11384
rect 8170 11328 8175 11384
rect 62 11326 8175 11328
rect 8109 11323 8175 11326
rect 4701 10912 5021 10913
rect 4701 10848 4709 10912
rect 4773 10848 4789 10912
rect 4853 10848 4869 10912
rect 4933 10848 4949 10912
rect 5013 10848 5021 10912
rect 4701 10847 5021 10848
rect 12217 10912 12537 10913
rect 12217 10848 12225 10912
rect 12289 10848 12305 10912
rect 12369 10848 12385 10912
rect 12449 10848 12465 10912
rect 12529 10848 12537 10912
rect 12217 10847 12537 10848
rect 19732 10912 20052 10913
rect 19732 10848 19740 10912
rect 19804 10848 19820 10912
rect 19884 10848 19900 10912
rect 19964 10848 19980 10912
rect 20044 10848 20052 10912
rect 19732 10847 20052 10848
rect 8459 10368 8779 10369
rect 0 10296 480 10328
rect 8459 10304 8467 10368
rect 8531 10304 8547 10368
rect 8611 10304 8627 10368
rect 8691 10304 8707 10368
rect 8771 10304 8779 10368
rect 8459 10303 8779 10304
rect 15974 10368 16294 10369
rect 15974 10304 15982 10368
rect 16046 10304 16062 10368
rect 16126 10304 16142 10368
rect 16206 10304 16222 10368
rect 16286 10304 16294 10368
rect 15974 10303 16294 10304
rect 0 10240 110 10296
rect 166 10240 480 10296
rect 0 10208 480 10240
rect 22066 10026 22546 10056
rect 22012 10024 22546 10026
rect 22012 9968 22098 10024
rect 22154 9968 22546 10024
rect 22012 9966 22546 9968
rect 22066 9936 22546 9966
rect 4701 9824 5021 9825
rect 4701 9760 4709 9824
rect 4773 9760 4789 9824
rect 4853 9760 4869 9824
rect 4933 9760 4949 9824
rect 5013 9760 5021 9824
rect 4701 9759 5021 9760
rect 12217 9824 12537 9825
rect 12217 9760 12225 9824
rect 12289 9760 12305 9824
rect 12369 9760 12385 9824
rect 12449 9760 12465 9824
rect 12529 9760 12537 9824
rect 12217 9759 12537 9760
rect 19732 9824 20052 9825
rect 19732 9760 19740 9824
rect 19804 9760 19820 9824
rect 19884 9760 19900 9824
rect 19964 9760 19980 9824
rect 20044 9760 20052 9824
rect 19732 9759 20052 9760
rect 8459 9280 8779 9281
rect 8459 9216 8467 9280
rect 8531 9216 8547 9280
rect 8611 9216 8627 9280
rect 8691 9216 8707 9280
rect 8771 9216 8779 9280
rect 8459 9215 8779 9216
rect 15974 9280 16294 9281
rect 15974 9216 15982 9280
rect 16046 9216 16062 9280
rect 16126 9216 16142 9280
rect 16206 9216 16222 9280
rect 16286 9216 16294 9280
rect 15974 9215 16294 9216
rect 0 8848 480 8968
rect 62 8394 122 8848
rect 4701 8736 5021 8737
rect 4701 8672 4709 8736
rect 4773 8672 4789 8736
rect 4853 8672 4869 8736
rect 4933 8672 4949 8736
rect 5013 8672 5021 8736
rect 4701 8671 5021 8672
rect 12217 8736 12537 8737
rect 12217 8672 12225 8736
rect 12289 8672 12305 8736
rect 12369 8672 12385 8736
rect 12449 8672 12465 8736
rect 12529 8672 12537 8736
rect 12217 8671 12537 8672
rect 19732 8736 20052 8737
rect 19732 8672 19740 8736
rect 19804 8672 19820 8736
rect 19884 8672 19900 8736
rect 19964 8672 19980 8736
rect 20044 8672 20052 8736
rect 19732 8671 20052 8672
rect 1853 8394 1919 8397
rect 62 8392 1919 8394
rect 62 8336 1858 8392
rect 1914 8336 1919 8392
rect 62 8334 1919 8336
rect 1853 8331 1919 8334
rect 22066 8304 22546 8424
rect 8459 8192 8779 8193
rect 8459 8128 8467 8192
rect 8531 8128 8547 8192
rect 8611 8128 8627 8192
rect 8691 8128 8707 8192
rect 8771 8128 8779 8192
rect 8459 8127 8779 8128
rect 15974 8192 16294 8193
rect 15974 8128 15982 8192
rect 16046 8128 16062 8192
rect 16126 8128 16142 8192
rect 16206 8128 16222 8192
rect 16286 8128 16294 8192
rect 15974 8127 16294 8128
rect 18689 7850 18755 7853
rect 22142 7850 22202 8304
rect 18689 7848 22202 7850
rect 18689 7792 18694 7848
rect 18750 7792 22202 7848
rect 18689 7790 22202 7792
rect 18689 7787 18755 7790
rect 4701 7648 5021 7649
rect 0 7488 480 7608
rect 4701 7584 4709 7648
rect 4773 7584 4789 7648
rect 4853 7584 4869 7648
rect 4933 7584 4949 7648
rect 5013 7584 5021 7648
rect 4701 7583 5021 7584
rect 12217 7648 12537 7649
rect 12217 7584 12225 7648
rect 12289 7584 12305 7648
rect 12369 7584 12385 7648
rect 12449 7584 12465 7648
rect 12529 7584 12537 7648
rect 12217 7583 12537 7584
rect 19732 7648 20052 7649
rect 19732 7584 19740 7648
rect 19804 7584 19820 7648
rect 19884 7584 19900 7648
rect 19964 7584 19980 7648
rect 20044 7584 20052 7648
rect 19732 7583 20052 7584
rect 62 7034 122 7488
rect 8459 7104 8779 7105
rect 8459 7040 8467 7104
rect 8531 7040 8547 7104
rect 8611 7040 8627 7104
rect 8691 7040 8707 7104
rect 8771 7040 8779 7104
rect 8459 7039 8779 7040
rect 15974 7104 16294 7105
rect 15974 7040 15982 7104
rect 16046 7040 16062 7104
rect 16126 7040 16142 7104
rect 16206 7040 16222 7104
rect 16286 7040 16294 7104
rect 15974 7039 16294 7040
rect 2497 7034 2563 7037
rect 62 7032 2563 7034
rect 62 6976 2502 7032
rect 2558 6976 2563 7032
rect 62 6974 2563 6976
rect 2497 6971 2563 6974
rect 22066 6900 22546 6928
rect 22066 6898 22140 6900
rect 22012 6838 22140 6898
rect 22066 6836 22140 6838
rect 22204 6836 22546 6900
rect 22066 6808 22546 6836
rect 13077 6762 13143 6765
rect 13077 6760 22018 6762
rect 13077 6704 13082 6760
rect 13138 6728 22018 6760
rect 22134 6728 22140 6730
rect 13138 6704 22140 6728
rect 13077 6702 22140 6704
rect 13077 6699 13143 6702
rect 21958 6668 22140 6702
rect 22134 6666 22140 6668
rect 22204 6666 22210 6730
rect 4701 6560 5021 6561
rect 4701 6496 4709 6560
rect 4773 6496 4789 6560
rect 4853 6496 4869 6560
rect 4933 6496 4949 6560
rect 5013 6496 5021 6560
rect 4701 6495 5021 6496
rect 12217 6560 12537 6561
rect 12217 6496 12225 6560
rect 12289 6496 12305 6560
rect 12369 6496 12385 6560
rect 12449 6496 12465 6560
rect 12529 6496 12537 6560
rect 12217 6495 12537 6496
rect 19732 6560 20052 6561
rect 19732 6496 19740 6560
rect 19804 6496 19820 6560
rect 19884 6496 19900 6560
rect 19964 6496 19980 6560
rect 20044 6496 20052 6560
rect 19732 6495 20052 6496
rect 0 6128 480 6248
rect 62 5674 122 6128
rect 8459 6016 8779 6017
rect 8459 5952 8467 6016
rect 8531 5952 8547 6016
rect 8611 5952 8627 6016
rect 8691 5952 8707 6016
rect 8771 5952 8779 6016
rect 8459 5951 8779 5952
rect 15974 6016 16294 6017
rect 15974 5952 15982 6016
rect 16046 5952 16062 6016
rect 16126 5952 16142 6016
rect 16206 5952 16222 6016
rect 16286 5952 16294 6016
rect 15974 5951 16294 5952
rect 1209 5674 1275 5677
rect 62 5672 1275 5674
rect 62 5616 1214 5672
rect 1270 5616 1275 5672
rect 62 5614 1275 5616
rect 1209 5611 1275 5614
rect 3417 5674 3483 5677
rect 18781 5674 18847 5677
rect 3417 5672 18847 5674
rect 3417 5616 3422 5672
rect 3478 5616 18786 5672
rect 18842 5616 18847 5672
rect 3417 5614 18847 5616
rect 3417 5611 3483 5614
rect 18781 5611 18847 5614
rect 4701 5472 5021 5473
rect 4701 5408 4709 5472
rect 4773 5408 4789 5472
rect 4853 5408 4869 5472
rect 4933 5408 4949 5472
rect 5013 5408 5021 5472
rect 4701 5407 5021 5408
rect 12217 5472 12537 5473
rect 12217 5408 12225 5472
rect 12289 5408 12305 5472
rect 12369 5408 12385 5472
rect 12449 5408 12465 5472
rect 12529 5408 12537 5472
rect 12217 5407 12537 5408
rect 19732 5472 20052 5473
rect 19732 5408 19740 5472
rect 19804 5408 19820 5472
rect 19884 5408 19900 5472
rect 19964 5408 19980 5472
rect 20044 5408 20052 5472
rect 19732 5407 20052 5408
rect 20161 5402 20227 5405
rect 22066 5402 22546 5432
rect 20161 5400 22546 5402
rect 20161 5344 20166 5400
rect 20222 5344 22546 5400
rect 20161 5342 22546 5344
rect 20161 5339 20227 5342
rect 22066 5312 22546 5342
rect 8459 4928 8779 4929
rect 0 4768 480 4888
rect 8459 4864 8467 4928
rect 8531 4864 8547 4928
rect 8611 4864 8627 4928
rect 8691 4864 8707 4928
rect 8771 4864 8779 4928
rect 8459 4863 8779 4864
rect 15974 4928 16294 4929
rect 15974 4864 15982 4928
rect 16046 4864 16062 4928
rect 16126 4864 16142 4928
rect 16206 4864 16222 4928
rect 16286 4864 16294 4928
rect 15974 4863 16294 4864
rect 62 4450 122 4768
rect 1853 4450 1919 4453
rect 62 4448 1919 4450
rect 62 4392 1858 4448
rect 1914 4392 1919 4448
rect 62 4390 1919 4392
rect 1853 4387 1919 4390
rect 4701 4384 5021 4385
rect 4701 4320 4709 4384
rect 4773 4320 4789 4384
rect 4853 4320 4869 4384
rect 4933 4320 4949 4384
rect 5013 4320 5021 4384
rect 4701 4319 5021 4320
rect 12217 4384 12537 4385
rect 12217 4320 12225 4384
rect 12289 4320 12305 4384
rect 12369 4320 12385 4384
rect 12449 4320 12465 4384
rect 12529 4320 12537 4384
rect 12217 4319 12537 4320
rect 19732 4384 20052 4385
rect 19732 4320 19740 4384
rect 19804 4320 19820 4384
rect 19884 4320 19900 4384
rect 19964 4320 19980 4384
rect 20044 4320 20052 4384
rect 19732 4319 20052 4320
rect 5073 4178 5139 4181
rect 6269 4178 6335 4181
rect 14457 4178 14523 4181
rect 5073 4176 14523 4178
rect 5073 4120 5078 4176
rect 5134 4120 6274 4176
rect 6330 4120 14462 4176
rect 14518 4120 14523 4176
rect 5073 4118 14523 4120
rect 5073 4115 5139 4118
rect 6269 4115 6335 4118
rect 14457 4115 14523 4118
rect 7833 4042 7899 4045
rect 20069 4042 20135 4045
rect 7833 4040 20135 4042
rect 7833 3984 7838 4040
rect 7894 3984 20074 4040
rect 20130 3984 20135 4040
rect 7833 3982 20135 3984
rect 7833 3979 7899 3982
rect 20069 3979 20135 3982
rect 8459 3840 8779 3841
rect 8459 3776 8467 3840
rect 8531 3776 8547 3840
rect 8611 3776 8627 3840
rect 8691 3776 8707 3840
rect 8771 3776 8779 3840
rect 8459 3775 8779 3776
rect 15974 3840 16294 3841
rect 15974 3776 15982 3840
rect 16046 3776 16062 3840
rect 16126 3776 16142 3840
rect 16206 3776 16222 3840
rect 16286 3776 16294 3840
rect 15974 3775 16294 3776
rect 22066 3680 22546 3800
rect 16481 3634 16547 3637
rect 13770 3632 16547 3634
rect 13770 3576 16486 3632
rect 16542 3576 16547 3632
rect 13770 3574 16547 3576
rect 0 3408 480 3528
rect 9581 3498 9647 3501
rect 13770 3498 13830 3574
rect 16481 3571 16547 3574
rect 9581 3496 13830 3498
rect 9581 3440 9586 3496
rect 9642 3440 13830 3496
rect 9581 3438 13830 3440
rect 14917 3498 14983 3501
rect 22142 3498 22202 3680
rect 14917 3496 22202 3498
rect 14917 3440 14922 3496
rect 14978 3440 22202 3496
rect 14917 3438 22202 3440
rect 9581 3435 9647 3438
rect 14917 3435 14983 3438
rect 4701 3296 5021 3297
rect 4701 3232 4709 3296
rect 4773 3232 4789 3296
rect 4853 3232 4869 3296
rect 4933 3232 4949 3296
rect 5013 3232 5021 3296
rect 4701 3231 5021 3232
rect 12217 3296 12537 3297
rect 12217 3232 12225 3296
rect 12289 3232 12305 3296
rect 12369 3232 12385 3296
rect 12449 3232 12465 3296
rect 12529 3232 12537 3296
rect 12217 3231 12537 3232
rect 19732 3296 20052 3297
rect 19732 3232 19740 3296
rect 19804 3232 19820 3296
rect 19884 3232 19900 3296
rect 19964 3232 19980 3296
rect 20044 3232 20052 3296
rect 19732 3231 20052 3232
rect 20621 2818 20687 2821
rect 20621 2816 22202 2818
rect 20621 2760 20626 2816
rect 20682 2760 22202 2816
rect 20621 2758 22202 2760
rect 20621 2755 20687 2758
rect 8459 2752 8779 2753
rect 8459 2688 8467 2752
rect 8531 2688 8547 2752
rect 8611 2688 8627 2752
rect 8691 2688 8707 2752
rect 8771 2688 8779 2752
rect 8459 2687 8779 2688
rect 15974 2752 16294 2753
rect 15974 2688 15982 2752
rect 16046 2688 16062 2752
rect 16126 2688 16142 2752
rect 16206 2688 16222 2752
rect 16286 2688 16294 2752
rect 15974 2687 16294 2688
rect 22142 2304 22202 2758
rect 4701 2208 5021 2209
rect 0 2048 480 2168
rect 4701 2144 4709 2208
rect 4773 2144 4789 2208
rect 4853 2144 4869 2208
rect 4933 2144 4949 2208
rect 5013 2144 5021 2208
rect 4701 2143 5021 2144
rect 12217 2208 12537 2209
rect 12217 2144 12225 2208
rect 12289 2144 12305 2208
rect 12369 2144 12385 2208
rect 12449 2144 12465 2208
rect 12529 2144 12537 2208
rect 12217 2143 12537 2144
rect 19732 2208 20052 2209
rect 19732 2144 19740 2208
rect 19804 2144 19820 2208
rect 19884 2144 19900 2208
rect 19964 2144 19980 2208
rect 20044 2144 20052 2208
rect 22066 2184 22546 2304
rect 19732 2143 20052 2144
rect 2497 2002 2563 2005
rect 10225 2002 10291 2005
rect 2497 2000 10291 2002
rect 2497 1944 2502 2000
rect 2558 1944 10230 2000
rect 10286 1944 10291 2000
rect 2497 1942 10291 1944
rect 2497 1939 2563 1942
rect 10225 1939 10291 1942
rect 20161 1322 20227 1325
rect 20161 1320 22202 1322
rect 20161 1264 20166 1320
rect 20222 1264 22202 1320
rect 20161 1262 22202 1264
rect 20161 1259 20227 1262
rect 22142 808 22202 1262
rect 0 688 480 808
rect 22066 688 22546 808
rect 6361 98 6427 101
rect 14273 98 14339 101
rect 6361 96 14339 98
rect 6361 40 6366 96
rect 6422 40 14278 96
rect 14334 40 14339 96
rect 6361 38 14339 40
rect 6361 35 6427 38
rect 14273 35 14339 38
<< via3 >>
rect 8467 22332 8531 22336
rect 8467 22276 8471 22332
rect 8471 22276 8527 22332
rect 8527 22276 8531 22332
rect 8467 22272 8531 22276
rect 8547 22332 8611 22336
rect 8547 22276 8551 22332
rect 8551 22276 8607 22332
rect 8607 22276 8611 22332
rect 8547 22272 8611 22276
rect 8627 22332 8691 22336
rect 8627 22276 8631 22332
rect 8631 22276 8687 22332
rect 8687 22276 8691 22332
rect 8627 22272 8691 22276
rect 8707 22332 8771 22336
rect 8707 22276 8711 22332
rect 8711 22276 8767 22332
rect 8767 22276 8771 22332
rect 8707 22272 8771 22276
rect 15982 22332 16046 22336
rect 15982 22276 15986 22332
rect 15986 22276 16042 22332
rect 16042 22276 16046 22332
rect 15982 22272 16046 22276
rect 16062 22332 16126 22336
rect 16062 22276 16066 22332
rect 16066 22276 16122 22332
rect 16122 22276 16126 22332
rect 16062 22272 16126 22276
rect 16142 22332 16206 22336
rect 16142 22276 16146 22332
rect 16146 22276 16202 22332
rect 16202 22276 16206 22332
rect 16142 22272 16206 22276
rect 16222 22332 16286 22336
rect 16222 22276 16226 22332
rect 16226 22276 16282 22332
rect 16282 22276 16286 22332
rect 16222 22272 16286 22276
rect 4709 21788 4773 21792
rect 4709 21732 4713 21788
rect 4713 21732 4769 21788
rect 4769 21732 4773 21788
rect 4709 21728 4773 21732
rect 4789 21788 4853 21792
rect 4789 21732 4793 21788
rect 4793 21732 4849 21788
rect 4849 21732 4853 21788
rect 4789 21728 4853 21732
rect 4869 21788 4933 21792
rect 4869 21732 4873 21788
rect 4873 21732 4929 21788
rect 4929 21732 4933 21788
rect 4869 21728 4933 21732
rect 4949 21788 5013 21792
rect 4949 21732 4953 21788
rect 4953 21732 5009 21788
rect 5009 21732 5013 21788
rect 4949 21728 5013 21732
rect 12225 21788 12289 21792
rect 12225 21732 12229 21788
rect 12229 21732 12285 21788
rect 12285 21732 12289 21788
rect 12225 21728 12289 21732
rect 12305 21788 12369 21792
rect 12305 21732 12309 21788
rect 12309 21732 12365 21788
rect 12365 21732 12369 21788
rect 12305 21728 12369 21732
rect 12385 21788 12449 21792
rect 12385 21732 12389 21788
rect 12389 21732 12445 21788
rect 12445 21732 12449 21788
rect 12385 21728 12449 21732
rect 12465 21788 12529 21792
rect 12465 21732 12469 21788
rect 12469 21732 12525 21788
rect 12525 21732 12529 21788
rect 12465 21728 12529 21732
rect 19740 21788 19804 21792
rect 19740 21732 19744 21788
rect 19744 21732 19800 21788
rect 19800 21732 19804 21788
rect 19740 21728 19804 21732
rect 19820 21788 19884 21792
rect 19820 21732 19824 21788
rect 19824 21732 19880 21788
rect 19880 21732 19884 21788
rect 19820 21728 19884 21732
rect 19900 21788 19964 21792
rect 19900 21732 19904 21788
rect 19904 21732 19960 21788
rect 19960 21732 19964 21788
rect 19900 21728 19964 21732
rect 19980 21788 20044 21792
rect 19980 21732 19984 21788
rect 19984 21732 20040 21788
rect 20040 21732 20044 21788
rect 19980 21728 20044 21732
rect 8467 21244 8531 21248
rect 8467 21188 8471 21244
rect 8471 21188 8527 21244
rect 8527 21188 8531 21244
rect 8467 21184 8531 21188
rect 8547 21244 8611 21248
rect 8547 21188 8551 21244
rect 8551 21188 8607 21244
rect 8607 21188 8611 21244
rect 8547 21184 8611 21188
rect 8627 21244 8691 21248
rect 8627 21188 8631 21244
rect 8631 21188 8687 21244
rect 8687 21188 8691 21244
rect 8627 21184 8691 21188
rect 8707 21244 8771 21248
rect 8707 21188 8711 21244
rect 8711 21188 8767 21244
rect 8767 21188 8771 21244
rect 8707 21184 8771 21188
rect 15982 21244 16046 21248
rect 15982 21188 15986 21244
rect 15986 21188 16042 21244
rect 16042 21188 16046 21244
rect 15982 21184 16046 21188
rect 16062 21244 16126 21248
rect 16062 21188 16066 21244
rect 16066 21188 16122 21244
rect 16122 21188 16126 21244
rect 16062 21184 16126 21188
rect 16142 21244 16206 21248
rect 16142 21188 16146 21244
rect 16146 21188 16202 21244
rect 16202 21188 16206 21244
rect 16142 21184 16206 21188
rect 16222 21244 16286 21248
rect 16222 21188 16226 21244
rect 16226 21188 16282 21244
rect 16282 21188 16286 21244
rect 16222 21184 16286 21188
rect 4709 20700 4773 20704
rect 4709 20644 4713 20700
rect 4713 20644 4769 20700
rect 4769 20644 4773 20700
rect 4709 20640 4773 20644
rect 4789 20700 4853 20704
rect 4789 20644 4793 20700
rect 4793 20644 4849 20700
rect 4849 20644 4853 20700
rect 4789 20640 4853 20644
rect 4869 20700 4933 20704
rect 4869 20644 4873 20700
rect 4873 20644 4929 20700
rect 4929 20644 4933 20700
rect 4869 20640 4933 20644
rect 4949 20700 5013 20704
rect 4949 20644 4953 20700
rect 4953 20644 5009 20700
rect 5009 20644 5013 20700
rect 4949 20640 5013 20644
rect 12225 20700 12289 20704
rect 12225 20644 12229 20700
rect 12229 20644 12285 20700
rect 12285 20644 12289 20700
rect 12225 20640 12289 20644
rect 12305 20700 12369 20704
rect 12305 20644 12309 20700
rect 12309 20644 12365 20700
rect 12365 20644 12369 20700
rect 12305 20640 12369 20644
rect 12385 20700 12449 20704
rect 12385 20644 12389 20700
rect 12389 20644 12445 20700
rect 12445 20644 12449 20700
rect 12385 20640 12449 20644
rect 12465 20700 12529 20704
rect 12465 20644 12469 20700
rect 12469 20644 12525 20700
rect 12525 20644 12529 20700
rect 12465 20640 12529 20644
rect 19740 20700 19804 20704
rect 19740 20644 19744 20700
rect 19744 20644 19800 20700
rect 19800 20644 19804 20700
rect 19740 20640 19804 20644
rect 19820 20700 19884 20704
rect 19820 20644 19824 20700
rect 19824 20644 19880 20700
rect 19880 20644 19884 20700
rect 19820 20640 19884 20644
rect 19900 20700 19964 20704
rect 19900 20644 19904 20700
rect 19904 20644 19960 20700
rect 19960 20644 19964 20700
rect 19900 20640 19964 20644
rect 19980 20700 20044 20704
rect 19980 20644 19984 20700
rect 19984 20644 20040 20700
rect 20040 20644 20044 20700
rect 19980 20640 20044 20644
rect 8467 20156 8531 20160
rect 8467 20100 8471 20156
rect 8471 20100 8527 20156
rect 8527 20100 8531 20156
rect 8467 20096 8531 20100
rect 8547 20156 8611 20160
rect 8547 20100 8551 20156
rect 8551 20100 8607 20156
rect 8607 20100 8611 20156
rect 8547 20096 8611 20100
rect 8627 20156 8691 20160
rect 8627 20100 8631 20156
rect 8631 20100 8687 20156
rect 8687 20100 8691 20156
rect 8627 20096 8691 20100
rect 8707 20156 8771 20160
rect 8707 20100 8711 20156
rect 8711 20100 8767 20156
rect 8767 20100 8771 20156
rect 8707 20096 8771 20100
rect 15982 20156 16046 20160
rect 15982 20100 15986 20156
rect 15986 20100 16042 20156
rect 16042 20100 16046 20156
rect 15982 20096 16046 20100
rect 16062 20156 16126 20160
rect 16062 20100 16066 20156
rect 16066 20100 16122 20156
rect 16122 20100 16126 20156
rect 16062 20096 16126 20100
rect 16142 20156 16206 20160
rect 16142 20100 16146 20156
rect 16146 20100 16202 20156
rect 16202 20100 16206 20156
rect 16142 20096 16206 20100
rect 16222 20156 16286 20160
rect 16222 20100 16226 20156
rect 16226 20100 16282 20156
rect 16282 20100 16286 20156
rect 16222 20096 16286 20100
rect 4709 19612 4773 19616
rect 4709 19556 4713 19612
rect 4713 19556 4769 19612
rect 4769 19556 4773 19612
rect 4709 19552 4773 19556
rect 4789 19612 4853 19616
rect 4789 19556 4793 19612
rect 4793 19556 4849 19612
rect 4849 19556 4853 19612
rect 4789 19552 4853 19556
rect 4869 19612 4933 19616
rect 4869 19556 4873 19612
rect 4873 19556 4929 19612
rect 4929 19556 4933 19612
rect 4869 19552 4933 19556
rect 4949 19612 5013 19616
rect 4949 19556 4953 19612
rect 4953 19556 5009 19612
rect 5009 19556 5013 19612
rect 4949 19552 5013 19556
rect 12225 19612 12289 19616
rect 12225 19556 12229 19612
rect 12229 19556 12285 19612
rect 12285 19556 12289 19612
rect 12225 19552 12289 19556
rect 12305 19612 12369 19616
rect 12305 19556 12309 19612
rect 12309 19556 12365 19612
rect 12365 19556 12369 19612
rect 12305 19552 12369 19556
rect 12385 19612 12449 19616
rect 12385 19556 12389 19612
rect 12389 19556 12445 19612
rect 12445 19556 12449 19612
rect 12385 19552 12449 19556
rect 12465 19612 12529 19616
rect 12465 19556 12469 19612
rect 12469 19556 12525 19612
rect 12525 19556 12529 19612
rect 12465 19552 12529 19556
rect 19740 19612 19804 19616
rect 19740 19556 19744 19612
rect 19744 19556 19800 19612
rect 19800 19556 19804 19612
rect 19740 19552 19804 19556
rect 19820 19612 19884 19616
rect 19820 19556 19824 19612
rect 19824 19556 19880 19612
rect 19880 19556 19884 19612
rect 19820 19552 19884 19556
rect 19900 19612 19964 19616
rect 19900 19556 19904 19612
rect 19904 19556 19960 19612
rect 19960 19556 19964 19612
rect 19900 19552 19964 19556
rect 19980 19612 20044 19616
rect 19980 19556 19984 19612
rect 19984 19556 20040 19612
rect 20040 19556 20044 19612
rect 19980 19552 20044 19556
rect 8467 19068 8531 19072
rect 8467 19012 8471 19068
rect 8471 19012 8527 19068
rect 8527 19012 8531 19068
rect 8467 19008 8531 19012
rect 8547 19068 8611 19072
rect 8547 19012 8551 19068
rect 8551 19012 8607 19068
rect 8607 19012 8611 19068
rect 8547 19008 8611 19012
rect 8627 19068 8691 19072
rect 8627 19012 8631 19068
rect 8631 19012 8687 19068
rect 8687 19012 8691 19068
rect 8627 19008 8691 19012
rect 8707 19068 8771 19072
rect 8707 19012 8711 19068
rect 8711 19012 8767 19068
rect 8767 19012 8771 19068
rect 8707 19008 8771 19012
rect 15982 19068 16046 19072
rect 15982 19012 15986 19068
rect 15986 19012 16042 19068
rect 16042 19012 16046 19068
rect 15982 19008 16046 19012
rect 16062 19068 16126 19072
rect 16062 19012 16066 19068
rect 16066 19012 16122 19068
rect 16122 19012 16126 19068
rect 16062 19008 16126 19012
rect 16142 19068 16206 19072
rect 16142 19012 16146 19068
rect 16146 19012 16202 19068
rect 16202 19012 16206 19068
rect 16142 19008 16206 19012
rect 16222 19068 16286 19072
rect 16222 19012 16226 19068
rect 16226 19012 16282 19068
rect 16282 19012 16286 19068
rect 16222 19008 16286 19012
rect 4709 18524 4773 18528
rect 4709 18468 4713 18524
rect 4713 18468 4769 18524
rect 4769 18468 4773 18524
rect 4709 18464 4773 18468
rect 4789 18524 4853 18528
rect 4789 18468 4793 18524
rect 4793 18468 4849 18524
rect 4849 18468 4853 18524
rect 4789 18464 4853 18468
rect 4869 18524 4933 18528
rect 4869 18468 4873 18524
rect 4873 18468 4929 18524
rect 4929 18468 4933 18524
rect 4869 18464 4933 18468
rect 4949 18524 5013 18528
rect 4949 18468 4953 18524
rect 4953 18468 5009 18524
rect 5009 18468 5013 18524
rect 4949 18464 5013 18468
rect 12225 18524 12289 18528
rect 12225 18468 12229 18524
rect 12229 18468 12285 18524
rect 12285 18468 12289 18524
rect 12225 18464 12289 18468
rect 12305 18524 12369 18528
rect 12305 18468 12309 18524
rect 12309 18468 12365 18524
rect 12365 18468 12369 18524
rect 12305 18464 12369 18468
rect 12385 18524 12449 18528
rect 12385 18468 12389 18524
rect 12389 18468 12445 18524
rect 12445 18468 12449 18524
rect 12385 18464 12449 18468
rect 12465 18524 12529 18528
rect 12465 18468 12469 18524
rect 12469 18468 12525 18524
rect 12525 18468 12529 18524
rect 12465 18464 12529 18468
rect 19740 18524 19804 18528
rect 19740 18468 19744 18524
rect 19744 18468 19800 18524
rect 19800 18468 19804 18524
rect 19740 18464 19804 18468
rect 19820 18524 19884 18528
rect 19820 18468 19824 18524
rect 19824 18468 19880 18524
rect 19880 18468 19884 18524
rect 19820 18464 19884 18468
rect 19900 18524 19964 18528
rect 19900 18468 19904 18524
rect 19904 18468 19960 18524
rect 19960 18468 19964 18524
rect 19900 18464 19964 18468
rect 19980 18524 20044 18528
rect 19980 18468 19984 18524
rect 19984 18468 20040 18524
rect 20040 18468 20044 18524
rect 19980 18464 20044 18468
rect 8467 17980 8531 17984
rect 8467 17924 8471 17980
rect 8471 17924 8527 17980
rect 8527 17924 8531 17980
rect 8467 17920 8531 17924
rect 8547 17980 8611 17984
rect 8547 17924 8551 17980
rect 8551 17924 8607 17980
rect 8607 17924 8611 17980
rect 8547 17920 8611 17924
rect 8627 17980 8691 17984
rect 8627 17924 8631 17980
rect 8631 17924 8687 17980
rect 8687 17924 8691 17980
rect 8627 17920 8691 17924
rect 8707 17980 8771 17984
rect 8707 17924 8711 17980
rect 8711 17924 8767 17980
rect 8767 17924 8771 17980
rect 8707 17920 8771 17924
rect 15982 17980 16046 17984
rect 15982 17924 15986 17980
rect 15986 17924 16042 17980
rect 16042 17924 16046 17980
rect 15982 17920 16046 17924
rect 16062 17980 16126 17984
rect 16062 17924 16066 17980
rect 16066 17924 16122 17980
rect 16122 17924 16126 17980
rect 16062 17920 16126 17924
rect 16142 17980 16206 17984
rect 16142 17924 16146 17980
rect 16146 17924 16202 17980
rect 16202 17924 16206 17980
rect 16142 17920 16206 17924
rect 16222 17980 16286 17984
rect 16222 17924 16226 17980
rect 16226 17924 16282 17980
rect 16282 17924 16286 17980
rect 16222 17920 16286 17924
rect 4709 17436 4773 17440
rect 4709 17380 4713 17436
rect 4713 17380 4769 17436
rect 4769 17380 4773 17436
rect 4709 17376 4773 17380
rect 4789 17436 4853 17440
rect 4789 17380 4793 17436
rect 4793 17380 4849 17436
rect 4849 17380 4853 17436
rect 4789 17376 4853 17380
rect 4869 17436 4933 17440
rect 4869 17380 4873 17436
rect 4873 17380 4929 17436
rect 4929 17380 4933 17436
rect 4869 17376 4933 17380
rect 4949 17436 5013 17440
rect 4949 17380 4953 17436
rect 4953 17380 5009 17436
rect 5009 17380 5013 17436
rect 4949 17376 5013 17380
rect 12225 17436 12289 17440
rect 12225 17380 12229 17436
rect 12229 17380 12285 17436
rect 12285 17380 12289 17436
rect 12225 17376 12289 17380
rect 12305 17436 12369 17440
rect 12305 17380 12309 17436
rect 12309 17380 12365 17436
rect 12365 17380 12369 17436
rect 12305 17376 12369 17380
rect 12385 17436 12449 17440
rect 12385 17380 12389 17436
rect 12389 17380 12445 17436
rect 12445 17380 12449 17436
rect 12385 17376 12449 17380
rect 12465 17436 12529 17440
rect 12465 17380 12469 17436
rect 12469 17380 12525 17436
rect 12525 17380 12529 17436
rect 12465 17376 12529 17380
rect 19740 17436 19804 17440
rect 19740 17380 19744 17436
rect 19744 17380 19800 17436
rect 19800 17380 19804 17436
rect 19740 17376 19804 17380
rect 19820 17436 19884 17440
rect 19820 17380 19824 17436
rect 19824 17380 19880 17436
rect 19880 17380 19884 17436
rect 19820 17376 19884 17380
rect 19900 17436 19964 17440
rect 19900 17380 19904 17436
rect 19904 17380 19960 17436
rect 19960 17380 19964 17436
rect 19900 17376 19964 17380
rect 19980 17436 20044 17440
rect 19980 17380 19984 17436
rect 19984 17380 20040 17436
rect 20040 17380 20044 17436
rect 19980 17376 20044 17380
rect 8467 16892 8531 16896
rect 8467 16836 8471 16892
rect 8471 16836 8527 16892
rect 8527 16836 8531 16892
rect 8467 16832 8531 16836
rect 8547 16892 8611 16896
rect 8547 16836 8551 16892
rect 8551 16836 8607 16892
rect 8607 16836 8611 16892
rect 8547 16832 8611 16836
rect 8627 16892 8691 16896
rect 8627 16836 8631 16892
rect 8631 16836 8687 16892
rect 8687 16836 8691 16892
rect 8627 16832 8691 16836
rect 8707 16892 8771 16896
rect 8707 16836 8711 16892
rect 8711 16836 8767 16892
rect 8767 16836 8771 16892
rect 8707 16832 8771 16836
rect 15982 16892 16046 16896
rect 15982 16836 15986 16892
rect 15986 16836 16042 16892
rect 16042 16836 16046 16892
rect 15982 16832 16046 16836
rect 16062 16892 16126 16896
rect 16062 16836 16066 16892
rect 16066 16836 16122 16892
rect 16122 16836 16126 16892
rect 16062 16832 16126 16836
rect 16142 16892 16206 16896
rect 16142 16836 16146 16892
rect 16146 16836 16202 16892
rect 16202 16836 16206 16892
rect 16142 16832 16206 16836
rect 16222 16892 16286 16896
rect 16222 16836 16226 16892
rect 16226 16836 16282 16892
rect 16282 16836 16286 16892
rect 16222 16832 16286 16836
rect 4709 16348 4773 16352
rect 4709 16292 4713 16348
rect 4713 16292 4769 16348
rect 4769 16292 4773 16348
rect 4709 16288 4773 16292
rect 4789 16348 4853 16352
rect 4789 16292 4793 16348
rect 4793 16292 4849 16348
rect 4849 16292 4853 16348
rect 4789 16288 4853 16292
rect 4869 16348 4933 16352
rect 4869 16292 4873 16348
rect 4873 16292 4929 16348
rect 4929 16292 4933 16348
rect 4869 16288 4933 16292
rect 4949 16348 5013 16352
rect 4949 16292 4953 16348
rect 4953 16292 5009 16348
rect 5009 16292 5013 16348
rect 4949 16288 5013 16292
rect 12225 16348 12289 16352
rect 12225 16292 12229 16348
rect 12229 16292 12285 16348
rect 12285 16292 12289 16348
rect 12225 16288 12289 16292
rect 12305 16348 12369 16352
rect 12305 16292 12309 16348
rect 12309 16292 12365 16348
rect 12365 16292 12369 16348
rect 12305 16288 12369 16292
rect 12385 16348 12449 16352
rect 12385 16292 12389 16348
rect 12389 16292 12445 16348
rect 12445 16292 12449 16348
rect 12385 16288 12449 16292
rect 12465 16348 12529 16352
rect 12465 16292 12469 16348
rect 12469 16292 12525 16348
rect 12525 16292 12529 16348
rect 12465 16288 12529 16292
rect 19740 16348 19804 16352
rect 19740 16292 19744 16348
rect 19744 16292 19800 16348
rect 19800 16292 19804 16348
rect 19740 16288 19804 16292
rect 19820 16348 19884 16352
rect 19820 16292 19824 16348
rect 19824 16292 19880 16348
rect 19880 16292 19884 16348
rect 19820 16288 19884 16292
rect 19900 16348 19964 16352
rect 19900 16292 19904 16348
rect 19904 16292 19960 16348
rect 19960 16292 19964 16348
rect 19900 16288 19964 16292
rect 19980 16348 20044 16352
rect 19980 16292 19984 16348
rect 19984 16292 20040 16348
rect 20040 16292 20044 16348
rect 19980 16288 20044 16292
rect 8467 15804 8531 15808
rect 8467 15748 8471 15804
rect 8471 15748 8527 15804
rect 8527 15748 8531 15804
rect 8467 15744 8531 15748
rect 8547 15804 8611 15808
rect 8547 15748 8551 15804
rect 8551 15748 8607 15804
rect 8607 15748 8611 15804
rect 8547 15744 8611 15748
rect 8627 15804 8691 15808
rect 8627 15748 8631 15804
rect 8631 15748 8687 15804
rect 8687 15748 8691 15804
rect 8627 15744 8691 15748
rect 8707 15804 8771 15808
rect 8707 15748 8711 15804
rect 8711 15748 8767 15804
rect 8767 15748 8771 15804
rect 8707 15744 8771 15748
rect 15982 15804 16046 15808
rect 15982 15748 15986 15804
rect 15986 15748 16042 15804
rect 16042 15748 16046 15804
rect 15982 15744 16046 15748
rect 16062 15804 16126 15808
rect 16062 15748 16066 15804
rect 16066 15748 16122 15804
rect 16122 15748 16126 15804
rect 16062 15744 16126 15748
rect 16142 15804 16206 15808
rect 16142 15748 16146 15804
rect 16146 15748 16202 15804
rect 16202 15748 16206 15804
rect 16142 15744 16206 15748
rect 16222 15804 16286 15808
rect 16222 15748 16226 15804
rect 16226 15748 16282 15804
rect 16282 15748 16286 15804
rect 16222 15744 16286 15748
rect 4709 15260 4773 15264
rect 4709 15204 4713 15260
rect 4713 15204 4769 15260
rect 4769 15204 4773 15260
rect 4709 15200 4773 15204
rect 4789 15260 4853 15264
rect 4789 15204 4793 15260
rect 4793 15204 4849 15260
rect 4849 15204 4853 15260
rect 4789 15200 4853 15204
rect 4869 15260 4933 15264
rect 4869 15204 4873 15260
rect 4873 15204 4929 15260
rect 4929 15204 4933 15260
rect 4869 15200 4933 15204
rect 4949 15260 5013 15264
rect 4949 15204 4953 15260
rect 4953 15204 5009 15260
rect 5009 15204 5013 15260
rect 4949 15200 5013 15204
rect 12225 15260 12289 15264
rect 12225 15204 12229 15260
rect 12229 15204 12285 15260
rect 12285 15204 12289 15260
rect 12225 15200 12289 15204
rect 12305 15260 12369 15264
rect 12305 15204 12309 15260
rect 12309 15204 12365 15260
rect 12365 15204 12369 15260
rect 12305 15200 12369 15204
rect 12385 15260 12449 15264
rect 12385 15204 12389 15260
rect 12389 15204 12445 15260
rect 12445 15204 12449 15260
rect 12385 15200 12449 15204
rect 12465 15260 12529 15264
rect 12465 15204 12469 15260
rect 12469 15204 12525 15260
rect 12525 15204 12529 15260
rect 12465 15200 12529 15204
rect 19740 15260 19804 15264
rect 19740 15204 19744 15260
rect 19744 15204 19800 15260
rect 19800 15204 19804 15260
rect 19740 15200 19804 15204
rect 19820 15260 19884 15264
rect 19820 15204 19824 15260
rect 19824 15204 19880 15260
rect 19880 15204 19884 15260
rect 19820 15200 19884 15204
rect 19900 15260 19964 15264
rect 19900 15204 19904 15260
rect 19904 15204 19960 15260
rect 19960 15204 19964 15260
rect 19900 15200 19964 15204
rect 19980 15260 20044 15264
rect 19980 15204 19984 15260
rect 19984 15204 20040 15260
rect 20040 15204 20044 15260
rect 19980 15200 20044 15204
rect 60 14860 124 14924
rect 8467 14716 8531 14720
rect 8467 14660 8471 14716
rect 8471 14660 8527 14716
rect 8527 14660 8531 14716
rect 8467 14656 8531 14660
rect 8547 14716 8611 14720
rect 8547 14660 8551 14716
rect 8551 14660 8607 14716
rect 8607 14660 8611 14716
rect 8547 14656 8611 14660
rect 8627 14716 8691 14720
rect 8627 14660 8631 14716
rect 8631 14660 8687 14716
rect 8687 14660 8691 14716
rect 8627 14656 8691 14660
rect 8707 14716 8771 14720
rect 8707 14660 8711 14716
rect 8711 14660 8767 14716
rect 8767 14660 8771 14716
rect 8707 14656 8771 14660
rect 15982 14716 16046 14720
rect 15982 14660 15986 14716
rect 15986 14660 16042 14716
rect 16042 14660 16046 14716
rect 15982 14656 16046 14660
rect 16062 14716 16126 14720
rect 16062 14660 16066 14716
rect 16066 14660 16122 14716
rect 16122 14660 16126 14716
rect 16062 14656 16126 14660
rect 16142 14716 16206 14720
rect 16142 14660 16146 14716
rect 16146 14660 16202 14716
rect 16202 14660 16206 14716
rect 16142 14656 16206 14660
rect 16222 14716 16286 14720
rect 16222 14660 16226 14716
rect 16226 14660 16282 14716
rect 16282 14660 16286 14716
rect 16222 14656 16286 14660
rect 22140 14588 22204 14652
rect 60 14452 124 14516
rect 22140 14316 22204 14380
rect 4709 14172 4773 14176
rect 4709 14116 4713 14172
rect 4713 14116 4769 14172
rect 4769 14116 4773 14172
rect 4709 14112 4773 14116
rect 4789 14172 4853 14176
rect 4789 14116 4793 14172
rect 4793 14116 4849 14172
rect 4849 14116 4853 14172
rect 4789 14112 4853 14116
rect 4869 14172 4933 14176
rect 4869 14116 4873 14172
rect 4873 14116 4929 14172
rect 4929 14116 4933 14172
rect 4869 14112 4933 14116
rect 4949 14172 5013 14176
rect 4949 14116 4953 14172
rect 4953 14116 5009 14172
rect 5009 14116 5013 14172
rect 4949 14112 5013 14116
rect 12225 14172 12289 14176
rect 12225 14116 12229 14172
rect 12229 14116 12285 14172
rect 12285 14116 12289 14172
rect 12225 14112 12289 14116
rect 12305 14172 12369 14176
rect 12305 14116 12309 14172
rect 12309 14116 12365 14172
rect 12365 14116 12369 14172
rect 12305 14112 12369 14116
rect 12385 14172 12449 14176
rect 12385 14116 12389 14172
rect 12389 14116 12445 14172
rect 12445 14116 12449 14172
rect 12385 14112 12449 14116
rect 12465 14172 12529 14176
rect 12465 14116 12469 14172
rect 12469 14116 12525 14172
rect 12525 14116 12529 14172
rect 12465 14112 12529 14116
rect 19740 14172 19804 14176
rect 19740 14116 19744 14172
rect 19744 14116 19800 14172
rect 19800 14116 19804 14172
rect 19740 14112 19804 14116
rect 19820 14172 19884 14176
rect 19820 14116 19824 14172
rect 19824 14116 19880 14172
rect 19880 14116 19884 14172
rect 19820 14112 19884 14116
rect 19900 14172 19964 14176
rect 19900 14116 19904 14172
rect 19904 14116 19960 14172
rect 19960 14116 19964 14172
rect 19900 14112 19964 14116
rect 19980 14172 20044 14176
rect 19980 14116 19984 14172
rect 19984 14116 20040 14172
rect 20040 14116 20044 14172
rect 19980 14112 20044 14116
rect 8467 13628 8531 13632
rect 8467 13572 8471 13628
rect 8471 13572 8527 13628
rect 8527 13572 8531 13628
rect 8467 13568 8531 13572
rect 8547 13628 8611 13632
rect 8547 13572 8551 13628
rect 8551 13572 8607 13628
rect 8607 13572 8611 13628
rect 8547 13568 8611 13572
rect 8627 13628 8691 13632
rect 8627 13572 8631 13628
rect 8631 13572 8687 13628
rect 8687 13572 8691 13628
rect 8627 13568 8691 13572
rect 8707 13628 8771 13632
rect 8707 13572 8711 13628
rect 8711 13572 8767 13628
rect 8767 13572 8771 13628
rect 8707 13568 8771 13572
rect 15982 13628 16046 13632
rect 15982 13572 15986 13628
rect 15986 13572 16042 13628
rect 16042 13572 16046 13628
rect 15982 13568 16046 13572
rect 16062 13628 16126 13632
rect 16062 13572 16066 13628
rect 16066 13572 16122 13628
rect 16122 13572 16126 13628
rect 16062 13568 16126 13572
rect 16142 13628 16206 13632
rect 16142 13572 16146 13628
rect 16146 13572 16202 13628
rect 16202 13572 16206 13628
rect 16142 13568 16206 13572
rect 16222 13628 16286 13632
rect 16222 13572 16226 13628
rect 16226 13572 16282 13628
rect 16282 13572 16286 13628
rect 16222 13568 16286 13572
rect 4709 13084 4773 13088
rect 4709 13028 4713 13084
rect 4713 13028 4769 13084
rect 4769 13028 4773 13084
rect 4709 13024 4773 13028
rect 4789 13084 4853 13088
rect 4789 13028 4793 13084
rect 4793 13028 4849 13084
rect 4849 13028 4853 13084
rect 4789 13024 4853 13028
rect 4869 13084 4933 13088
rect 4869 13028 4873 13084
rect 4873 13028 4929 13084
rect 4929 13028 4933 13084
rect 4869 13024 4933 13028
rect 4949 13084 5013 13088
rect 4949 13028 4953 13084
rect 4953 13028 5009 13084
rect 5009 13028 5013 13084
rect 4949 13024 5013 13028
rect 12225 13084 12289 13088
rect 12225 13028 12229 13084
rect 12229 13028 12285 13084
rect 12285 13028 12289 13084
rect 12225 13024 12289 13028
rect 12305 13084 12369 13088
rect 12305 13028 12309 13084
rect 12309 13028 12365 13084
rect 12365 13028 12369 13084
rect 12305 13024 12369 13028
rect 12385 13084 12449 13088
rect 12385 13028 12389 13084
rect 12389 13028 12445 13084
rect 12445 13028 12449 13084
rect 12385 13024 12449 13028
rect 12465 13084 12529 13088
rect 12465 13028 12469 13084
rect 12469 13028 12525 13084
rect 12525 13028 12529 13084
rect 12465 13024 12529 13028
rect 19740 13084 19804 13088
rect 19740 13028 19744 13084
rect 19744 13028 19800 13084
rect 19800 13028 19804 13084
rect 19740 13024 19804 13028
rect 19820 13084 19884 13088
rect 19820 13028 19824 13084
rect 19824 13028 19880 13084
rect 19880 13028 19884 13084
rect 19820 13024 19884 13028
rect 19900 13084 19964 13088
rect 19900 13028 19904 13084
rect 19904 13028 19960 13084
rect 19960 13028 19964 13084
rect 19900 13024 19964 13028
rect 19980 13084 20044 13088
rect 19980 13028 19984 13084
rect 19984 13028 20040 13084
rect 20040 13028 20044 13084
rect 19980 13024 20044 13028
rect 8467 12540 8531 12544
rect 8467 12484 8471 12540
rect 8471 12484 8527 12540
rect 8527 12484 8531 12540
rect 8467 12480 8531 12484
rect 8547 12540 8611 12544
rect 8547 12484 8551 12540
rect 8551 12484 8607 12540
rect 8607 12484 8611 12540
rect 8547 12480 8611 12484
rect 8627 12540 8691 12544
rect 8627 12484 8631 12540
rect 8631 12484 8687 12540
rect 8687 12484 8691 12540
rect 8627 12480 8691 12484
rect 8707 12540 8771 12544
rect 8707 12484 8711 12540
rect 8711 12484 8767 12540
rect 8767 12484 8771 12540
rect 8707 12480 8771 12484
rect 15982 12540 16046 12544
rect 15982 12484 15986 12540
rect 15986 12484 16042 12540
rect 16042 12484 16046 12540
rect 15982 12480 16046 12484
rect 16062 12540 16126 12544
rect 16062 12484 16066 12540
rect 16066 12484 16122 12540
rect 16122 12484 16126 12540
rect 16062 12480 16126 12484
rect 16142 12540 16206 12544
rect 16142 12484 16146 12540
rect 16146 12484 16202 12540
rect 16202 12484 16206 12540
rect 16142 12480 16206 12484
rect 16222 12540 16286 12544
rect 16222 12484 16226 12540
rect 16226 12484 16282 12540
rect 16282 12484 16286 12540
rect 16222 12480 16286 12484
rect 4709 11996 4773 12000
rect 4709 11940 4713 11996
rect 4713 11940 4769 11996
rect 4769 11940 4773 11996
rect 4709 11936 4773 11940
rect 4789 11996 4853 12000
rect 4789 11940 4793 11996
rect 4793 11940 4849 11996
rect 4849 11940 4853 11996
rect 4789 11936 4853 11940
rect 4869 11996 4933 12000
rect 4869 11940 4873 11996
rect 4873 11940 4929 11996
rect 4929 11940 4933 11996
rect 4869 11936 4933 11940
rect 4949 11996 5013 12000
rect 4949 11940 4953 11996
rect 4953 11940 5009 11996
rect 5009 11940 5013 11996
rect 4949 11936 5013 11940
rect 12225 11996 12289 12000
rect 12225 11940 12229 11996
rect 12229 11940 12285 11996
rect 12285 11940 12289 11996
rect 12225 11936 12289 11940
rect 12305 11996 12369 12000
rect 12305 11940 12309 11996
rect 12309 11940 12365 11996
rect 12365 11940 12369 11996
rect 12305 11936 12369 11940
rect 12385 11996 12449 12000
rect 12385 11940 12389 11996
rect 12389 11940 12445 11996
rect 12445 11940 12449 11996
rect 12385 11936 12449 11940
rect 12465 11996 12529 12000
rect 12465 11940 12469 11996
rect 12469 11940 12525 11996
rect 12525 11940 12529 11996
rect 12465 11936 12529 11940
rect 19740 11996 19804 12000
rect 19740 11940 19744 11996
rect 19744 11940 19800 11996
rect 19800 11940 19804 11996
rect 19740 11936 19804 11940
rect 19820 11996 19884 12000
rect 19820 11940 19824 11996
rect 19824 11940 19880 11996
rect 19880 11940 19884 11996
rect 19820 11936 19884 11940
rect 19900 11996 19964 12000
rect 19900 11940 19904 11996
rect 19904 11940 19960 11996
rect 19960 11940 19964 11996
rect 19900 11936 19964 11940
rect 19980 11996 20044 12000
rect 19980 11940 19984 11996
rect 19984 11940 20040 11996
rect 20040 11940 20044 11996
rect 19980 11936 20044 11940
rect 8467 11452 8531 11456
rect 8467 11396 8471 11452
rect 8471 11396 8527 11452
rect 8527 11396 8531 11452
rect 8467 11392 8531 11396
rect 8547 11452 8611 11456
rect 8547 11396 8551 11452
rect 8551 11396 8607 11452
rect 8607 11396 8611 11452
rect 8547 11392 8611 11396
rect 8627 11452 8691 11456
rect 8627 11396 8631 11452
rect 8631 11396 8687 11452
rect 8687 11396 8691 11452
rect 8627 11392 8691 11396
rect 8707 11452 8771 11456
rect 8707 11396 8711 11452
rect 8711 11396 8767 11452
rect 8767 11396 8771 11452
rect 8707 11392 8771 11396
rect 15982 11452 16046 11456
rect 15982 11396 15986 11452
rect 15986 11396 16042 11452
rect 16042 11396 16046 11452
rect 15982 11392 16046 11396
rect 16062 11452 16126 11456
rect 16062 11396 16066 11452
rect 16066 11396 16122 11452
rect 16122 11396 16126 11452
rect 16062 11392 16126 11396
rect 16142 11452 16206 11456
rect 16142 11396 16146 11452
rect 16146 11396 16202 11452
rect 16202 11396 16206 11452
rect 16142 11392 16206 11396
rect 16222 11452 16286 11456
rect 16222 11396 16226 11452
rect 16226 11396 16282 11452
rect 16282 11396 16286 11452
rect 16222 11392 16286 11396
rect 4709 10908 4773 10912
rect 4709 10852 4713 10908
rect 4713 10852 4769 10908
rect 4769 10852 4773 10908
rect 4709 10848 4773 10852
rect 4789 10908 4853 10912
rect 4789 10852 4793 10908
rect 4793 10852 4849 10908
rect 4849 10852 4853 10908
rect 4789 10848 4853 10852
rect 4869 10908 4933 10912
rect 4869 10852 4873 10908
rect 4873 10852 4929 10908
rect 4929 10852 4933 10908
rect 4869 10848 4933 10852
rect 4949 10908 5013 10912
rect 4949 10852 4953 10908
rect 4953 10852 5009 10908
rect 5009 10852 5013 10908
rect 4949 10848 5013 10852
rect 12225 10908 12289 10912
rect 12225 10852 12229 10908
rect 12229 10852 12285 10908
rect 12285 10852 12289 10908
rect 12225 10848 12289 10852
rect 12305 10908 12369 10912
rect 12305 10852 12309 10908
rect 12309 10852 12365 10908
rect 12365 10852 12369 10908
rect 12305 10848 12369 10852
rect 12385 10908 12449 10912
rect 12385 10852 12389 10908
rect 12389 10852 12445 10908
rect 12445 10852 12449 10908
rect 12385 10848 12449 10852
rect 12465 10908 12529 10912
rect 12465 10852 12469 10908
rect 12469 10852 12525 10908
rect 12525 10852 12529 10908
rect 12465 10848 12529 10852
rect 19740 10908 19804 10912
rect 19740 10852 19744 10908
rect 19744 10852 19800 10908
rect 19800 10852 19804 10908
rect 19740 10848 19804 10852
rect 19820 10908 19884 10912
rect 19820 10852 19824 10908
rect 19824 10852 19880 10908
rect 19880 10852 19884 10908
rect 19820 10848 19884 10852
rect 19900 10908 19964 10912
rect 19900 10852 19904 10908
rect 19904 10852 19960 10908
rect 19960 10852 19964 10908
rect 19900 10848 19964 10852
rect 19980 10908 20044 10912
rect 19980 10852 19984 10908
rect 19984 10852 20040 10908
rect 20040 10852 20044 10908
rect 19980 10848 20044 10852
rect 8467 10364 8531 10368
rect 8467 10308 8471 10364
rect 8471 10308 8527 10364
rect 8527 10308 8531 10364
rect 8467 10304 8531 10308
rect 8547 10364 8611 10368
rect 8547 10308 8551 10364
rect 8551 10308 8607 10364
rect 8607 10308 8611 10364
rect 8547 10304 8611 10308
rect 8627 10364 8691 10368
rect 8627 10308 8631 10364
rect 8631 10308 8687 10364
rect 8687 10308 8691 10364
rect 8627 10304 8691 10308
rect 8707 10364 8771 10368
rect 8707 10308 8711 10364
rect 8711 10308 8767 10364
rect 8767 10308 8771 10364
rect 8707 10304 8771 10308
rect 15982 10364 16046 10368
rect 15982 10308 15986 10364
rect 15986 10308 16042 10364
rect 16042 10308 16046 10364
rect 15982 10304 16046 10308
rect 16062 10364 16126 10368
rect 16062 10308 16066 10364
rect 16066 10308 16122 10364
rect 16122 10308 16126 10364
rect 16062 10304 16126 10308
rect 16142 10364 16206 10368
rect 16142 10308 16146 10364
rect 16146 10308 16202 10364
rect 16202 10308 16206 10364
rect 16142 10304 16206 10308
rect 16222 10364 16286 10368
rect 16222 10308 16226 10364
rect 16226 10308 16282 10364
rect 16282 10308 16286 10364
rect 16222 10304 16286 10308
rect 4709 9820 4773 9824
rect 4709 9764 4713 9820
rect 4713 9764 4769 9820
rect 4769 9764 4773 9820
rect 4709 9760 4773 9764
rect 4789 9820 4853 9824
rect 4789 9764 4793 9820
rect 4793 9764 4849 9820
rect 4849 9764 4853 9820
rect 4789 9760 4853 9764
rect 4869 9820 4933 9824
rect 4869 9764 4873 9820
rect 4873 9764 4929 9820
rect 4929 9764 4933 9820
rect 4869 9760 4933 9764
rect 4949 9820 5013 9824
rect 4949 9764 4953 9820
rect 4953 9764 5009 9820
rect 5009 9764 5013 9820
rect 4949 9760 5013 9764
rect 12225 9820 12289 9824
rect 12225 9764 12229 9820
rect 12229 9764 12285 9820
rect 12285 9764 12289 9820
rect 12225 9760 12289 9764
rect 12305 9820 12369 9824
rect 12305 9764 12309 9820
rect 12309 9764 12365 9820
rect 12365 9764 12369 9820
rect 12305 9760 12369 9764
rect 12385 9820 12449 9824
rect 12385 9764 12389 9820
rect 12389 9764 12445 9820
rect 12445 9764 12449 9820
rect 12385 9760 12449 9764
rect 12465 9820 12529 9824
rect 12465 9764 12469 9820
rect 12469 9764 12525 9820
rect 12525 9764 12529 9820
rect 12465 9760 12529 9764
rect 19740 9820 19804 9824
rect 19740 9764 19744 9820
rect 19744 9764 19800 9820
rect 19800 9764 19804 9820
rect 19740 9760 19804 9764
rect 19820 9820 19884 9824
rect 19820 9764 19824 9820
rect 19824 9764 19880 9820
rect 19880 9764 19884 9820
rect 19820 9760 19884 9764
rect 19900 9820 19964 9824
rect 19900 9764 19904 9820
rect 19904 9764 19960 9820
rect 19960 9764 19964 9820
rect 19900 9760 19964 9764
rect 19980 9820 20044 9824
rect 19980 9764 19984 9820
rect 19984 9764 20040 9820
rect 20040 9764 20044 9820
rect 19980 9760 20044 9764
rect 8467 9276 8531 9280
rect 8467 9220 8471 9276
rect 8471 9220 8527 9276
rect 8527 9220 8531 9276
rect 8467 9216 8531 9220
rect 8547 9276 8611 9280
rect 8547 9220 8551 9276
rect 8551 9220 8607 9276
rect 8607 9220 8611 9276
rect 8547 9216 8611 9220
rect 8627 9276 8691 9280
rect 8627 9220 8631 9276
rect 8631 9220 8687 9276
rect 8687 9220 8691 9276
rect 8627 9216 8691 9220
rect 8707 9276 8771 9280
rect 8707 9220 8711 9276
rect 8711 9220 8767 9276
rect 8767 9220 8771 9276
rect 8707 9216 8771 9220
rect 15982 9276 16046 9280
rect 15982 9220 15986 9276
rect 15986 9220 16042 9276
rect 16042 9220 16046 9276
rect 15982 9216 16046 9220
rect 16062 9276 16126 9280
rect 16062 9220 16066 9276
rect 16066 9220 16122 9276
rect 16122 9220 16126 9276
rect 16062 9216 16126 9220
rect 16142 9276 16206 9280
rect 16142 9220 16146 9276
rect 16146 9220 16202 9276
rect 16202 9220 16206 9276
rect 16142 9216 16206 9220
rect 16222 9276 16286 9280
rect 16222 9220 16226 9276
rect 16226 9220 16282 9276
rect 16282 9220 16286 9276
rect 16222 9216 16286 9220
rect 4709 8732 4773 8736
rect 4709 8676 4713 8732
rect 4713 8676 4769 8732
rect 4769 8676 4773 8732
rect 4709 8672 4773 8676
rect 4789 8732 4853 8736
rect 4789 8676 4793 8732
rect 4793 8676 4849 8732
rect 4849 8676 4853 8732
rect 4789 8672 4853 8676
rect 4869 8732 4933 8736
rect 4869 8676 4873 8732
rect 4873 8676 4929 8732
rect 4929 8676 4933 8732
rect 4869 8672 4933 8676
rect 4949 8732 5013 8736
rect 4949 8676 4953 8732
rect 4953 8676 5009 8732
rect 5009 8676 5013 8732
rect 4949 8672 5013 8676
rect 12225 8732 12289 8736
rect 12225 8676 12229 8732
rect 12229 8676 12285 8732
rect 12285 8676 12289 8732
rect 12225 8672 12289 8676
rect 12305 8732 12369 8736
rect 12305 8676 12309 8732
rect 12309 8676 12365 8732
rect 12365 8676 12369 8732
rect 12305 8672 12369 8676
rect 12385 8732 12449 8736
rect 12385 8676 12389 8732
rect 12389 8676 12445 8732
rect 12445 8676 12449 8732
rect 12385 8672 12449 8676
rect 12465 8732 12529 8736
rect 12465 8676 12469 8732
rect 12469 8676 12525 8732
rect 12525 8676 12529 8732
rect 12465 8672 12529 8676
rect 19740 8732 19804 8736
rect 19740 8676 19744 8732
rect 19744 8676 19800 8732
rect 19800 8676 19804 8732
rect 19740 8672 19804 8676
rect 19820 8732 19884 8736
rect 19820 8676 19824 8732
rect 19824 8676 19880 8732
rect 19880 8676 19884 8732
rect 19820 8672 19884 8676
rect 19900 8732 19964 8736
rect 19900 8676 19904 8732
rect 19904 8676 19960 8732
rect 19960 8676 19964 8732
rect 19900 8672 19964 8676
rect 19980 8732 20044 8736
rect 19980 8676 19984 8732
rect 19984 8676 20040 8732
rect 20040 8676 20044 8732
rect 19980 8672 20044 8676
rect 8467 8188 8531 8192
rect 8467 8132 8471 8188
rect 8471 8132 8527 8188
rect 8527 8132 8531 8188
rect 8467 8128 8531 8132
rect 8547 8188 8611 8192
rect 8547 8132 8551 8188
rect 8551 8132 8607 8188
rect 8607 8132 8611 8188
rect 8547 8128 8611 8132
rect 8627 8188 8691 8192
rect 8627 8132 8631 8188
rect 8631 8132 8687 8188
rect 8687 8132 8691 8188
rect 8627 8128 8691 8132
rect 8707 8188 8771 8192
rect 8707 8132 8711 8188
rect 8711 8132 8767 8188
rect 8767 8132 8771 8188
rect 8707 8128 8771 8132
rect 15982 8188 16046 8192
rect 15982 8132 15986 8188
rect 15986 8132 16042 8188
rect 16042 8132 16046 8188
rect 15982 8128 16046 8132
rect 16062 8188 16126 8192
rect 16062 8132 16066 8188
rect 16066 8132 16122 8188
rect 16122 8132 16126 8188
rect 16062 8128 16126 8132
rect 16142 8188 16206 8192
rect 16142 8132 16146 8188
rect 16146 8132 16202 8188
rect 16202 8132 16206 8188
rect 16142 8128 16206 8132
rect 16222 8188 16286 8192
rect 16222 8132 16226 8188
rect 16226 8132 16282 8188
rect 16282 8132 16286 8188
rect 16222 8128 16286 8132
rect 4709 7644 4773 7648
rect 4709 7588 4713 7644
rect 4713 7588 4769 7644
rect 4769 7588 4773 7644
rect 4709 7584 4773 7588
rect 4789 7644 4853 7648
rect 4789 7588 4793 7644
rect 4793 7588 4849 7644
rect 4849 7588 4853 7644
rect 4789 7584 4853 7588
rect 4869 7644 4933 7648
rect 4869 7588 4873 7644
rect 4873 7588 4929 7644
rect 4929 7588 4933 7644
rect 4869 7584 4933 7588
rect 4949 7644 5013 7648
rect 4949 7588 4953 7644
rect 4953 7588 5009 7644
rect 5009 7588 5013 7644
rect 4949 7584 5013 7588
rect 12225 7644 12289 7648
rect 12225 7588 12229 7644
rect 12229 7588 12285 7644
rect 12285 7588 12289 7644
rect 12225 7584 12289 7588
rect 12305 7644 12369 7648
rect 12305 7588 12309 7644
rect 12309 7588 12365 7644
rect 12365 7588 12369 7644
rect 12305 7584 12369 7588
rect 12385 7644 12449 7648
rect 12385 7588 12389 7644
rect 12389 7588 12445 7644
rect 12445 7588 12449 7644
rect 12385 7584 12449 7588
rect 12465 7644 12529 7648
rect 12465 7588 12469 7644
rect 12469 7588 12525 7644
rect 12525 7588 12529 7644
rect 12465 7584 12529 7588
rect 19740 7644 19804 7648
rect 19740 7588 19744 7644
rect 19744 7588 19800 7644
rect 19800 7588 19804 7644
rect 19740 7584 19804 7588
rect 19820 7644 19884 7648
rect 19820 7588 19824 7644
rect 19824 7588 19880 7644
rect 19880 7588 19884 7644
rect 19820 7584 19884 7588
rect 19900 7644 19964 7648
rect 19900 7588 19904 7644
rect 19904 7588 19960 7644
rect 19960 7588 19964 7644
rect 19900 7584 19964 7588
rect 19980 7644 20044 7648
rect 19980 7588 19984 7644
rect 19984 7588 20040 7644
rect 20040 7588 20044 7644
rect 19980 7584 20044 7588
rect 8467 7100 8531 7104
rect 8467 7044 8471 7100
rect 8471 7044 8527 7100
rect 8527 7044 8531 7100
rect 8467 7040 8531 7044
rect 8547 7100 8611 7104
rect 8547 7044 8551 7100
rect 8551 7044 8607 7100
rect 8607 7044 8611 7100
rect 8547 7040 8611 7044
rect 8627 7100 8691 7104
rect 8627 7044 8631 7100
rect 8631 7044 8687 7100
rect 8687 7044 8691 7100
rect 8627 7040 8691 7044
rect 8707 7100 8771 7104
rect 8707 7044 8711 7100
rect 8711 7044 8767 7100
rect 8767 7044 8771 7100
rect 8707 7040 8771 7044
rect 15982 7100 16046 7104
rect 15982 7044 15986 7100
rect 15986 7044 16042 7100
rect 16042 7044 16046 7100
rect 15982 7040 16046 7044
rect 16062 7100 16126 7104
rect 16062 7044 16066 7100
rect 16066 7044 16122 7100
rect 16122 7044 16126 7100
rect 16062 7040 16126 7044
rect 16142 7100 16206 7104
rect 16142 7044 16146 7100
rect 16146 7044 16202 7100
rect 16202 7044 16206 7100
rect 16142 7040 16206 7044
rect 16222 7100 16286 7104
rect 16222 7044 16226 7100
rect 16226 7044 16282 7100
rect 16282 7044 16286 7100
rect 16222 7040 16286 7044
rect 22140 6836 22204 6900
rect 22140 6666 22204 6730
rect 4709 6556 4773 6560
rect 4709 6500 4713 6556
rect 4713 6500 4769 6556
rect 4769 6500 4773 6556
rect 4709 6496 4773 6500
rect 4789 6556 4853 6560
rect 4789 6500 4793 6556
rect 4793 6500 4849 6556
rect 4849 6500 4853 6556
rect 4789 6496 4853 6500
rect 4869 6556 4933 6560
rect 4869 6500 4873 6556
rect 4873 6500 4929 6556
rect 4929 6500 4933 6556
rect 4869 6496 4933 6500
rect 4949 6556 5013 6560
rect 4949 6500 4953 6556
rect 4953 6500 5009 6556
rect 5009 6500 5013 6556
rect 4949 6496 5013 6500
rect 12225 6556 12289 6560
rect 12225 6500 12229 6556
rect 12229 6500 12285 6556
rect 12285 6500 12289 6556
rect 12225 6496 12289 6500
rect 12305 6556 12369 6560
rect 12305 6500 12309 6556
rect 12309 6500 12365 6556
rect 12365 6500 12369 6556
rect 12305 6496 12369 6500
rect 12385 6556 12449 6560
rect 12385 6500 12389 6556
rect 12389 6500 12445 6556
rect 12445 6500 12449 6556
rect 12385 6496 12449 6500
rect 12465 6556 12529 6560
rect 12465 6500 12469 6556
rect 12469 6500 12525 6556
rect 12525 6500 12529 6556
rect 12465 6496 12529 6500
rect 19740 6556 19804 6560
rect 19740 6500 19744 6556
rect 19744 6500 19800 6556
rect 19800 6500 19804 6556
rect 19740 6496 19804 6500
rect 19820 6556 19884 6560
rect 19820 6500 19824 6556
rect 19824 6500 19880 6556
rect 19880 6500 19884 6556
rect 19820 6496 19884 6500
rect 19900 6556 19964 6560
rect 19900 6500 19904 6556
rect 19904 6500 19960 6556
rect 19960 6500 19964 6556
rect 19900 6496 19964 6500
rect 19980 6556 20044 6560
rect 19980 6500 19984 6556
rect 19984 6500 20040 6556
rect 20040 6500 20044 6556
rect 19980 6496 20044 6500
rect 8467 6012 8531 6016
rect 8467 5956 8471 6012
rect 8471 5956 8527 6012
rect 8527 5956 8531 6012
rect 8467 5952 8531 5956
rect 8547 6012 8611 6016
rect 8547 5956 8551 6012
rect 8551 5956 8607 6012
rect 8607 5956 8611 6012
rect 8547 5952 8611 5956
rect 8627 6012 8691 6016
rect 8627 5956 8631 6012
rect 8631 5956 8687 6012
rect 8687 5956 8691 6012
rect 8627 5952 8691 5956
rect 8707 6012 8771 6016
rect 8707 5956 8711 6012
rect 8711 5956 8767 6012
rect 8767 5956 8771 6012
rect 8707 5952 8771 5956
rect 15982 6012 16046 6016
rect 15982 5956 15986 6012
rect 15986 5956 16042 6012
rect 16042 5956 16046 6012
rect 15982 5952 16046 5956
rect 16062 6012 16126 6016
rect 16062 5956 16066 6012
rect 16066 5956 16122 6012
rect 16122 5956 16126 6012
rect 16062 5952 16126 5956
rect 16142 6012 16206 6016
rect 16142 5956 16146 6012
rect 16146 5956 16202 6012
rect 16202 5956 16206 6012
rect 16142 5952 16206 5956
rect 16222 6012 16286 6016
rect 16222 5956 16226 6012
rect 16226 5956 16282 6012
rect 16282 5956 16286 6012
rect 16222 5952 16286 5956
rect 4709 5468 4773 5472
rect 4709 5412 4713 5468
rect 4713 5412 4769 5468
rect 4769 5412 4773 5468
rect 4709 5408 4773 5412
rect 4789 5468 4853 5472
rect 4789 5412 4793 5468
rect 4793 5412 4849 5468
rect 4849 5412 4853 5468
rect 4789 5408 4853 5412
rect 4869 5468 4933 5472
rect 4869 5412 4873 5468
rect 4873 5412 4929 5468
rect 4929 5412 4933 5468
rect 4869 5408 4933 5412
rect 4949 5468 5013 5472
rect 4949 5412 4953 5468
rect 4953 5412 5009 5468
rect 5009 5412 5013 5468
rect 4949 5408 5013 5412
rect 12225 5468 12289 5472
rect 12225 5412 12229 5468
rect 12229 5412 12285 5468
rect 12285 5412 12289 5468
rect 12225 5408 12289 5412
rect 12305 5468 12369 5472
rect 12305 5412 12309 5468
rect 12309 5412 12365 5468
rect 12365 5412 12369 5468
rect 12305 5408 12369 5412
rect 12385 5468 12449 5472
rect 12385 5412 12389 5468
rect 12389 5412 12445 5468
rect 12445 5412 12449 5468
rect 12385 5408 12449 5412
rect 12465 5468 12529 5472
rect 12465 5412 12469 5468
rect 12469 5412 12525 5468
rect 12525 5412 12529 5468
rect 12465 5408 12529 5412
rect 19740 5468 19804 5472
rect 19740 5412 19744 5468
rect 19744 5412 19800 5468
rect 19800 5412 19804 5468
rect 19740 5408 19804 5412
rect 19820 5468 19884 5472
rect 19820 5412 19824 5468
rect 19824 5412 19880 5468
rect 19880 5412 19884 5468
rect 19820 5408 19884 5412
rect 19900 5468 19964 5472
rect 19900 5412 19904 5468
rect 19904 5412 19960 5468
rect 19960 5412 19964 5468
rect 19900 5408 19964 5412
rect 19980 5468 20044 5472
rect 19980 5412 19984 5468
rect 19984 5412 20040 5468
rect 20040 5412 20044 5468
rect 19980 5408 20044 5412
rect 8467 4924 8531 4928
rect 8467 4868 8471 4924
rect 8471 4868 8527 4924
rect 8527 4868 8531 4924
rect 8467 4864 8531 4868
rect 8547 4924 8611 4928
rect 8547 4868 8551 4924
rect 8551 4868 8607 4924
rect 8607 4868 8611 4924
rect 8547 4864 8611 4868
rect 8627 4924 8691 4928
rect 8627 4868 8631 4924
rect 8631 4868 8687 4924
rect 8687 4868 8691 4924
rect 8627 4864 8691 4868
rect 8707 4924 8771 4928
rect 8707 4868 8711 4924
rect 8711 4868 8767 4924
rect 8767 4868 8771 4924
rect 8707 4864 8771 4868
rect 15982 4924 16046 4928
rect 15982 4868 15986 4924
rect 15986 4868 16042 4924
rect 16042 4868 16046 4924
rect 15982 4864 16046 4868
rect 16062 4924 16126 4928
rect 16062 4868 16066 4924
rect 16066 4868 16122 4924
rect 16122 4868 16126 4924
rect 16062 4864 16126 4868
rect 16142 4924 16206 4928
rect 16142 4868 16146 4924
rect 16146 4868 16202 4924
rect 16202 4868 16206 4924
rect 16142 4864 16206 4868
rect 16222 4924 16286 4928
rect 16222 4868 16226 4924
rect 16226 4868 16282 4924
rect 16282 4868 16286 4924
rect 16222 4864 16286 4868
rect 4709 4380 4773 4384
rect 4709 4324 4713 4380
rect 4713 4324 4769 4380
rect 4769 4324 4773 4380
rect 4709 4320 4773 4324
rect 4789 4380 4853 4384
rect 4789 4324 4793 4380
rect 4793 4324 4849 4380
rect 4849 4324 4853 4380
rect 4789 4320 4853 4324
rect 4869 4380 4933 4384
rect 4869 4324 4873 4380
rect 4873 4324 4929 4380
rect 4929 4324 4933 4380
rect 4869 4320 4933 4324
rect 4949 4380 5013 4384
rect 4949 4324 4953 4380
rect 4953 4324 5009 4380
rect 5009 4324 5013 4380
rect 4949 4320 5013 4324
rect 12225 4380 12289 4384
rect 12225 4324 12229 4380
rect 12229 4324 12285 4380
rect 12285 4324 12289 4380
rect 12225 4320 12289 4324
rect 12305 4380 12369 4384
rect 12305 4324 12309 4380
rect 12309 4324 12365 4380
rect 12365 4324 12369 4380
rect 12305 4320 12369 4324
rect 12385 4380 12449 4384
rect 12385 4324 12389 4380
rect 12389 4324 12445 4380
rect 12445 4324 12449 4380
rect 12385 4320 12449 4324
rect 12465 4380 12529 4384
rect 12465 4324 12469 4380
rect 12469 4324 12525 4380
rect 12525 4324 12529 4380
rect 12465 4320 12529 4324
rect 19740 4380 19804 4384
rect 19740 4324 19744 4380
rect 19744 4324 19800 4380
rect 19800 4324 19804 4380
rect 19740 4320 19804 4324
rect 19820 4380 19884 4384
rect 19820 4324 19824 4380
rect 19824 4324 19880 4380
rect 19880 4324 19884 4380
rect 19820 4320 19884 4324
rect 19900 4380 19964 4384
rect 19900 4324 19904 4380
rect 19904 4324 19960 4380
rect 19960 4324 19964 4380
rect 19900 4320 19964 4324
rect 19980 4380 20044 4384
rect 19980 4324 19984 4380
rect 19984 4324 20040 4380
rect 20040 4324 20044 4380
rect 19980 4320 20044 4324
rect 8467 3836 8531 3840
rect 8467 3780 8471 3836
rect 8471 3780 8527 3836
rect 8527 3780 8531 3836
rect 8467 3776 8531 3780
rect 8547 3836 8611 3840
rect 8547 3780 8551 3836
rect 8551 3780 8607 3836
rect 8607 3780 8611 3836
rect 8547 3776 8611 3780
rect 8627 3836 8691 3840
rect 8627 3780 8631 3836
rect 8631 3780 8687 3836
rect 8687 3780 8691 3836
rect 8627 3776 8691 3780
rect 8707 3836 8771 3840
rect 8707 3780 8711 3836
rect 8711 3780 8767 3836
rect 8767 3780 8771 3836
rect 8707 3776 8771 3780
rect 15982 3836 16046 3840
rect 15982 3780 15986 3836
rect 15986 3780 16042 3836
rect 16042 3780 16046 3836
rect 15982 3776 16046 3780
rect 16062 3836 16126 3840
rect 16062 3780 16066 3836
rect 16066 3780 16122 3836
rect 16122 3780 16126 3836
rect 16062 3776 16126 3780
rect 16142 3836 16206 3840
rect 16142 3780 16146 3836
rect 16146 3780 16202 3836
rect 16202 3780 16206 3836
rect 16142 3776 16206 3780
rect 16222 3836 16286 3840
rect 16222 3780 16226 3836
rect 16226 3780 16282 3836
rect 16282 3780 16286 3836
rect 16222 3776 16286 3780
rect 4709 3292 4773 3296
rect 4709 3236 4713 3292
rect 4713 3236 4769 3292
rect 4769 3236 4773 3292
rect 4709 3232 4773 3236
rect 4789 3292 4853 3296
rect 4789 3236 4793 3292
rect 4793 3236 4849 3292
rect 4849 3236 4853 3292
rect 4789 3232 4853 3236
rect 4869 3292 4933 3296
rect 4869 3236 4873 3292
rect 4873 3236 4929 3292
rect 4929 3236 4933 3292
rect 4869 3232 4933 3236
rect 4949 3292 5013 3296
rect 4949 3236 4953 3292
rect 4953 3236 5009 3292
rect 5009 3236 5013 3292
rect 4949 3232 5013 3236
rect 12225 3292 12289 3296
rect 12225 3236 12229 3292
rect 12229 3236 12285 3292
rect 12285 3236 12289 3292
rect 12225 3232 12289 3236
rect 12305 3292 12369 3296
rect 12305 3236 12309 3292
rect 12309 3236 12365 3292
rect 12365 3236 12369 3292
rect 12305 3232 12369 3236
rect 12385 3292 12449 3296
rect 12385 3236 12389 3292
rect 12389 3236 12445 3292
rect 12445 3236 12449 3292
rect 12385 3232 12449 3236
rect 12465 3292 12529 3296
rect 12465 3236 12469 3292
rect 12469 3236 12525 3292
rect 12525 3236 12529 3292
rect 12465 3232 12529 3236
rect 19740 3292 19804 3296
rect 19740 3236 19744 3292
rect 19744 3236 19800 3292
rect 19800 3236 19804 3292
rect 19740 3232 19804 3236
rect 19820 3292 19884 3296
rect 19820 3236 19824 3292
rect 19824 3236 19880 3292
rect 19880 3236 19884 3292
rect 19820 3232 19884 3236
rect 19900 3292 19964 3296
rect 19900 3236 19904 3292
rect 19904 3236 19960 3292
rect 19960 3236 19964 3292
rect 19900 3232 19964 3236
rect 19980 3292 20044 3296
rect 19980 3236 19984 3292
rect 19984 3236 20040 3292
rect 20040 3236 20044 3292
rect 19980 3232 20044 3236
rect 8467 2748 8531 2752
rect 8467 2692 8471 2748
rect 8471 2692 8527 2748
rect 8527 2692 8531 2748
rect 8467 2688 8531 2692
rect 8547 2748 8611 2752
rect 8547 2692 8551 2748
rect 8551 2692 8607 2748
rect 8607 2692 8611 2748
rect 8547 2688 8611 2692
rect 8627 2748 8691 2752
rect 8627 2692 8631 2748
rect 8631 2692 8687 2748
rect 8687 2692 8691 2748
rect 8627 2688 8691 2692
rect 8707 2748 8771 2752
rect 8707 2692 8711 2748
rect 8711 2692 8767 2748
rect 8767 2692 8771 2748
rect 8707 2688 8771 2692
rect 15982 2748 16046 2752
rect 15982 2692 15986 2748
rect 15986 2692 16042 2748
rect 16042 2692 16046 2748
rect 15982 2688 16046 2692
rect 16062 2748 16126 2752
rect 16062 2692 16066 2748
rect 16066 2692 16122 2748
rect 16122 2692 16126 2748
rect 16062 2688 16126 2692
rect 16142 2748 16206 2752
rect 16142 2692 16146 2748
rect 16146 2692 16202 2748
rect 16202 2692 16206 2748
rect 16142 2688 16206 2692
rect 16222 2748 16286 2752
rect 16222 2692 16226 2748
rect 16226 2692 16282 2748
rect 16282 2692 16286 2748
rect 16222 2688 16286 2692
rect 4709 2204 4773 2208
rect 4709 2148 4713 2204
rect 4713 2148 4769 2204
rect 4769 2148 4773 2204
rect 4709 2144 4773 2148
rect 4789 2204 4853 2208
rect 4789 2148 4793 2204
rect 4793 2148 4849 2204
rect 4849 2148 4853 2204
rect 4789 2144 4853 2148
rect 4869 2204 4933 2208
rect 4869 2148 4873 2204
rect 4873 2148 4929 2204
rect 4929 2148 4933 2204
rect 4869 2144 4933 2148
rect 4949 2204 5013 2208
rect 4949 2148 4953 2204
rect 4953 2148 5009 2204
rect 5009 2148 5013 2204
rect 4949 2144 5013 2148
rect 12225 2204 12289 2208
rect 12225 2148 12229 2204
rect 12229 2148 12285 2204
rect 12285 2148 12289 2204
rect 12225 2144 12289 2148
rect 12305 2204 12369 2208
rect 12305 2148 12309 2204
rect 12309 2148 12365 2204
rect 12365 2148 12369 2204
rect 12305 2144 12369 2148
rect 12385 2204 12449 2208
rect 12385 2148 12389 2204
rect 12389 2148 12445 2204
rect 12445 2148 12449 2204
rect 12385 2144 12449 2148
rect 12465 2204 12529 2208
rect 12465 2148 12469 2204
rect 12469 2148 12525 2204
rect 12525 2148 12529 2204
rect 12465 2144 12529 2148
rect 19740 2204 19804 2208
rect 19740 2148 19744 2204
rect 19744 2148 19800 2204
rect 19800 2148 19804 2204
rect 19740 2144 19804 2148
rect 19820 2204 19884 2208
rect 19820 2148 19824 2204
rect 19824 2148 19880 2204
rect 19880 2148 19884 2204
rect 19820 2144 19884 2148
rect 19900 2204 19964 2208
rect 19900 2148 19904 2204
rect 19904 2148 19960 2204
rect 19960 2148 19964 2204
rect 19900 2144 19964 2148
rect 19980 2204 20044 2208
rect 19980 2148 19984 2204
rect 19984 2148 20040 2204
rect 20040 2148 20044 2204
rect 19980 2144 20044 2148
<< metal4 >>
rect 4701 21792 5022 22352
rect 4701 21728 4709 21792
rect 4773 21728 4789 21792
rect 4853 21728 4869 21792
rect 4933 21728 4949 21792
rect 5013 21728 5022 21792
rect 4701 20704 5022 21728
rect 4701 20640 4709 20704
rect 4773 20640 4789 20704
rect 4853 20640 4869 20704
rect 4933 20640 4949 20704
rect 5013 20640 5022 20704
rect 4701 19616 5022 20640
rect 4701 19552 4709 19616
rect 4773 19552 4789 19616
rect 4853 19552 4869 19616
rect 4933 19552 4949 19616
rect 5013 19552 5022 19616
rect 4701 18528 5022 19552
rect 4701 18464 4709 18528
rect 4773 18464 4789 18528
rect 4853 18464 4869 18528
rect 4933 18464 4949 18528
rect 5013 18464 5022 18528
rect 4701 17440 5022 18464
rect 4701 17376 4709 17440
rect 4773 17376 4789 17440
rect 4853 17376 4869 17440
rect 4933 17376 4949 17440
rect 5013 17376 5022 17440
rect 4701 16352 5022 17376
rect 4701 16288 4709 16352
rect 4773 16288 4789 16352
rect 4853 16288 4869 16352
rect 4933 16288 4949 16352
rect 5013 16288 5022 16352
rect 4701 15264 5022 16288
rect 4701 15200 4709 15264
rect 4773 15200 4789 15264
rect 4853 15200 4869 15264
rect 4933 15200 4949 15264
rect 5013 15200 5022 15264
rect 59 14924 125 14925
rect 59 14860 60 14924
rect 124 14860 125 14924
rect 59 14859 125 14860
rect 62 14517 122 14859
rect 59 14516 125 14517
rect 59 14452 60 14516
rect 124 14452 125 14516
rect 59 14451 125 14452
rect 4701 14176 5022 15200
rect 4701 14112 4709 14176
rect 4773 14112 4789 14176
rect 4853 14112 4869 14176
rect 4933 14112 4949 14176
rect 5013 14112 5022 14176
rect 4701 13088 5022 14112
rect 4701 13024 4709 13088
rect 4773 13024 4789 13088
rect 4853 13024 4869 13088
rect 4933 13024 4949 13088
rect 5013 13024 5022 13088
rect 4701 12000 5022 13024
rect 4701 11936 4709 12000
rect 4773 11936 4789 12000
rect 4853 11936 4869 12000
rect 4933 11936 4949 12000
rect 5013 11936 5022 12000
rect 4701 10912 5022 11936
rect 4701 10848 4709 10912
rect 4773 10848 4789 10912
rect 4853 10848 4869 10912
rect 4933 10848 4949 10912
rect 5013 10848 5022 10912
rect 4701 9824 5022 10848
rect 4701 9760 4709 9824
rect 4773 9760 4789 9824
rect 4853 9760 4869 9824
rect 4933 9760 4949 9824
rect 5013 9760 5022 9824
rect 4701 8736 5022 9760
rect 4701 8672 4709 8736
rect 4773 8672 4789 8736
rect 4853 8672 4869 8736
rect 4933 8672 4949 8736
rect 5013 8672 5022 8736
rect 4701 7648 5022 8672
rect 4701 7584 4709 7648
rect 4773 7584 4789 7648
rect 4853 7584 4869 7648
rect 4933 7584 4949 7648
rect 5013 7584 5022 7648
rect 4701 6560 5022 7584
rect 4701 6496 4709 6560
rect 4773 6496 4789 6560
rect 4853 6496 4869 6560
rect 4933 6496 4949 6560
rect 5013 6496 5022 6560
rect 4701 5472 5022 6496
rect 4701 5408 4709 5472
rect 4773 5408 4789 5472
rect 4853 5408 4869 5472
rect 4933 5408 4949 5472
rect 5013 5408 5022 5472
rect 4701 4384 5022 5408
rect 4701 4320 4709 4384
rect 4773 4320 4789 4384
rect 4853 4320 4869 4384
rect 4933 4320 4949 4384
rect 5013 4320 5022 4384
rect 4701 3296 5022 4320
rect 4701 3232 4709 3296
rect 4773 3232 4789 3296
rect 4853 3232 4869 3296
rect 4933 3232 4949 3296
rect 5013 3232 5022 3296
rect 4701 2208 5022 3232
rect 4701 2144 4709 2208
rect 4773 2144 4789 2208
rect 4853 2144 4869 2208
rect 4933 2144 4949 2208
rect 5013 2144 5022 2208
rect 4701 2128 5022 2144
rect 8459 22336 8779 22352
rect 8459 22272 8467 22336
rect 8531 22272 8547 22336
rect 8611 22272 8627 22336
rect 8691 22272 8707 22336
rect 8771 22272 8779 22336
rect 8459 21248 8779 22272
rect 8459 21184 8467 21248
rect 8531 21184 8547 21248
rect 8611 21184 8627 21248
rect 8691 21184 8707 21248
rect 8771 21184 8779 21248
rect 8459 20160 8779 21184
rect 8459 20096 8467 20160
rect 8531 20096 8547 20160
rect 8611 20096 8627 20160
rect 8691 20096 8707 20160
rect 8771 20096 8779 20160
rect 8459 19072 8779 20096
rect 8459 19008 8467 19072
rect 8531 19008 8547 19072
rect 8611 19008 8627 19072
rect 8691 19008 8707 19072
rect 8771 19008 8779 19072
rect 8459 17984 8779 19008
rect 8459 17920 8467 17984
rect 8531 17920 8547 17984
rect 8611 17920 8627 17984
rect 8691 17920 8707 17984
rect 8771 17920 8779 17984
rect 8459 16896 8779 17920
rect 8459 16832 8467 16896
rect 8531 16832 8547 16896
rect 8611 16832 8627 16896
rect 8691 16832 8707 16896
rect 8771 16832 8779 16896
rect 8459 15808 8779 16832
rect 8459 15744 8467 15808
rect 8531 15744 8547 15808
rect 8611 15744 8627 15808
rect 8691 15744 8707 15808
rect 8771 15744 8779 15808
rect 8459 14720 8779 15744
rect 8459 14656 8467 14720
rect 8531 14656 8547 14720
rect 8611 14656 8627 14720
rect 8691 14656 8707 14720
rect 8771 14656 8779 14720
rect 8459 13632 8779 14656
rect 8459 13568 8467 13632
rect 8531 13568 8547 13632
rect 8611 13568 8627 13632
rect 8691 13568 8707 13632
rect 8771 13568 8779 13632
rect 8459 12544 8779 13568
rect 8459 12480 8467 12544
rect 8531 12480 8547 12544
rect 8611 12480 8627 12544
rect 8691 12480 8707 12544
rect 8771 12480 8779 12544
rect 8459 11456 8779 12480
rect 8459 11392 8467 11456
rect 8531 11392 8547 11456
rect 8611 11392 8627 11456
rect 8691 11392 8707 11456
rect 8771 11392 8779 11456
rect 8459 10368 8779 11392
rect 8459 10304 8467 10368
rect 8531 10304 8547 10368
rect 8611 10304 8627 10368
rect 8691 10304 8707 10368
rect 8771 10304 8779 10368
rect 8459 9280 8779 10304
rect 8459 9216 8467 9280
rect 8531 9216 8547 9280
rect 8611 9216 8627 9280
rect 8691 9216 8707 9280
rect 8771 9216 8779 9280
rect 8459 8192 8779 9216
rect 8459 8128 8467 8192
rect 8531 8128 8547 8192
rect 8611 8128 8627 8192
rect 8691 8128 8707 8192
rect 8771 8128 8779 8192
rect 8459 7104 8779 8128
rect 8459 7040 8467 7104
rect 8531 7040 8547 7104
rect 8611 7040 8627 7104
rect 8691 7040 8707 7104
rect 8771 7040 8779 7104
rect 8459 6016 8779 7040
rect 8459 5952 8467 6016
rect 8531 5952 8547 6016
rect 8611 5952 8627 6016
rect 8691 5952 8707 6016
rect 8771 5952 8779 6016
rect 8459 4928 8779 5952
rect 8459 4864 8467 4928
rect 8531 4864 8547 4928
rect 8611 4864 8627 4928
rect 8691 4864 8707 4928
rect 8771 4864 8779 4928
rect 8459 3840 8779 4864
rect 8459 3776 8467 3840
rect 8531 3776 8547 3840
rect 8611 3776 8627 3840
rect 8691 3776 8707 3840
rect 8771 3776 8779 3840
rect 8459 2752 8779 3776
rect 8459 2688 8467 2752
rect 8531 2688 8547 2752
rect 8611 2688 8627 2752
rect 8691 2688 8707 2752
rect 8771 2688 8779 2752
rect 8459 2128 8779 2688
rect 12217 21792 12537 22352
rect 12217 21728 12225 21792
rect 12289 21728 12305 21792
rect 12369 21728 12385 21792
rect 12449 21728 12465 21792
rect 12529 21728 12537 21792
rect 12217 20704 12537 21728
rect 12217 20640 12225 20704
rect 12289 20640 12305 20704
rect 12369 20640 12385 20704
rect 12449 20640 12465 20704
rect 12529 20640 12537 20704
rect 12217 19616 12537 20640
rect 12217 19552 12225 19616
rect 12289 19552 12305 19616
rect 12369 19552 12385 19616
rect 12449 19552 12465 19616
rect 12529 19552 12537 19616
rect 12217 18528 12537 19552
rect 12217 18464 12225 18528
rect 12289 18464 12305 18528
rect 12369 18464 12385 18528
rect 12449 18464 12465 18528
rect 12529 18464 12537 18528
rect 12217 17440 12537 18464
rect 12217 17376 12225 17440
rect 12289 17376 12305 17440
rect 12369 17376 12385 17440
rect 12449 17376 12465 17440
rect 12529 17376 12537 17440
rect 12217 16352 12537 17376
rect 12217 16288 12225 16352
rect 12289 16288 12305 16352
rect 12369 16288 12385 16352
rect 12449 16288 12465 16352
rect 12529 16288 12537 16352
rect 12217 15264 12537 16288
rect 12217 15200 12225 15264
rect 12289 15200 12305 15264
rect 12369 15200 12385 15264
rect 12449 15200 12465 15264
rect 12529 15200 12537 15264
rect 12217 14176 12537 15200
rect 12217 14112 12225 14176
rect 12289 14112 12305 14176
rect 12369 14112 12385 14176
rect 12449 14112 12465 14176
rect 12529 14112 12537 14176
rect 12217 13088 12537 14112
rect 12217 13024 12225 13088
rect 12289 13024 12305 13088
rect 12369 13024 12385 13088
rect 12449 13024 12465 13088
rect 12529 13024 12537 13088
rect 12217 12000 12537 13024
rect 12217 11936 12225 12000
rect 12289 11936 12305 12000
rect 12369 11936 12385 12000
rect 12449 11936 12465 12000
rect 12529 11936 12537 12000
rect 12217 10912 12537 11936
rect 12217 10848 12225 10912
rect 12289 10848 12305 10912
rect 12369 10848 12385 10912
rect 12449 10848 12465 10912
rect 12529 10848 12537 10912
rect 12217 9824 12537 10848
rect 12217 9760 12225 9824
rect 12289 9760 12305 9824
rect 12369 9760 12385 9824
rect 12449 9760 12465 9824
rect 12529 9760 12537 9824
rect 12217 8736 12537 9760
rect 12217 8672 12225 8736
rect 12289 8672 12305 8736
rect 12369 8672 12385 8736
rect 12449 8672 12465 8736
rect 12529 8672 12537 8736
rect 12217 7648 12537 8672
rect 12217 7584 12225 7648
rect 12289 7584 12305 7648
rect 12369 7584 12385 7648
rect 12449 7584 12465 7648
rect 12529 7584 12537 7648
rect 12217 6560 12537 7584
rect 12217 6496 12225 6560
rect 12289 6496 12305 6560
rect 12369 6496 12385 6560
rect 12449 6496 12465 6560
rect 12529 6496 12537 6560
rect 12217 5472 12537 6496
rect 12217 5408 12225 5472
rect 12289 5408 12305 5472
rect 12369 5408 12385 5472
rect 12449 5408 12465 5472
rect 12529 5408 12537 5472
rect 12217 4384 12537 5408
rect 12217 4320 12225 4384
rect 12289 4320 12305 4384
rect 12369 4320 12385 4384
rect 12449 4320 12465 4384
rect 12529 4320 12537 4384
rect 12217 3296 12537 4320
rect 12217 3232 12225 3296
rect 12289 3232 12305 3296
rect 12369 3232 12385 3296
rect 12449 3232 12465 3296
rect 12529 3232 12537 3296
rect 12217 2208 12537 3232
rect 12217 2144 12225 2208
rect 12289 2144 12305 2208
rect 12369 2144 12385 2208
rect 12449 2144 12465 2208
rect 12529 2144 12537 2208
rect 12217 2128 12537 2144
rect 15974 22336 16294 22352
rect 15974 22272 15982 22336
rect 16046 22272 16062 22336
rect 16126 22272 16142 22336
rect 16206 22272 16222 22336
rect 16286 22272 16294 22336
rect 15974 21248 16294 22272
rect 15974 21184 15982 21248
rect 16046 21184 16062 21248
rect 16126 21184 16142 21248
rect 16206 21184 16222 21248
rect 16286 21184 16294 21248
rect 15974 20160 16294 21184
rect 15974 20096 15982 20160
rect 16046 20096 16062 20160
rect 16126 20096 16142 20160
rect 16206 20096 16222 20160
rect 16286 20096 16294 20160
rect 15974 19072 16294 20096
rect 15974 19008 15982 19072
rect 16046 19008 16062 19072
rect 16126 19008 16142 19072
rect 16206 19008 16222 19072
rect 16286 19008 16294 19072
rect 15974 17984 16294 19008
rect 15974 17920 15982 17984
rect 16046 17920 16062 17984
rect 16126 17920 16142 17984
rect 16206 17920 16222 17984
rect 16286 17920 16294 17984
rect 15974 16896 16294 17920
rect 15974 16832 15982 16896
rect 16046 16832 16062 16896
rect 16126 16832 16142 16896
rect 16206 16832 16222 16896
rect 16286 16832 16294 16896
rect 15974 15808 16294 16832
rect 15974 15744 15982 15808
rect 16046 15744 16062 15808
rect 16126 15744 16142 15808
rect 16206 15744 16222 15808
rect 16286 15744 16294 15808
rect 15974 14720 16294 15744
rect 15974 14656 15982 14720
rect 16046 14656 16062 14720
rect 16126 14656 16142 14720
rect 16206 14656 16222 14720
rect 16286 14656 16294 14720
rect 15974 13632 16294 14656
rect 15974 13568 15982 13632
rect 16046 13568 16062 13632
rect 16126 13568 16142 13632
rect 16206 13568 16222 13632
rect 16286 13568 16294 13632
rect 15974 12544 16294 13568
rect 15974 12480 15982 12544
rect 16046 12480 16062 12544
rect 16126 12480 16142 12544
rect 16206 12480 16222 12544
rect 16286 12480 16294 12544
rect 15974 11456 16294 12480
rect 15974 11392 15982 11456
rect 16046 11392 16062 11456
rect 16126 11392 16142 11456
rect 16206 11392 16222 11456
rect 16286 11392 16294 11456
rect 15974 10368 16294 11392
rect 15974 10304 15982 10368
rect 16046 10304 16062 10368
rect 16126 10304 16142 10368
rect 16206 10304 16222 10368
rect 16286 10304 16294 10368
rect 15974 9280 16294 10304
rect 15974 9216 15982 9280
rect 16046 9216 16062 9280
rect 16126 9216 16142 9280
rect 16206 9216 16222 9280
rect 16286 9216 16294 9280
rect 15974 8192 16294 9216
rect 15974 8128 15982 8192
rect 16046 8128 16062 8192
rect 16126 8128 16142 8192
rect 16206 8128 16222 8192
rect 16286 8128 16294 8192
rect 15974 7104 16294 8128
rect 15974 7040 15982 7104
rect 16046 7040 16062 7104
rect 16126 7040 16142 7104
rect 16206 7040 16222 7104
rect 16286 7040 16294 7104
rect 15974 6016 16294 7040
rect 15974 5952 15982 6016
rect 16046 5952 16062 6016
rect 16126 5952 16142 6016
rect 16206 5952 16222 6016
rect 16286 5952 16294 6016
rect 15974 4928 16294 5952
rect 15974 4864 15982 4928
rect 16046 4864 16062 4928
rect 16126 4864 16142 4928
rect 16206 4864 16222 4928
rect 16286 4864 16294 4928
rect 15974 3840 16294 4864
rect 15974 3776 15982 3840
rect 16046 3776 16062 3840
rect 16126 3776 16142 3840
rect 16206 3776 16222 3840
rect 16286 3776 16294 3840
rect 15974 2752 16294 3776
rect 15974 2688 15982 2752
rect 16046 2688 16062 2752
rect 16126 2688 16142 2752
rect 16206 2688 16222 2752
rect 16286 2688 16294 2752
rect 15974 2128 16294 2688
rect 19732 21792 20052 22352
rect 19732 21728 19740 21792
rect 19804 21728 19820 21792
rect 19884 21728 19900 21792
rect 19964 21728 19980 21792
rect 20044 21728 20052 21792
rect 19732 20704 20052 21728
rect 19732 20640 19740 20704
rect 19804 20640 19820 20704
rect 19884 20640 19900 20704
rect 19964 20640 19980 20704
rect 20044 20640 20052 20704
rect 19732 19616 20052 20640
rect 19732 19552 19740 19616
rect 19804 19552 19820 19616
rect 19884 19552 19900 19616
rect 19964 19552 19980 19616
rect 20044 19552 20052 19616
rect 19732 18528 20052 19552
rect 19732 18464 19740 18528
rect 19804 18464 19820 18528
rect 19884 18464 19900 18528
rect 19964 18464 19980 18528
rect 20044 18464 20052 18528
rect 19732 17440 20052 18464
rect 19732 17376 19740 17440
rect 19804 17376 19820 17440
rect 19884 17376 19900 17440
rect 19964 17376 19980 17440
rect 20044 17376 20052 17440
rect 19732 16352 20052 17376
rect 19732 16288 19740 16352
rect 19804 16288 19820 16352
rect 19884 16288 19900 16352
rect 19964 16288 19980 16352
rect 20044 16288 20052 16352
rect 19732 15264 20052 16288
rect 19732 15200 19740 15264
rect 19804 15200 19820 15264
rect 19884 15200 19900 15264
rect 19964 15200 19980 15264
rect 20044 15200 20052 15264
rect 19732 14176 20052 15200
rect 22139 14652 22205 14653
rect 22139 14588 22140 14652
rect 22204 14588 22205 14652
rect 22139 14587 22205 14588
rect 22142 14381 22202 14587
rect 22139 14380 22205 14381
rect 22139 14316 22140 14380
rect 22204 14316 22205 14380
rect 22139 14315 22205 14316
rect 19732 14112 19740 14176
rect 19804 14112 19820 14176
rect 19884 14112 19900 14176
rect 19964 14112 19980 14176
rect 20044 14112 20052 14176
rect 19732 13088 20052 14112
rect 19732 13024 19740 13088
rect 19804 13024 19820 13088
rect 19884 13024 19900 13088
rect 19964 13024 19980 13088
rect 20044 13024 20052 13088
rect 19732 12000 20052 13024
rect 19732 11936 19740 12000
rect 19804 11936 19820 12000
rect 19884 11936 19900 12000
rect 19964 11936 19980 12000
rect 20044 11936 20052 12000
rect 19732 10912 20052 11936
rect 19732 10848 19740 10912
rect 19804 10848 19820 10912
rect 19884 10848 19900 10912
rect 19964 10848 19980 10912
rect 20044 10848 20052 10912
rect 19732 9824 20052 10848
rect 19732 9760 19740 9824
rect 19804 9760 19820 9824
rect 19884 9760 19900 9824
rect 19964 9760 19980 9824
rect 20044 9760 20052 9824
rect 19732 8736 20052 9760
rect 19732 8672 19740 8736
rect 19804 8672 19820 8736
rect 19884 8672 19900 8736
rect 19964 8672 19980 8736
rect 20044 8672 20052 8736
rect 19732 7648 20052 8672
rect 19732 7584 19740 7648
rect 19804 7584 19820 7648
rect 19884 7584 19900 7648
rect 19964 7584 19980 7648
rect 20044 7584 20052 7648
rect 19732 6560 20052 7584
rect 22139 6900 22205 6901
rect 22139 6836 22140 6900
rect 22204 6836 22205 6900
rect 22139 6835 22205 6836
rect 22142 6731 22202 6835
rect 22139 6730 22205 6731
rect 22139 6666 22140 6730
rect 22204 6666 22205 6730
rect 22139 6665 22205 6666
rect 19732 6496 19740 6560
rect 19804 6496 19820 6560
rect 19884 6496 19900 6560
rect 19964 6496 19980 6560
rect 20044 6496 20052 6560
rect 19732 5472 20052 6496
rect 19732 5408 19740 5472
rect 19804 5408 19820 5472
rect 19884 5408 19900 5472
rect 19964 5408 19980 5472
rect 20044 5408 20052 5472
rect 19732 4384 20052 5408
rect 19732 4320 19740 4384
rect 19804 4320 19820 4384
rect 19884 4320 19900 4384
rect 19964 4320 19980 4384
rect 20044 4320 20052 4384
rect 19732 3296 20052 4320
rect 19732 3232 19740 3296
rect 19804 3232 19820 3296
rect 19884 3232 19900 3296
rect 19964 3232 19980 3296
rect 20044 3232 20052 3296
rect 19732 2208 20052 3232
rect 19732 2144 19740 2208
rect 19804 2144 19820 2208
rect 19884 2144 19900 2208
rect 19964 2144 19980 2208
rect 20044 2144 20052 2208
rect 19732 2128 20052 2144
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_12 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_9 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_12
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_16
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_16 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_20
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_74 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_48
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_54 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_54
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_78 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_83
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_90
timestamp 1586364061
transform 1 0 9384 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _42_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_111
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_107
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_111
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_115
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_151
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_158
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_162
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_164
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_172
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 590 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 21436 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 21436 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_9
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_39
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_43
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _32_
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_55
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_61
timestamp 1586364061
transform 1 0 6716 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_12  FILLER_2_78
timestamp 1586364061
transform 1 0 8280 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_114
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_137
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use scs8hd_conb_1  _18_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_180
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_191
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_204
timestamp 1586364061
transform 1 0 19872 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 21436 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_212
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_6
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_18
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_26
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_69
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_91
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 774 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_108
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_119
timestamp 1586364061
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 866 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_167
timestamp 1586364061
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_181
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 21436 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_216
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_62
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_12  FILLER_4_79
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_130
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_137
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_174
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  FILLER_4_194
timestamp 1586364061
transform 1 0 18952 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 21436 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_6
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_49
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_81
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_85
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_89
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_93
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_106
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_182
timestamp 1586364061
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_192
timestamp 1586364061
transform 1 0 18768 0 1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_200
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 21436 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_216
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_9
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_9
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_19
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_13
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 590 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_58
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_73
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_106
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_120
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_134
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_129
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_146
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_146
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_162
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_158
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_165
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_174
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _16_
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_185
timestamp 1586364061
transform 1 0 18124 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_187
timestamp 1586364061
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_191
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 21436 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 21436 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_216
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _17_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_17
timestamp 1586364061
transform 1 0 2668 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_21
timestamp 1586364061
transform 1 0 3036 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_29
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_73
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use scs8hd_conb_1  _15_
timestamp 1586364061
transform 1 0 9752 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_109
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_130
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_162
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_188
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_194
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 21436 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_68
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_102
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_137
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 130 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_165
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_169
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_192
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 21436 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_28
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_38
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_42
timestamp 1586364061
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_79
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_113
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_157
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_168
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_173
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_184
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_201
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 21436 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_20
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_52
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_84
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_121
timestamp 1586364061
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 21436 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_20
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_28
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_35
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_12_47
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_63
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_12_66
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_76
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_108
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12328 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_142
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_176
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_193
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_12_204
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 21436 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_13
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_13
timestamp 1586364061
transform 1 0 2300 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_25
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_51
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_78
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_84
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_111
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_128
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_135
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_165
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 774 592
use scs8hd_conb_1  _19_
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_174
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_179
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_205
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_196
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 21436 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 21436 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_209
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_208
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_6
timestamp 1586364061
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_10
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_17
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_21
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_45
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_81
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_93
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 1142 592
use scs8hd_conb_1  _22_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_117
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_121
timestamp 1586364061
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_126
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_130
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_162
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_203
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 21436 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_209
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_213
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 130 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_18
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_6  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_126
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  FILLER_16_162
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_174
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_2  _33_
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_205
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 21436 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_70
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_78
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _30_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_127
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_131
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_155
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_163
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_167
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 406 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_17_187
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_198
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_203
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 21436 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_215
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_114
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_150
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_198
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_204
timestamp 1586364061
transform 1 0 19872 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 21436 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_212
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 774 592
use scs8hd_decap_4  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_155
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_161
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_177
timestamp 1586364061
transform 1 0 17388 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_189
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_201
timestamp 1586364061
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 21436 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 21436 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_215
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_213
timestamp 1586364061
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_103
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_21_115
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_150
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_158
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_180
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_21_192
timestamp 1586364061
transform 1 0 18768 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 21436 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_206
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_96
timestamp 1586364061
transform 1 0 9936 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_120
timestamp 1586364061
transform 1 0 12144 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_132
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_171
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_195
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 21436 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_207
timestamp 1586364061
transform 1 0 20148 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_70
timestamp 1586364061
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_104
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_148
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_152
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_202
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 21436 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_206
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_210
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_75
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_198
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 21436 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_72
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_107
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_25_192
timestamp 1586364061
transform 1 0 18768 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 21436 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_8
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_20
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_32
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_44
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_52
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_65
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_69
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_82
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_94
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_109
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_106
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_121
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_133
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_198
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 21436 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 21436 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_216
timestamp 1586364061
transform 1 0 20976 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_9
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_21
timestamp 1586364061
transform 1 0 3036 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_29
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 774 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 6072 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_58
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 1142 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_70
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 21436 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_19
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_31
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_43
timestamp 1586364061
transform 1 0 5060 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_75
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 406 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_111
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_119
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_200
timestamp 1586364061
transform 1 0 19504 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_203
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 21436 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_215
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 314 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_62
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_74
timestamp 1586364061
transform 1 0 7912 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_86
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_198
timestamp 1586364061
transform 1 0 19320 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_204
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 21436 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_208
timestamp 1586364061
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_153
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_157
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_161
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_169
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 21436 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_144
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_12  FILLER_32_180
timestamp 1586364061
transform 1 0 17664 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_192
timestamp 1586364061
transform 1 0 18768 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_32_196
timestamp 1586364061
transform 1 0 19136 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 21436 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_206
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_20
timestamp 1586364061
transform 1 0 2944 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_18
timestamp 1586364061
transform 1 0 2760 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_32
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_30
timestamp 1586364061
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_44
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_56
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _31_
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_82
timestamp 1586364061
transform 1 0 8648 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_90
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_96
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_107
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_108
timestamp 1586364061
transform 1 0 11040 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_124
timestamp 1586364061
transform 1 0 12512 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14076 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_131
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_134
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_138
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_135
timestamp 1586364061
transform 1 0 13524 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_33_150
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 590 592
use scs8hd_decap_6  FILLER_34_147
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_8  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_162
timestamp 1586364061
transform 1 0 16008 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_167
timestamp 1586364061
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_173
timestamp 1586364061
transform 1 0 17020 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_188
timestamp 1586364061
transform 1 0 18400 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_192
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_185
timestamp 1586364061
transform 1 0 18124 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_189
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_195
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_199
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 21436 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 21436 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_209
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_217
timestamp 1586364061
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_206
timestamp 1586364061
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_35_152
timestamp 1586364061
transform 1 0 15088 0 1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_163
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_167
timestamp 1586364061
transform 1 0 16468 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_174
timestamp 1586364061
transform 1 0 17112 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_178
timestamp 1586364061
transform 1 0 17480 0 1 21216
box -38 -48 406 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_182
timestamp 1586364061
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_190
timestamp 1586364061
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_195
timestamp 1586364061
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 21436 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_206
timestamp 1586364061
transform 1 0 20056 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_210
timestamp 1586364061
transform 1 0 20424 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_36_63
timestamp 1586364061
transform 1 0 6900 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_75
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_87
timestamp 1586364061
transform 1 0 9108 0 -1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_94
timestamp 1586364061
transform 1 0 9752 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 12512 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_118
timestamp 1586364061
transform 1 0 11960 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 15364 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_156
timestamp 1586364061
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_168
timestamp 1586364061
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 18216 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_180
timestamp 1586364061
transform 1 0 17664 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_36_187
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_199
timestamp 1586364061
transform 1 0 19412 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_204
timestamp 1586364061
transform 1 0 19872 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 21436 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 21068 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_216
timestamp 1586364061
transform 1 0 20976 0 -1 22304
box -38 -48 130 592
<< labels >>
rlabel metal2 s 1858 0 1914 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 2594 0 2650 480 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 688 480 808 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 2048 480 2168 6 address[3]
port 3 nsew default input
rlabel metal2 s 570 24210 626 24690 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 3408 480 3528 6 address[5]
port 5 nsew default input
rlabel metal2 s 1674 24210 1730 24690 6 address[6]
port 6 nsew default input
rlabel metal3 s 22066 688 22546 808 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal3 s 0 6128 480 6248 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal3 s 22066 3680 22546 3800 6 bottom_right_grid_pin_13_
port 9 nsew default input
rlabel metal2 s 4066 0 4122 480 6 bottom_right_grid_pin_15_
port 10 nsew default input
rlabel metal2 s 2870 24210 2926 24690 6 bottom_right_grid_pin_1_
port 11 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_right_grid_pin_3_
port 12 nsew default input
rlabel metal3 s 22066 2184 22546 2304 6 bottom_right_grid_pin_5_
port 13 nsew default input
rlabel metal3 s 0 4768 480 4888 6 bottom_right_grid_pin_7_
port 14 nsew default input
rlabel metal2 s 4066 24210 4122 24690 6 bottom_right_grid_pin_9_
port 15 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[0]
port 16 nsew default input
rlabel metal2 s 4894 0 4950 480 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal2 s 5630 0 5686 480 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 22066 5312 22546 5432 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal3 s 22066 6808 22546 6928 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal3 s 22066 8304 22546 8424 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal2 s 5262 24210 5318 24690 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal3 s 0 10208 480 10328 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chanx_left_out[0]
port 25 nsew default tristate
rlabel metal2 s 6458 24210 6514 24690 6 chanx_left_out[1]
port 26 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[2]
port 27 nsew default tristate
rlabel metal2 s 7654 24210 7710 24690 6 chanx_left_out[3]
port 28 nsew default tristate
rlabel metal3 s 22066 9936 22546 10056 6 chanx_left_out[4]
port 29 nsew default tristate
rlabel metal3 s 22066 11432 22546 11552 6 chanx_left_out[5]
port 30 nsew default tristate
rlabel metal2 s 7102 0 7158 480 6 chanx_left_out[6]
port 31 nsew default tristate
rlabel metal2 s 8850 24210 8906 24690 6 chanx_left_out[7]
port 32 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[8]
port 33 nsew default tristate
rlabel metal3 s 0 14424 480 14544 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal3 s 22066 13064 22546 13184 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal2 s 10046 24210 10102 24690 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal2 s 11242 24210 11298 24690 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal3 s 22066 14560 22546 14680 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal2 s 12346 24210 12402 24690 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal2 s 12346 0 12402 480 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal3 s 22066 16056 22546 16176 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal2 s 13542 24210 13598 24690 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal3 s 22066 17688 22546 17808 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chany_top_in[0]
port 52 nsew default input
rlabel metal2 s 14738 24210 14794 24690 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 15934 24210 15990 24690 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 17130 24210 17186 24690 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 14646 0 14702 480 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 16118 0 16174 480 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 18326 24210 18382 24690 6 chany_top_in[8]
port 60 nsew default input
rlabel metal3 s 0 18504 480 18624 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal3 s 22066 19184 22546 19304 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal2 s 16854 0 16910 480 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal2 s 19522 24210 19578 24690 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal2 s 20718 24210 20774 24690 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal2 s 18418 0 18474 480 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal2 s 1122 0 1178 480 6 data_in
port 70 nsew default input
rlabel metal2 s 386 0 442 480 6 enable
port 71 nsew default input
rlabel metal2 s 19890 0 19946 480 6 left_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal2 s 20626 0 20682 480 6 left_top_grid_pin_10_
port 73 nsew default input
rlabel metal2 s 21914 24210 21970 24690 6 top_left_grid_pin_13_
port 74 nsew default input
rlabel metal3 s 22066 20680 22546 20800 6 top_right_grid_pin_11_
port 75 nsew default input
rlabel metal3 s 22066 22312 22546 22432 6 top_right_grid_pin_13_
port 76 nsew default input
rlabel metal3 s 22066 23808 22546 23928 6 top_right_grid_pin_15_
port 77 nsew default input
rlabel metal3 s 0 21224 480 21344 6 top_right_grid_pin_1_
port 78 nsew default input
rlabel metal3 s 0 22584 480 22704 6 top_right_grid_pin_3_
port 79 nsew default input
rlabel metal3 s 0 23944 480 24064 6 top_right_grid_pin_5_
port 80 nsew default input
rlabel metal2 s 21362 0 21418 480 6 top_right_grid_pin_7_
port 81 nsew default input
rlabel metal2 s 22098 0 22154 480 6 top_right_grid_pin_9_
port 82 nsew default input
rlabel metal4 s 4702 2128 5022 22352 6 vpwr
port 83 nsew default input
rlabel metal4 s 8459 2128 8779 22352 6 vgnd
port 84 nsew default input
<< end >>
