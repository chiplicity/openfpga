magic
tech sky130A
magscale 1 2
timestamp 1605120228
<< locali >>
rect 3893 12699 3927 12801
rect 12081 8347 12115 8585
rect 4169 6715 4203 6953
<< viali >>
rect 18429 21097 18463 21131
rect 18245 20961 18279 20995
rect 19349 20961 19383 20995
rect 21649 20961 21683 20995
rect 19533 20825 19567 20859
rect 21833 20825 21867 20859
rect 8769 20553 8803 20587
rect 10241 20553 10275 20587
rect 13001 20553 13035 20587
rect 19349 20553 19383 20587
rect 21649 20553 21683 20587
rect 20545 20485 20579 20519
rect 23857 20485 23891 20519
rect 8585 20349 8619 20383
rect 12449 20349 12483 20383
rect 16313 20349 16347 20383
rect 16957 20349 16991 20383
rect 18061 20349 18095 20383
rect 18613 20349 18647 20383
rect 19165 20349 19199 20383
rect 19717 20349 19751 20383
rect 20361 20349 20395 20383
rect 20913 20349 20947 20383
rect 21833 20349 21867 20383
rect 23673 20349 23707 20383
rect 24225 20349 24259 20383
rect 20177 20281 20211 20315
rect 9229 20213 9263 20247
rect 12633 20213 12667 20247
rect 16497 20213 16531 20247
rect 18245 20213 18279 20247
rect 19073 20213 19107 20247
rect 22017 20213 22051 20247
rect 22385 20213 22419 20247
rect 21097 20009 21131 20043
rect 17325 19873 17359 19907
rect 19441 19873 19475 19907
rect 20913 19873 20947 19907
rect 17509 19737 17543 19771
rect 19625 19737 19659 19771
rect 17417 19397 17451 19431
rect 19441 19125 19475 19159
rect 20913 19125 20947 19159
rect 7665 14433 7699 14467
rect 8125 14433 8159 14467
rect 8217 14365 8251 14399
rect 8309 14365 8343 14399
rect 7757 14229 7791 14263
rect 8033 14025 8067 14059
rect 9413 14025 9447 14059
rect 8585 13889 8619 13923
rect 9045 13889 9079 13923
rect 7849 13821 7883 13855
rect 8493 13821 8527 13855
rect 7021 13753 7055 13787
rect 7573 13753 7607 13787
rect 8401 13753 8435 13787
rect 7113 13481 7147 13515
rect 7849 13481 7883 13515
rect 8033 13481 8067 13515
rect 8493 13481 8527 13515
rect 1409 13345 1443 13379
rect 8401 13345 8435 13379
rect 10241 13345 10275 13379
rect 10793 13345 10827 13379
rect 11060 13345 11094 13379
rect 13257 13345 13291 13379
rect 2329 13277 2363 13311
rect 2513 13277 2547 13311
rect 8585 13277 8619 13311
rect 13001 13277 13035 13311
rect 1593 13141 1627 13175
rect 9137 13141 9171 13175
rect 12173 13141 12207 13175
rect 14381 13141 14415 13175
rect 15485 13141 15519 13175
rect 1685 12937 1719 12971
rect 8125 12937 8159 12971
rect 8493 12937 8527 12971
rect 12725 12937 12759 12971
rect 15117 12937 15151 12971
rect 8585 12869 8619 12903
rect 2881 12801 2915 12835
rect 3249 12801 3283 12835
rect 3893 12801 3927 12835
rect 3985 12801 4019 12835
rect 7481 12801 7515 12835
rect 7573 12801 7607 12835
rect 9137 12801 9171 12835
rect 10149 12801 10183 12835
rect 13553 12801 13587 12835
rect 14105 12801 14139 12835
rect 14289 12801 14323 12835
rect 14657 12801 14691 12835
rect 15301 12801 15335 12835
rect 2605 12733 2639 12767
rect 3709 12733 3743 12767
rect 4169 12733 4203 12767
rect 7389 12733 7423 12767
rect 15557 12733 15591 12767
rect 2145 12665 2179 12699
rect 2697 12665 2731 12699
rect 3893 12665 3927 12699
rect 4414 12665 4448 12699
rect 6653 12665 6687 12699
rect 8953 12665 8987 12699
rect 10057 12665 10091 12699
rect 10394 12665 10428 12699
rect 13185 12665 13219 12699
rect 2237 12597 2271 12631
rect 5549 12597 5583 12631
rect 7021 12597 7055 12631
rect 9045 12597 9079 12631
rect 11529 12597 11563 12631
rect 13645 12597 13679 12631
rect 14013 12597 14047 12631
rect 16681 12597 16715 12631
rect 2789 12393 2823 12427
rect 7113 12393 7147 12427
rect 8125 12393 8159 12427
rect 8677 12393 8711 12427
rect 10885 12393 10919 12427
rect 11253 12393 11287 12427
rect 15301 12393 15335 12427
rect 17233 12393 17267 12427
rect 5150 12325 5184 12359
rect 14013 12325 14047 12359
rect 2697 12257 2731 12291
rect 10057 12257 10091 12291
rect 17785 12257 17819 12291
rect 2973 12189 3007 12223
rect 4905 12189 4939 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 17877 12189 17911 12223
rect 17969 12189 18003 12223
rect 18429 12189 18463 12223
rect 9045 12121 9079 12155
rect 9689 12121 9723 12155
rect 2053 12053 2087 12087
rect 2329 12053 2363 12087
rect 6285 12053 6319 12087
rect 13093 12053 13127 12087
rect 13645 12053 13679 12087
rect 16497 12053 16531 12087
rect 17417 12053 17451 12087
rect 1869 11849 1903 11883
rect 5273 11849 5307 11883
rect 11161 11849 11195 11883
rect 13185 11849 13219 11883
rect 13461 11849 13495 11883
rect 15301 11849 15335 11883
rect 16313 11849 16347 11883
rect 19073 11849 19107 11883
rect 4905 11781 4939 11815
rect 10793 11781 10827 11815
rect 2421 11713 2455 11747
rect 2605 11713 2639 11747
rect 6837 11713 6871 11747
rect 10333 11713 10367 11747
rect 13645 11713 13679 11747
rect 16957 11713 16991 11747
rect 17785 11713 17819 11747
rect 18613 11713 18647 11747
rect 2329 11645 2363 11679
rect 3709 11645 3743 11679
rect 10149 11645 10183 11679
rect 15945 11645 15979 11679
rect 16773 11645 16807 11679
rect 18521 11645 18555 11679
rect 26433 11645 26467 11679
rect 26985 11645 27019 11679
rect 6561 11577 6595 11611
rect 7082 11577 7116 11611
rect 9689 11577 9723 11611
rect 12817 11577 12851 11611
rect 13912 11577 13946 11611
rect 16865 11577 16899 11611
rect 1961 11509 1995 11543
rect 3065 11509 3099 11543
rect 3433 11509 3467 11543
rect 8217 11509 8251 11543
rect 8861 11509 8895 11543
rect 9229 11509 9263 11543
rect 9781 11509 9815 11543
rect 10241 11509 10275 11543
rect 15025 11509 15059 11543
rect 16405 11509 16439 11543
rect 17417 11509 17451 11543
rect 18061 11509 18095 11543
rect 18429 11509 18463 11543
rect 26617 11509 26651 11543
rect 2145 11305 2179 11339
rect 4537 11305 4571 11339
rect 6837 11305 6871 11339
rect 8769 11305 8803 11339
rect 9505 11305 9539 11339
rect 10149 11305 10183 11339
rect 13277 11305 13311 11339
rect 13737 11305 13771 11339
rect 16221 11305 16255 11339
rect 17325 11305 17359 11339
rect 2053 11237 2087 11271
rect 16129 11237 16163 11271
rect 18337 11237 18371 11271
rect 1685 11169 1719 11203
rect 2513 11169 2547 11203
rect 4445 11169 4479 11203
rect 7389 11169 7423 11203
rect 7645 11169 7679 11203
rect 13829 11169 13863 11203
rect 14473 11169 14507 11203
rect 17693 11169 17727 11203
rect 26525 11169 26559 11203
rect 2605 11101 2639 11135
rect 2697 11101 2731 11135
rect 4629 11101 4663 11135
rect 10241 11101 10275 11135
rect 10333 11101 10367 11135
rect 13921 11101 13955 11135
rect 16405 11101 16439 11135
rect 17785 11101 17819 11135
rect 17969 11101 18003 11135
rect 4077 11033 4111 11067
rect 9781 11033 9815 11067
rect 26709 11033 26743 11067
rect 3249 10965 3283 10999
rect 13369 10965 13403 10999
rect 15761 10965 15795 10999
rect 1593 10761 1627 10795
rect 2421 10761 2455 10795
rect 2881 10761 2915 10795
rect 4169 10761 4203 10795
rect 7481 10761 7515 10795
rect 8953 10761 8987 10795
rect 9689 10761 9723 10795
rect 9781 10761 9815 10795
rect 14381 10761 14415 10795
rect 15209 10761 15243 10795
rect 17049 10761 17083 10795
rect 27353 10761 27387 10795
rect 4445 10693 4479 10727
rect 7757 10693 7791 10727
rect 2053 10625 2087 10659
rect 2789 10625 2823 10659
rect 3525 10625 3559 10659
rect 4813 10625 4847 10659
rect 10333 10625 10367 10659
rect 11161 10625 11195 10659
rect 11529 10625 11563 10659
rect 13277 10625 13311 10659
rect 13921 10625 13955 10659
rect 14841 10625 14875 10659
rect 16221 10625 16255 10659
rect 1409 10557 1443 10591
rect 10241 10557 10275 10591
rect 15577 10557 15611 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 26433 10557 26467 10591
rect 26985 10557 27019 10591
rect 3249 10489 3283 10523
rect 10793 10489 10827 10523
rect 13829 10489 13863 10523
rect 3341 10421 3375 10455
rect 9229 10421 9263 10455
rect 10149 10421 10183 10455
rect 12909 10421 12943 10455
rect 13369 10421 13403 10455
rect 13737 10421 13771 10455
rect 15669 10421 15703 10455
rect 17417 10421 17451 10455
rect 17693 10421 17727 10455
rect 26617 10421 26651 10455
rect 2329 10217 2363 10251
rect 6101 10217 6135 10251
rect 6929 10217 6963 10251
rect 9689 10217 9723 10251
rect 10149 10217 10183 10251
rect 12909 10217 12943 10251
rect 14381 10217 14415 10251
rect 16497 10217 16531 10251
rect 1869 10149 1903 10183
rect 15853 10149 15887 10183
rect 16221 10149 16255 10183
rect 2697 10081 2731 10115
rect 4988 10081 5022 10115
rect 7113 10081 7147 10115
rect 10057 10081 10091 10115
rect 13001 10081 13035 10115
rect 13257 10081 13291 10115
rect 2237 10013 2271 10047
rect 2789 10013 2823 10047
rect 2973 10013 3007 10047
rect 4721 10013 4755 10047
rect 10333 10013 10367 10047
rect 3433 9877 3467 9911
rect 4629 9877 4663 9911
rect 8585 9877 8619 9911
rect 10425 9673 10459 9707
rect 13093 9673 13127 9707
rect 13461 9673 13495 9707
rect 14105 9673 14139 9707
rect 1593 9605 1627 9639
rect 2053 9605 2087 9639
rect 2973 9605 3007 9639
rect 4537 9605 4571 9639
rect 6009 9605 6043 9639
rect 10149 9605 10183 9639
rect 3617 9537 3651 9571
rect 4077 9537 4111 9571
rect 5181 9537 5215 9571
rect 9045 9537 9079 9571
rect 9229 9537 9263 9571
rect 14197 9537 14231 9571
rect 1409 9469 1443 9503
rect 4445 9469 4479 9503
rect 4997 9469 5031 9503
rect 8125 9469 8159 9503
rect 12265 9469 12299 9503
rect 12633 9469 12667 9503
rect 2881 9401 2915 9435
rect 8401 9401 8435 9435
rect 14442 9401 14476 9435
rect 2421 9333 2455 9367
rect 3341 9333 3375 9367
rect 3433 9333 3467 9367
rect 4905 9333 4939 9367
rect 5549 9333 5583 9367
rect 7021 9333 7055 9367
rect 8585 9333 8619 9367
rect 8953 9333 8987 9367
rect 9781 9333 9815 9367
rect 12081 9333 12115 9367
rect 15577 9333 15611 9367
rect 1593 9129 1627 9163
rect 2421 9129 2455 9163
rect 4077 9129 4111 9163
rect 4537 9129 4571 9163
rect 8493 9129 8527 9163
rect 9689 9129 9723 9163
rect 13461 9129 13495 9163
rect 14197 9129 14231 9163
rect 26709 9129 26743 9163
rect 3433 9061 3467 9095
rect 8401 9061 8435 9095
rect 1409 8993 1443 9027
rect 4445 8993 4479 9027
rect 10057 8993 10091 9027
rect 11345 8993 11379 9027
rect 11612 8993 11646 9027
rect 26525 8993 26559 9027
rect 4721 8925 4755 8959
rect 5641 8925 5675 8959
rect 8585 8925 8619 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 13093 8857 13127 8891
rect 3065 8789 3099 8823
rect 5181 8789 5215 8823
rect 8033 8789 8067 8823
rect 9229 8789 9263 8823
rect 12725 8789 12759 8823
rect 1593 8585 1627 8619
rect 2329 8585 2363 8619
rect 3157 8585 3191 8619
rect 3801 8585 3835 8619
rect 4169 8585 4203 8619
rect 7481 8585 7515 8619
rect 8125 8585 8159 8619
rect 8493 8585 8527 8619
rect 12081 8585 12115 8619
rect 12173 8585 12207 8619
rect 27353 8585 27387 8619
rect 2697 8517 2731 8551
rect 7573 8517 7607 8551
rect 2053 8449 2087 8483
rect 5825 8449 5859 8483
rect 9045 8449 9079 8483
rect 1409 8381 1443 8415
rect 2513 8381 2547 8415
rect 5089 8381 5123 8415
rect 5549 8381 5583 8415
rect 7757 8381 7791 8415
rect 26617 8517 26651 8551
rect 27721 8517 27755 8551
rect 13369 8449 13403 8483
rect 13093 8381 13127 8415
rect 26433 8381 26467 8415
rect 26985 8381 27019 8415
rect 27537 8381 27571 8415
rect 28089 8381 28123 8415
rect 4445 8313 4479 8347
rect 5641 8313 5675 8347
rect 9229 8313 9263 8347
rect 10977 8313 11011 8347
rect 12081 8313 12115 8347
rect 13185 8313 13219 8347
rect 5181 8245 5215 8279
rect 6285 8245 6319 8279
rect 11437 8245 11471 8279
rect 11805 8245 11839 8279
rect 12725 8245 12759 8279
rect 16129 8245 16163 8279
rect 1593 8041 1627 8075
rect 5457 8041 5491 8075
rect 6653 8041 6687 8075
rect 7665 8041 7699 8075
rect 7849 8041 7883 8075
rect 9873 8041 9907 8075
rect 11437 8041 11471 8075
rect 12081 8041 12115 8075
rect 12541 8041 12575 8075
rect 13093 8041 13127 8075
rect 16221 8041 16255 8075
rect 26709 8041 26743 8075
rect 6745 7973 6779 8007
rect 1409 7905 1443 7939
rect 4333 7905 4367 7939
rect 8392 7905 8426 7939
rect 13185 7905 13219 7939
rect 26525 7905 26559 7939
rect 4077 7837 4111 7871
rect 6929 7837 6963 7871
rect 8125 7837 8159 7871
rect 11529 7837 11563 7871
rect 11621 7837 11655 7871
rect 13369 7837 13403 7871
rect 16313 7837 16347 7871
rect 16497 7837 16531 7871
rect 10333 7769 10367 7803
rect 2973 7701 3007 7735
rect 6285 7701 6319 7735
rect 9505 7701 9539 7735
rect 10701 7701 10735 7735
rect 11069 7701 11103 7735
rect 12725 7701 12759 7735
rect 15853 7701 15887 7735
rect 2421 7497 2455 7531
rect 6377 7497 6411 7531
rect 7021 7497 7055 7531
rect 7849 7497 7883 7531
rect 8585 7497 8619 7531
rect 11621 7497 11655 7531
rect 11805 7497 11839 7531
rect 15117 7497 15151 7531
rect 27353 7497 27387 7531
rect 1593 7429 1627 7463
rect 9781 7429 9815 7463
rect 15393 7429 15427 7463
rect 15761 7429 15795 7463
rect 2973 7361 3007 7395
rect 5089 7361 5123 7395
rect 5825 7361 5859 7395
rect 9229 7361 9263 7395
rect 10701 7361 10735 7395
rect 10885 7361 10919 7395
rect 12909 7361 12943 7395
rect 13001 7361 13035 7395
rect 16405 7361 16439 7395
rect 16589 7361 16623 7395
rect 1409 7293 1443 7327
rect 3240 7293 3274 7327
rect 5549 7293 5583 7327
rect 8217 7293 8251 7327
rect 9137 7293 9171 7327
rect 10149 7293 10183 7327
rect 10609 7293 10643 7327
rect 11989 7293 12023 7327
rect 12817 7293 12851 7327
rect 13829 7293 13863 7327
rect 16313 7293 16347 7327
rect 26433 7293 26467 7327
rect 26985 7293 27019 7327
rect 2881 7225 2915 7259
rect 9045 7225 9079 7259
rect 14197 7225 14231 7259
rect 2053 7157 2087 7191
rect 4353 7157 4387 7191
rect 4629 7157 4663 7191
rect 5181 7157 5215 7191
rect 5641 7157 5675 7191
rect 7389 7157 7423 7191
rect 8677 7157 8711 7191
rect 10241 7157 10275 7191
rect 11345 7157 11379 7191
rect 12449 7157 12483 7191
rect 13461 7157 13495 7191
rect 15945 7157 15979 7191
rect 16957 7157 16991 7191
rect 26617 7157 26651 7191
rect 4169 6953 4203 6987
rect 4261 6953 4295 6987
rect 5641 6953 5675 6987
rect 9045 6953 9079 6987
rect 10057 6953 10091 6987
rect 11161 6953 11195 6987
rect 11897 6953 11931 6987
rect 12817 6953 12851 6987
rect 13185 6953 13219 6987
rect 15117 6953 15151 6987
rect 15669 6953 15703 6987
rect 16313 6953 16347 6987
rect 1409 6817 1443 6851
rect 2513 6817 2547 6851
rect 3157 6817 3191 6851
rect 15761 6885 15795 6919
rect 5181 6817 5215 6851
rect 6193 6817 6227 6851
rect 6633 6817 6667 6851
rect 8769 6817 8803 6851
rect 26525 6817 26559 6851
rect 6377 6749 6411 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 15853 6749 15887 6783
rect 1593 6681 1627 6715
rect 4169 6681 4203 6715
rect 6009 6681 6043 6715
rect 7757 6681 7791 6715
rect 26709 6681 26743 6715
rect 2697 6613 2731 6647
rect 9689 6613 9723 6647
rect 13737 6613 13771 6647
rect 15301 6613 15335 6647
rect 16681 6613 16715 6647
rect 17049 6613 17083 6647
rect 1961 6409 1995 6443
rect 2513 6409 2547 6443
rect 6101 6409 6135 6443
rect 8769 6409 8803 6443
rect 10333 6409 10367 6443
rect 15117 6409 15151 6443
rect 15485 6409 15519 6443
rect 7021 6341 7055 6375
rect 10609 6341 10643 6375
rect 2973 6273 3007 6307
rect 3617 6273 3651 6307
rect 10977 6273 11011 6307
rect 13737 6273 13771 6307
rect 16773 6273 16807 6307
rect 1409 6205 1443 6239
rect 3433 6205 3467 6239
rect 8953 6205 8987 6239
rect 9209 6205 9243 6239
rect 12265 6205 12299 6239
rect 12633 6205 12667 6239
rect 16589 6205 16623 6239
rect 26525 6205 26559 6239
rect 13645 6137 13679 6171
rect 13982 6137 14016 6171
rect 1593 6069 1627 6103
rect 3065 6069 3099 6103
rect 3525 6069 3559 6103
rect 6377 6069 6411 6103
rect 12081 6069 12115 6103
rect 16037 6069 16071 6103
rect 16221 6069 16255 6103
rect 16681 6069 16715 6103
rect 17233 6069 17267 6103
rect 2053 5865 2087 5899
rect 3157 5865 3191 5899
rect 4077 5865 4111 5899
rect 6101 5865 6135 5899
rect 8953 5865 8987 5899
rect 9965 5865 9999 5899
rect 13921 5865 13955 5899
rect 15117 5865 15151 5899
rect 16865 5865 16899 5899
rect 17325 5865 17359 5899
rect 26709 5865 26743 5899
rect 6009 5797 6043 5831
rect 10578 5797 10612 5831
rect 12786 5797 12820 5831
rect 1409 5729 1443 5763
rect 3893 5729 3927 5763
rect 4445 5729 4479 5763
rect 10333 5729 10367 5763
rect 15669 5729 15703 5763
rect 17233 5729 17267 5763
rect 26525 5729 26559 5763
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 6285 5661 6319 5695
rect 12541 5661 12575 5695
rect 15761 5661 15795 5695
rect 15853 5661 15887 5695
rect 17417 5661 17451 5695
rect 16405 5593 16439 5627
rect 1593 5525 1627 5559
rect 5181 5525 5215 5559
rect 5641 5525 5675 5559
rect 11713 5525 11747 5559
rect 14197 5525 14231 5559
rect 15301 5525 15335 5559
rect 2421 5321 2455 5355
rect 3525 5321 3559 5355
rect 4353 5321 4387 5355
rect 5733 5321 5767 5355
rect 6377 5321 6411 5355
rect 10333 5321 10367 5355
rect 10701 5321 10735 5355
rect 12633 5321 12667 5355
rect 15761 5321 15795 5355
rect 16405 5321 16439 5355
rect 17785 5321 17819 5355
rect 26617 5321 26651 5355
rect 3893 5253 3927 5287
rect 6101 5253 6135 5287
rect 16313 5253 16347 5287
rect 17509 5253 17543 5287
rect 4813 5185 4847 5219
rect 4905 5185 4939 5219
rect 13553 5185 13587 5219
rect 16957 5185 16991 5219
rect 1409 5117 1443 5151
rect 4261 5117 4295 5151
rect 4721 5117 4755 5151
rect 13645 5117 13679 5151
rect 13912 5117 13946 5151
rect 16773 5117 16807 5151
rect 26433 5117 26467 5151
rect 26985 5117 27019 5151
rect 16865 5049 16899 5083
rect 1593 4981 1627 5015
rect 2053 4981 2087 5015
rect 13093 4981 13127 5015
rect 15025 4981 15059 5015
rect 15393 4981 15427 5015
rect 26341 4981 26375 5015
rect 2053 4777 2087 4811
rect 3893 4777 3927 4811
rect 4261 4777 4295 4811
rect 7389 4777 7423 4811
rect 10241 4777 10275 4811
rect 14013 4777 14047 4811
rect 15577 4777 15611 4811
rect 16681 4777 16715 4811
rect 17141 4777 17175 4811
rect 26709 4777 26743 4811
rect 4629 4709 4663 4743
rect 5365 4709 5399 4743
rect 6276 4709 6310 4743
rect 16405 4709 16439 4743
rect 17049 4709 17083 4743
rect 1409 4641 1443 4675
rect 2513 4641 2547 4675
rect 6009 4641 6043 4675
rect 10517 4641 10551 4675
rect 17693 4641 17727 4675
rect 26525 4641 26559 4675
rect 4721 4573 4755 4607
rect 4905 4573 4939 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 17233 4573 17267 4607
rect 2697 4505 2731 4539
rect 1593 4437 1627 4471
rect 10701 4437 10735 4471
rect 13645 4437 13679 4471
rect 6193 4233 6227 4267
rect 6469 4233 6503 4267
rect 14105 4233 14139 4267
rect 15209 4233 15243 4267
rect 17049 4233 17083 4267
rect 17417 4233 17451 4267
rect 27353 4233 27387 4267
rect 15117 4165 15151 4199
rect 16773 4165 16807 4199
rect 2421 4097 2455 4131
rect 3065 4097 3099 4131
rect 4261 4097 4295 4131
rect 5365 4097 5399 4131
rect 13737 4097 13771 4131
rect 14749 4097 14783 4131
rect 15761 4097 15795 4131
rect 1409 4029 1443 4063
rect 2513 4029 2547 4063
rect 3617 4029 3651 4063
rect 4537 4029 4571 4063
rect 5089 4029 5123 4063
rect 5733 4029 5767 4063
rect 10149 4029 10183 4063
rect 10416 4029 10450 4063
rect 15577 4029 15611 4063
rect 15669 4029 15703 4063
rect 26433 4029 26467 4063
rect 26985 4029 27019 4063
rect 2053 3961 2087 3995
rect 3525 3961 3559 3995
rect 5181 3961 5215 3995
rect 10057 3961 10091 3995
rect 13369 3961 13403 3995
rect 1593 3893 1627 3927
rect 2697 3893 2731 3927
rect 3801 3893 3835 3927
rect 4721 3893 4755 3927
rect 11529 3893 11563 3927
rect 26617 3893 26651 3927
rect 3893 3689 3927 3723
rect 5089 3689 5123 3723
rect 10609 3689 10643 3723
rect 15485 3689 15519 3723
rect 26709 3689 26743 3723
rect 4353 3621 4387 3655
rect 1409 3553 1443 3587
rect 2697 3553 2731 3587
rect 11529 3553 11563 3587
rect 11796 3553 11830 3587
rect 15853 3553 15887 3587
rect 25329 3553 25363 3587
rect 26525 3553 26559 3587
rect 1593 3485 1627 3519
rect 5181 3485 5215 3519
rect 5365 3485 5399 3519
rect 4721 3417 4755 3451
rect 9873 3417 9907 3451
rect 2881 3349 2915 3383
rect 12909 3349 12943 3383
rect 13185 3349 13219 3383
rect 16037 3349 16071 3383
rect 25513 3349 25547 3383
rect 1777 3145 1811 3179
rect 2789 3145 2823 3179
rect 3801 3145 3835 3179
rect 4813 3145 4847 3179
rect 5825 3145 5859 3179
rect 8861 3145 8895 3179
rect 25145 3145 25179 3179
rect 25881 3145 25915 3179
rect 26617 3145 26651 3179
rect 27353 3145 27387 3179
rect 4445 3077 4479 3111
rect 12173 3077 12207 3111
rect 6285 3009 6319 3043
rect 1869 2941 1903 2975
rect 3157 2941 3191 2975
rect 5089 2941 5123 2975
rect 8033 2941 8067 2975
rect 10149 2941 10183 2975
rect 13093 2941 13127 2975
rect 15209 2941 15243 2975
rect 15301 2941 15335 2975
rect 18245 2941 18279 2975
rect 18797 2941 18831 2975
rect 25329 2941 25363 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 27537 2941 27571 2975
rect 28089 2941 28123 2975
rect 2145 2873 2179 2907
rect 5365 2873 5399 2907
rect 8309 2873 8343 2907
rect 10057 2873 10091 2907
rect 10416 2873 10450 2907
rect 12909 2873 12943 2907
rect 13338 2873 13372 2907
rect 15546 2873 15580 2907
rect 3341 2805 3375 2839
rect 11529 2805 11563 2839
rect 11805 2805 11839 2839
rect 14473 2805 14507 2839
rect 14749 2805 14783 2839
rect 16681 2805 16715 2839
rect 17049 2805 17083 2839
rect 18429 2805 18463 2839
rect 25513 2805 25547 2839
rect 27721 2805 27755 2839
rect 1685 2601 1719 2635
rect 2789 2601 2823 2635
rect 6009 2601 6043 2635
rect 8309 2601 8343 2635
rect 10241 2601 10275 2635
rect 10885 2601 10919 2635
rect 11621 2601 11655 2635
rect 13829 2601 13863 2635
rect 16865 2601 16899 2635
rect 17141 2601 17175 2635
rect 19625 2601 19659 2635
rect 23029 2601 23063 2635
rect 7757 2533 7791 2567
rect 14933 2533 14967 2567
rect 15301 2533 15335 2567
rect 15752 2533 15786 2567
rect 1961 2465 1995 2499
rect 4537 2465 4571 2499
rect 4896 2465 4930 2499
rect 7481 2465 7515 2499
rect 10333 2465 10367 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 13185 2465 13219 2499
rect 14289 2465 14323 2499
rect 15485 2465 15519 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 19441 2465 19475 2499
rect 19993 2465 20027 2499
rect 22845 2465 22879 2499
rect 23397 2465 23431 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 25697 2465 25731 2499
rect 26249 2465 26283 2499
rect 26893 2465 26927 2499
rect 27445 2465 27479 2499
rect 2237 2397 2271 2431
rect 3893 2397 3927 2431
rect 4629 2397 4663 2431
rect 10517 2329 10551 2363
rect 14473 2329 14507 2363
rect 18521 2329 18555 2363
rect 13369 2261 13403 2295
rect 24777 2261 24811 2295
rect 25881 2261 25915 2295
rect 27077 2261 27111 2295
<< metal1 >>
rect 3326 22516 3332 22568
rect 3384 22556 3390 22568
rect 7650 22556 7656 22568
rect 3384 22528 7656 22556
rect 3384 22516 3390 22528
rect 7650 22516 7656 22528
rect 7708 22516 7714 22568
rect 4062 22108 4068 22160
rect 4120 22148 4126 22160
rect 13446 22148 13452 22160
rect 4120 22120 13452 22148
rect 4120 22108 4126 22120
rect 13446 22108 13452 22120
rect 13504 22108 13510 22160
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 3694 21088 3700 21140
rect 3752 21128 3758 21140
rect 18417 21131 18475 21137
rect 18417 21128 18429 21131
rect 3752 21100 18429 21128
rect 3752 21088 3758 21100
rect 18417 21097 18429 21100
rect 18463 21097 18475 21131
rect 18417 21091 18475 21097
rect 6362 21020 6368 21072
rect 6420 21060 6426 21072
rect 25590 21060 25596 21072
rect 6420 21032 25596 21060
rect 6420 21020 6426 21032
rect 25590 21020 25596 21032
rect 25648 21020 25654 21072
rect 3878 20952 3884 21004
rect 3936 20992 3942 21004
rect 15838 20992 15844 21004
rect 3936 20964 15844 20992
rect 3936 20952 3942 20964
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 18233 20995 18291 21001
rect 18233 20961 18245 20995
rect 18279 20992 18291 20995
rect 19058 20992 19064 21004
rect 18279 20964 19064 20992
rect 18279 20961 18291 20964
rect 18233 20955 18291 20961
rect 19058 20952 19064 20964
rect 19116 20952 19122 21004
rect 19337 20995 19395 21001
rect 19337 20961 19349 20995
rect 19383 20992 19395 20995
rect 19518 20992 19524 21004
rect 19383 20964 19524 20992
rect 19383 20961 19395 20964
rect 19337 20955 19395 20961
rect 19518 20952 19524 20964
rect 19576 20952 19582 21004
rect 21634 20992 21640 21004
rect 21595 20964 21640 20992
rect 21634 20952 21640 20964
rect 21692 20952 21698 21004
rect 8202 20884 8208 20936
rect 8260 20924 8266 20936
rect 8260 20896 21864 20924
rect 8260 20884 8266 20896
rect 5166 20816 5172 20868
rect 5224 20856 5230 20868
rect 21836 20865 21864 20896
rect 19521 20859 19579 20865
rect 19521 20856 19533 20859
rect 5224 20828 19533 20856
rect 5224 20816 5230 20828
rect 19521 20825 19533 20828
rect 19567 20825 19579 20859
rect 19521 20819 19579 20825
rect 21821 20859 21879 20865
rect 21821 20825 21833 20859
rect 21867 20825 21879 20859
rect 21821 20819 21879 20825
rect 3326 20748 3332 20800
rect 3384 20788 3390 20800
rect 5074 20788 5080 20800
rect 3384 20760 5080 20788
rect 3384 20748 3390 20760
rect 5074 20748 5080 20760
rect 5132 20748 5138 20800
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 8757 20587 8815 20593
rect 8757 20553 8769 20587
rect 8803 20584 8815 20587
rect 9582 20584 9588 20596
rect 8803 20556 9588 20584
rect 8803 20553 8815 20556
rect 8757 20547 8815 20553
rect 9582 20544 9588 20556
rect 9640 20544 9646 20596
rect 10229 20587 10287 20593
rect 10229 20553 10241 20587
rect 10275 20584 10287 20587
rect 11330 20584 11336 20596
rect 10275 20556 11336 20584
rect 10275 20553 10287 20556
rect 10229 20547 10287 20553
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 12710 20544 12716 20596
rect 12768 20584 12774 20596
rect 12989 20587 13047 20593
rect 12989 20584 13001 20587
rect 12768 20556 13001 20584
rect 12768 20544 12774 20556
rect 12989 20553 13001 20556
rect 13035 20553 13047 20587
rect 12989 20547 13047 20553
rect 19337 20587 19395 20593
rect 19337 20553 19349 20587
rect 19383 20584 19395 20587
rect 19426 20584 19432 20596
rect 19383 20556 19432 20584
rect 19383 20553 19395 20556
rect 19337 20547 19395 20553
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 21634 20584 21640 20596
rect 21595 20556 21640 20584
rect 21634 20544 21640 20556
rect 21692 20544 21698 20596
rect 20530 20516 20536 20528
rect 20491 20488 20536 20516
rect 20530 20476 20536 20488
rect 20588 20476 20594 20528
rect 23842 20516 23848 20528
rect 23803 20488 23848 20516
rect 23842 20476 23848 20488
rect 23900 20476 23906 20528
rect 25130 20408 25136 20460
rect 25188 20448 25194 20460
rect 25866 20448 25872 20460
rect 25188 20420 25872 20448
rect 25188 20408 25194 20420
rect 25866 20408 25872 20420
rect 25924 20408 25930 20460
rect 8573 20383 8631 20389
rect 8573 20349 8585 20383
rect 8619 20380 8631 20383
rect 12437 20383 12495 20389
rect 8619 20352 9260 20380
rect 8619 20349 8631 20352
rect 8573 20343 8631 20349
rect 9232 20256 9260 20352
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 12710 20380 12716 20392
rect 12483 20352 12716 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 12710 20340 12716 20352
rect 12768 20340 12774 20392
rect 16301 20383 16359 20389
rect 16301 20349 16313 20383
rect 16347 20380 16359 20383
rect 16945 20383 17003 20389
rect 16945 20380 16957 20383
rect 16347 20352 16957 20380
rect 16347 20349 16359 20352
rect 16301 20343 16359 20349
rect 16945 20349 16957 20352
rect 16991 20380 17003 20383
rect 18046 20380 18052 20392
rect 16991 20352 18052 20380
rect 16991 20349 17003 20352
rect 16945 20343 17003 20349
rect 18046 20340 18052 20352
rect 18104 20380 18110 20392
rect 18601 20383 18659 20389
rect 18601 20380 18613 20383
rect 18104 20352 18613 20380
rect 18104 20340 18110 20352
rect 18601 20349 18613 20352
rect 18647 20349 18659 20383
rect 19150 20380 19156 20392
rect 19111 20352 19156 20380
rect 18601 20343 18659 20349
rect 19150 20340 19156 20352
rect 19208 20380 19214 20392
rect 19705 20383 19763 20389
rect 19705 20380 19717 20383
rect 19208 20352 19717 20380
rect 19208 20340 19214 20352
rect 19705 20349 19717 20352
rect 19751 20349 19763 20383
rect 19705 20343 19763 20349
rect 20349 20383 20407 20389
rect 20349 20349 20361 20383
rect 20395 20380 20407 20383
rect 20901 20383 20959 20389
rect 20901 20380 20913 20383
rect 20395 20352 20913 20380
rect 20395 20349 20407 20352
rect 20349 20343 20407 20349
rect 20901 20349 20913 20352
rect 20947 20380 20959 20383
rect 21821 20383 21879 20389
rect 21821 20380 21833 20383
rect 20947 20352 21833 20380
rect 20947 20349 20959 20352
rect 20901 20343 20959 20349
rect 21821 20349 21833 20352
rect 21867 20380 21879 20383
rect 23658 20380 23664 20392
rect 21867 20352 22416 20380
rect 23619 20352 23664 20380
rect 21867 20349 21879 20352
rect 21821 20343 21879 20349
rect 19518 20272 19524 20324
rect 19576 20312 19582 20324
rect 20165 20315 20223 20321
rect 20165 20312 20177 20315
rect 19576 20284 20177 20312
rect 19576 20272 19582 20284
rect 20165 20281 20177 20284
rect 20211 20312 20223 20315
rect 20714 20312 20720 20324
rect 20211 20284 20720 20312
rect 20211 20281 20223 20284
rect 20165 20275 20223 20281
rect 20714 20272 20720 20284
rect 20772 20272 20778 20324
rect 21634 20272 21640 20324
rect 21692 20312 21698 20324
rect 22094 20312 22100 20324
rect 21692 20284 22100 20312
rect 21692 20272 21698 20284
rect 22094 20272 22100 20284
rect 22152 20272 22158 20324
rect 22388 20256 22416 20352
rect 23658 20340 23664 20352
rect 23716 20380 23722 20392
rect 24213 20383 24271 20389
rect 24213 20380 24225 20383
rect 23716 20352 24225 20380
rect 23716 20340 23722 20352
rect 24213 20349 24225 20352
rect 24259 20349 24271 20383
rect 24213 20343 24271 20349
rect 9214 20244 9220 20256
rect 9175 20216 9220 20244
rect 9214 20204 9220 20216
rect 9272 20204 9278 20256
rect 12621 20247 12679 20253
rect 12621 20213 12633 20247
rect 12667 20244 12679 20247
rect 13078 20244 13084 20256
rect 12667 20216 13084 20244
rect 12667 20213 12679 20216
rect 12621 20207 12679 20213
rect 13078 20204 13084 20216
rect 13136 20204 13142 20256
rect 16482 20244 16488 20256
rect 16443 20216 16488 20244
rect 16482 20204 16488 20216
rect 16540 20204 16546 20256
rect 18230 20244 18236 20256
rect 18191 20216 18236 20244
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 19058 20244 19064 20256
rect 18971 20216 19064 20244
rect 19058 20204 19064 20216
rect 19116 20244 19122 20256
rect 19426 20244 19432 20256
rect 19116 20216 19432 20244
rect 19116 20204 19122 20216
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 22002 20244 22008 20256
rect 21963 20216 22008 20244
rect 22002 20204 22008 20216
rect 22060 20204 22066 20256
rect 22370 20244 22376 20256
rect 22331 20216 22376 20244
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 21085 20043 21143 20049
rect 21085 20009 21097 20043
rect 21131 20040 21143 20043
rect 21542 20040 21548 20052
rect 21131 20012 21548 20040
rect 21131 20009 21143 20012
rect 21085 20003 21143 20009
rect 21542 20000 21548 20012
rect 21600 20000 21606 20052
rect 17310 19904 17316 19916
rect 17271 19876 17316 19904
rect 17310 19864 17316 19876
rect 17368 19864 17374 19916
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 20714 19864 20720 19916
rect 20772 19904 20778 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20772 19876 20913 19904
rect 20772 19864 20778 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 17494 19768 17500 19780
rect 17455 19740 17500 19768
rect 17494 19728 17500 19740
rect 17552 19728 17558 19780
rect 19610 19768 19616 19780
rect 19571 19740 19616 19768
rect 19610 19728 19616 19740
rect 19668 19728 19674 19780
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 17310 19388 17316 19440
rect 17368 19428 17374 19440
rect 17405 19431 17463 19437
rect 17405 19428 17417 19431
rect 17368 19400 17417 19428
rect 17368 19388 17374 19400
rect 17405 19397 17417 19400
rect 17451 19428 17463 19431
rect 19150 19428 19156 19440
rect 17451 19400 19156 19428
rect 17451 19397 17463 19400
rect 17405 19391 17463 19397
rect 19150 19388 19156 19400
rect 19208 19388 19214 19440
rect 15746 19320 15752 19372
rect 15804 19360 15810 19372
rect 16482 19360 16488 19372
rect 15804 19332 16488 19360
rect 15804 19320 15810 19332
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 17218 19320 17224 19372
rect 17276 19360 17282 19372
rect 17862 19360 17868 19372
rect 17276 19332 17868 19360
rect 17276 19320 17282 19332
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 18690 19320 18696 19372
rect 18748 19360 18754 19372
rect 19242 19360 19248 19372
rect 18748 19332 19248 19360
rect 18748 19320 18754 19332
rect 19242 19320 19248 19332
rect 19300 19320 19306 19372
rect 19426 19156 19432 19168
rect 19339 19128 19432 19156
rect 19426 19116 19432 19128
rect 19484 19156 19490 19168
rect 19702 19156 19708 19168
rect 19484 19128 19708 19156
rect 19484 19116 19490 19128
rect 19702 19116 19708 19128
rect 19760 19116 19766 19168
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 20901 19159 20959 19165
rect 20901 19156 20913 19159
rect 20772 19128 20913 19156
rect 20772 19116 20778 19128
rect 20901 19125 20913 19128
rect 20947 19125 20959 19159
rect 20901 19119 20959 19125
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 29362 18748 29368 18760
rect 19392 18720 29368 18748
rect 19392 18708 19398 18720
rect 29362 18708 29368 18720
rect 29420 18708 29426 18760
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 7653 14467 7711 14473
rect 7653 14433 7665 14467
rect 7699 14464 7711 14467
rect 8018 14464 8024 14476
rect 7699 14436 8024 14464
rect 7699 14433 7711 14436
rect 7653 14427 7711 14433
rect 8018 14424 8024 14436
rect 8076 14464 8082 14476
rect 8113 14467 8171 14473
rect 8113 14464 8125 14467
rect 8076 14436 8125 14464
rect 8076 14424 8082 14436
rect 8113 14433 8125 14436
rect 8159 14433 8171 14467
rect 8113 14427 8171 14433
rect 8202 14396 8208 14408
rect 8163 14368 8208 14396
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14365 8355 14399
rect 8297 14359 8355 14365
rect 7926 14288 7932 14340
rect 7984 14328 7990 14340
rect 8312 14328 8340 14359
rect 7984 14300 8340 14328
rect 7984 14288 7990 14300
rect 7742 14260 7748 14272
rect 7703 14232 7748 14260
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 8018 14056 8024 14068
rect 7979 14028 8024 14056
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 8260 14028 9413 14056
rect 8260 14016 8266 14028
rect 9401 14025 9413 14028
rect 9447 14025 9459 14059
rect 9401 14019 9459 14025
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 8573 13923 8631 13929
rect 8573 13920 8585 13923
rect 8352 13892 8585 13920
rect 8352 13880 8358 13892
rect 8573 13889 8585 13892
rect 8619 13920 8631 13923
rect 9033 13923 9091 13929
rect 9033 13920 9045 13923
rect 8619 13892 9045 13920
rect 8619 13889 8631 13892
rect 8573 13883 8631 13889
rect 9033 13889 9045 13892
rect 9079 13889 9091 13923
rect 9033 13883 9091 13889
rect 7834 13852 7840 13864
rect 7795 13824 7840 13852
rect 7834 13812 7840 13824
rect 7892 13852 7898 13864
rect 8478 13852 8484 13864
rect 7892 13824 8484 13852
rect 7892 13812 7898 13824
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 7009 13787 7067 13793
rect 7009 13753 7021 13787
rect 7055 13784 7067 13787
rect 7561 13787 7619 13793
rect 7561 13784 7573 13787
rect 7055 13756 7573 13784
rect 7055 13753 7067 13756
rect 7009 13747 7067 13753
rect 7561 13753 7573 13756
rect 7607 13784 7619 13787
rect 8389 13787 8447 13793
rect 8389 13784 8401 13787
rect 7607 13756 8401 13784
rect 7607 13753 7619 13756
rect 7561 13747 7619 13753
rect 8389 13753 8401 13756
rect 8435 13753 8447 13787
rect 8389 13747 8447 13753
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 7101 13515 7159 13521
rect 7101 13481 7113 13515
rect 7147 13512 7159 13515
rect 7374 13512 7380 13524
rect 7147 13484 7380 13512
rect 7147 13481 7159 13484
rect 7101 13475 7159 13481
rect 7374 13472 7380 13484
rect 7432 13512 7438 13524
rect 7742 13512 7748 13524
rect 7432 13484 7748 13512
rect 7432 13472 7438 13484
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 7837 13515 7895 13521
rect 7837 13481 7849 13515
rect 7883 13512 7895 13515
rect 7926 13512 7932 13524
rect 7883 13484 7932 13512
rect 7883 13481 7895 13484
rect 7837 13475 7895 13481
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 8021 13515 8079 13521
rect 8021 13481 8033 13515
rect 8067 13512 8079 13515
rect 8202 13512 8208 13524
rect 8067 13484 8208 13512
rect 8067 13481 8079 13484
rect 8021 13475 8079 13481
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 8754 13512 8760 13524
rect 8527 13484 8760 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 7944 13444 7972 13472
rect 8570 13444 8576 13456
rect 7944 13416 8576 13444
rect 8570 13404 8576 13416
rect 8628 13404 8634 13456
rect 11330 13444 11336 13456
rect 10796 13416 11336 13444
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1670 13376 1676 13388
rect 1443 13348 1676 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1670 13336 1676 13348
rect 1728 13376 1734 13388
rect 2682 13376 2688 13388
rect 1728 13348 2688 13376
rect 1728 13336 1734 13348
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 8110 13376 8116 13388
rect 7708 13348 8116 13376
rect 7708 13336 7714 13348
rect 8110 13336 8116 13348
rect 8168 13376 8174 13388
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 8168 13348 8401 13376
rect 8168 13336 8174 13348
rect 8389 13345 8401 13348
rect 8435 13376 8447 13379
rect 9490 13376 9496 13388
rect 8435 13348 9496 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 10134 13336 10140 13388
rect 10192 13376 10198 13388
rect 10796 13385 10824 13416
rect 11330 13404 11336 13416
rect 11388 13404 11394 13456
rect 11054 13385 11060 13388
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 10192 13348 10241 13376
rect 10192 13336 10198 13348
rect 10229 13345 10241 13348
rect 10275 13376 10287 13379
rect 10781 13379 10839 13385
rect 10781 13376 10793 13379
rect 10275 13348 10793 13376
rect 10275 13345 10287 13348
rect 10229 13339 10287 13345
rect 10781 13345 10793 13348
rect 10827 13345 10839 13379
rect 11048 13376 11060 13385
rect 11015 13348 11060 13376
rect 10781 13339 10839 13345
rect 11048 13339 11060 13348
rect 11054 13336 11060 13339
rect 11112 13336 11118 13388
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 13245 13379 13303 13385
rect 13245 13376 13257 13379
rect 12216 13348 13257 13376
rect 12216 13336 12222 13348
rect 13245 13345 13257 13348
rect 13291 13345 13303 13379
rect 13245 13339 13303 13345
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13308 2375 13311
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 2363 13280 2513 13308
rect 2363 13277 2375 13280
rect 2317 13271 2375 13277
rect 2501 13277 2513 13280
rect 2547 13308 2559 13311
rect 2590 13308 2596 13320
rect 2547 13280 2596 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2590 13268 2596 13280
rect 2648 13268 2654 13320
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 8294 13200 8300 13252
rect 8352 13240 8358 13252
rect 8588 13240 8616 13271
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 12989 13311 13047 13317
rect 12989 13308 13001 13311
rect 12952 13280 13001 13308
rect 12952 13268 12958 13280
rect 12989 13277 13001 13280
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 8352 13212 8616 13240
rect 8352 13200 8358 13212
rect 1394 13132 1400 13184
rect 1452 13172 1458 13184
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 1452 13144 1593 13172
rect 1452 13132 1458 13144
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 9122 13172 9128 13184
rect 9083 13144 9128 13172
rect 1581 13135 1639 13141
rect 9122 13132 9128 13144
rect 9180 13132 9186 13184
rect 12158 13172 12164 13184
rect 12119 13144 12164 13172
rect 12158 13132 12164 13144
rect 12216 13132 12222 13184
rect 14369 13175 14427 13181
rect 14369 13141 14381 13175
rect 14415 13172 14427 13175
rect 15102 13172 15108 13184
rect 14415 13144 15108 13172
rect 14415 13141 14427 13144
rect 14369 13135 14427 13141
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 15286 13132 15292 13184
rect 15344 13172 15350 13184
rect 15473 13175 15531 13181
rect 15473 13172 15485 13175
rect 15344 13144 15485 13172
rect 15344 13132 15350 13144
rect 15473 13141 15485 13144
rect 15519 13141 15531 13175
rect 15473 13135 15531 13141
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 1670 12968 1676 12980
rect 1631 12940 1676 12968
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 8110 12968 8116 12980
rect 8071 12940 8116 12968
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 8481 12971 8539 12977
rect 8481 12937 8493 12971
rect 8527 12968 8539 12971
rect 8754 12968 8760 12980
rect 8527 12940 8760 12968
rect 8527 12937 8539 12940
rect 8481 12931 8539 12937
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12713 12971 12771 12977
rect 12713 12968 12725 12971
rect 12216 12940 12725 12968
rect 12216 12928 12222 12940
rect 12713 12937 12725 12940
rect 12759 12937 12771 12971
rect 15102 12968 15108 12980
rect 15063 12940 15108 12968
rect 12713 12931 12771 12937
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 8573 12903 8631 12909
rect 8573 12900 8585 12903
rect 7484 12872 8585 12900
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 2915 12804 3249 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 3237 12801 3249 12804
rect 3283 12832 3295 12835
rect 3510 12832 3516 12844
rect 3283 12804 3516 12832
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 3510 12792 3516 12804
rect 3568 12832 3574 12844
rect 3881 12835 3939 12841
rect 3881 12832 3893 12835
rect 3568 12804 3893 12832
rect 3568 12792 3574 12804
rect 3881 12801 3893 12804
rect 3927 12832 3939 12835
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 3927 12804 3985 12832
rect 3927 12801 3939 12804
rect 3881 12795 3939 12801
rect 3973 12801 3985 12804
rect 4019 12801 4031 12835
rect 3973 12795 4031 12801
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7484 12841 7512 12872
rect 8573 12869 8585 12872
rect 8619 12869 8631 12903
rect 8573 12863 8631 12869
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 7156 12804 7481 12832
rect 7156 12792 7162 12804
rect 7469 12801 7481 12804
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 9125 12835 9183 12841
rect 9125 12832 9137 12835
rect 7616 12804 7709 12832
rect 8588 12804 9137 12832
rect 7616 12792 7622 12804
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3697 12767 3755 12773
rect 3697 12733 3709 12767
rect 3743 12764 3755 12767
rect 4154 12764 4160 12776
rect 3743 12736 4160 12764
rect 3743 12733 3755 12736
rect 3697 12727 3755 12733
rect 4154 12724 4160 12736
rect 4212 12724 4218 12776
rect 7374 12764 7380 12776
rect 7335 12736 7380 12764
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 2130 12696 2136 12708
rect 2043 12668 2136 12696
rect 2130 12656 2136 12668
rect 2188 12696 2194 12708
rect 2682 12696 2688 12708
rect 2188 12668 2688 12696
rect 2188 12656 2194 12668
rect 2682 12656 2688 12668
rect 2740 12656 2746 12708
rect 3881 12699 3939 12705
rect 3881 12665 3893 12699
rect 3927 12696 3939 12699
rect 4402 12699 4460 12705
rect 4402 12696 4414 12699
rect 3927 12668 4414 12696
rect 3927 12665 3939 12668
rect 3881 12659 3939 12665
rect 4402 12665 4414 12668
rect 4448 12665 4460 12699
rect 4402 12659 4460 12665
rect 6641 12699 6699 12705
rect 6641 12665 6653 12699
rect 6687 12696 6699 12699
rect 7576 12696 7604 12792
rect 8588 12776 8616 12804
rect 9125 12801 9137 12804
rect 9171 12801 9183 12835
rect 10134 12832 10140 12844
rect 10095 12804 10140 12832
rect 9125 12795 9183 12801
rect 10134 12792 10140 12804
rect 10192 12792 10198 12844
rect 13541 12835 13599 12841
rect 13541 12801 13553 12835
rect 13587 12832 13599 12835
rect 14090 12832 14096 12844
rect 13587 12804 14096 12832
rect 13587 12801 13599 12804
rect 13541 12795 13599 12801
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12832 14335 12835
rect 14458 12832 14464 12844
rect 14323 12804 14464 12832
rect 14323 12801 14335 12804
rect 14277 12795 14335 12801
rect 14458 12792 14464 12804
rect 14516 12832 14522 12844
rect 14645 12835 14703 12841
rect 14645 12832 14657 12835
rect 14516 12804 14657 12832
rect 14516 12792 14522 12804
rect 14645 12801 14657 12804
rect 14691 12801 14703 12835
rect 15286 12832 15292 12844
rect 15247 12804 15292 12832
rect 14645 12795 14703 12801
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 8570 12724 8576 12776
rect 8628 12724 8634 12776
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15545 12767 15603 12773
rect 15545 12764 15557 12767
rect 15252 12736 15557 12764
rect 15252 12724 15258 12736
rect 15545 12733 15557 12736
rect 15591 12764 15603 12767
rect 16390 12764 16396 12776
rect 15591 12736 16396 12764
rect 15591 12733 15603 12736
rect 15545 12727 15603 12733
rect 16390 12724 16396 12736
rect 16448 12724 16454 12776
rect 6687 12668 7604 12696
rect 8941 12699 8999 12705
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 8941 12665 8953 12699
rect 8987 12696 8999 12699
rect 9122 12696 9128 12708
rect 8987 12668 9128 12696
rect 8987 12665 8999 12668
rect 8941 12659 8999 12665
rect 9122 12656 9128 12668
rect 9180 12696 9186 12708
rect 9582 12696 9588 12708
rect 9180 12668 9588 12696
rect 9180 12656 9186 12668
rect 9582 12656 9588 12668
rect 9640 12656 9646 12708
rect 10045 12699 10103 12705
rect 10045 12665 10057 12699
rect 10091 12696 10103 12699
rect 10318 12696 10324 12708
rect 10091 12668 10324 12696
rect 10091 12665 10103 12668
rect 10045 12659 10103 12665
rect 10318 12656 10324 12668
rect 10376 12705 10382 12708
rect 10376 12699 10440 12705
rect 10376 12665 10394 12699
rect 10428 12665 10440 12699
rect 10376 12659 10440 12665
rect 10376 12656 10382 12659
rect 11054 12656 11060 12708
rect 11112 12656 11118 12708
rect 13173 12699 13231 12705
rect 13173 12665 13185 12699
rect 13219 12696 13231 12699
rect 13219 12668 14044 12696
rect 13219 12665 13231 12668
rect 13173 12659 13231 12665
rect 2222 12628 2228 12640
rect 2183 12600 2228 12628
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 5534 12628 5540 12640
rect 5495 12600 5540 12628
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 7009 12631 7067 12637
rect 7009 12597 7021 12631
rect 7055 12628 7067 12631
rect 7190 12628 7196 12640
rect 7055 12600 7196 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 9030 12628 9036 12640
rect 8991 12600 9036 12628
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 10870 12588 10876 12640
rect 10928 12628 10934 12640
rect 11072 12628 11100 12656
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 10928 12600 11529 12628
rect 10928 12588 10934 12600
rect 11517 12597 11529 12600
rect 11563 12597 11575 12631
rect 13630 12628 13636 12640
rect 13591 12600 13636 12628
rect 11517 12591 11575 12597
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 14016 12637 14044 12668
rect 14001 12631 14059 12637
rect 14001 12597 14013 12631
rect 14047 12628 14059 12631
rect 15194 12628 15200 12640
rect 14047 12600 15200 12628
rect 14047 12597 14059 12600
rect 14001 12591 14059 12597
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 16666 12628 16672 12640
rect 16627 12600 16672 12628
rect 16666 12588 16672 12600
rect 16724 12588 16730 12640
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 2774 12424 2780 12436
rect 2687 12396 2780 12424
rect 2774 12384 2780 12396
rect 2832 12424 2838 12436
rect 6270 12424 6276 12436
rect 2832 12396 6276 12424
rect 2832 12384 2838 12396
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 7098 12424 7104 12436
rect 7059 12396 7104 12424
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 8113 12427 8171 12433
rect 8113 12393 8125 12427
rect 8159 12424 8171 12427
rect 8294 12424 8300 12436
rect 8159 12396 8300 12424
rect 8159 12393 8171 12396
rect 8113 12387 8171 12393
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 8665 12427 8723 12433
rect 8665 12424 8677 12427
rect 8628 12396 8677 12424
rect 8628 12384 8634 12396
rect 8665 12393 8677 12396
rect 8711 12424 8723 12427
rect 10870 12424 10876 12436
rect 8711 12396 10876 12424
rect 8711 12393 8723 12396
rect 8665 12387 8723 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 11330 12424 11336 12436
rect 11287 12396 11336 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 15252 12396 15301 12424
rect 15252 12384 15258 12396
rect 15289 12393 15301 12396
rect 15335 12393 15347 12427
rect 15289 12387 15347 12393
rect 16390 12384 16396 12436
rect 16448 12424 16454 12436
rect 17221 12427 17279 12433
rect 17221 12424 17233 12427
rect 16448 12396 17233 12424
rect 16448 12384 16454 12396
rect 17221 12393 17233 12396
rect 17267 12393 17279 12427
rect 17221 12387 17279 12393
rect 4890 12316 4896 12368
rect 4948 12356 4954 12368
rect 5138 12359 5196 12365
rect 5138 12356 5150 12359
rect 4948 12328 5150 12356
rect 4948 12316 4954 12328
rect 5138 12325 5150 12328
rect 5184 12356 5196 12359
rect 5534 12356 5540 12368
rect 5184 12328 5540 12356
rect 5184 12325 5196 12328
rect 5138 12319 5196 12325
rect 5534 12316 5540 12328
rect 5592 12316 5598 12368
rect 8312 12356 8340 12384
rect 8312 12328 10180 12356
rect 2685 12291 2743 12297
rect 2685 12257 2697 12291
rect 2731 12288 2743 12291
rect 2866 12288 2872 12300
rect 2731 12260 2872 12288
rect 2731 12257 2743 12260
rect 2685 12251 2743 12257
rect 2866 12248 2872 12260
rect 2924 12288 2930 12300
rect 3050 12288 3056 12300
rect 2924 12260 3056 12288
rect 2924 12248 2930 12260
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 10152 12288 10180 12328
rect 13446 12316 13452 12368
rect 13504 12356 13510 12368
rect 14001 12359 14059 12365
rect 14001 12356 14013 12359
rect 13504 12328 14013 12356
rect 13504 12316 13510 12328
rect 14001 12325 14013 12328
rect 14047 12325 14059 12359
rect 17236 12356 17264 12387
rect 17236 12328 17908 12356
rect 14001 12319 14059 12325
rect 10318 12288 10324 12300
rect 10152 12260 10324 12288
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3510 12220 3516 12232
rect 3007 12192 3516 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 3510 12180 3516 12192
rect 3568 12180 3574 12232
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 4706 12220 4712 12232
rect 4212 12192 4712 12220
rect 4212 12180 4218 12192
rect 4706 12180 4712 12192
rect 4764 12220 4770 12232
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4764 12192 4905 12220
rect 4764 12180 4770 12192
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 10134 12220 10140 12232
rect 10095 12192 10140 12220
rect 4893 12183 4951 12189
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10244 12229 10272 12260
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 16758 12248 16764 12300
rect 16816 12288 16822 12300
rect 17678 12288 17684 12300
rect 16816 12260 17684 12288
rect 16816 12248 16822 12260
rect 17678 12248 17684 12260
rect 17736 12288 17742 12300
rect 17773 12291 17831 12297
rect 17773 12288 17785 12291
rect 17736 12260 17785 12288
rect 17736 12248 17742 12260
rect 17773 12257 17785 12260
rect 17819 12257 17831 12291
rect 17880 12288 17908 12328
rect 17880 12260 18000 12288
rect 17773 12251 17831 12257
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 13170 12180 13176 12232
rect 13228 12220 13234 12232
rect 14090 12220 14096 12232
rect 13228 12192 14096 12220
rect 13228 12180 13234 12192
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 14458 12220 14464 12232
rect 14323 12192 14464 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 17494 12180 17500 12232
rect 17552 12220 17558 12232
rect 17972 12229 18000 12260
rect 17865 12223 17923 12229
rect 17865 12220 17877 12223
rect 17552 12192 17877 12220
rect 17552 12180 17558 12192
rect 17865 12189 17877 12192
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18417 12223 18475 12229
rect 18417 12220 18429 12223
rect 18003 12192 18429 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18417 12189 18429 12192
rect 18463 12220 18475 12223
rect 18598 12220 18604 12232
rect 18463 12192 18604 12220
rect 18463 12189 18475 12192
rect 18417 12183 18475 12189
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 9030 12152 9036 12164
rect 8943 12124 9036 12152
rect 9030 12112 9036 12124
rect 9088 12152 9094 12164
rect 9677 12155 9735 12161
rect 9677 12152 9689 12155
rect 9088 12124 9689 12152
rect 9088 12112 9094 12124
rect 9677 12121 9689 12124
rect 9723 12121 9735 12155
rect 9677 12115 9735 12121
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12084 2099 12087
rect 2317 12087 2375 12093
rect 2317 12084 2329 12087
rect 2087 12056 2329 12084
rect 2087 12053 2099 12056
rect 2041 12047 2099 12053
rect 2317 12053 2329 12056
rect 2363 12084 2375 12087
rect 2406 12084 2412 12096
rect 2363 12056 2412 12084
rect 2363 12053 2375 12056
rect 2317 12047 2375 12053
rect 2406 12044 2412 12056
rect 2464 12044 2470 12096
rect 6270 12084 6276 12096
rect 6231 12056 6276 12084
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 12894 12084 12900 12096
rect 11388 12056 12900 12084
rect 11388 12044 11394 12056
rect 12894 12044 12900 12056
rect 12952 12084 12958 12096
rect 13081 12087 13139 12093
rect 13081 12084 13093 12087
rect 12952 12056 13093 12084
rect 12952 12044 12958 12056
rect 13081 12053 13093 12056
rect 13127 12084 13139 12087
rect 13538 12084 13544 12096
rect 13127 12056 13544 12084
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 13633 12087 13691 12093
rect 13633 12053 13645 12087
rect 13679 12084 13691 12087
rect 13722 12084 13728 12096
rect 13679 12056 13728 12084
rect 13679 12053 13691 12056
rect 13633 12047 13691 12053
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 16485 12087 16543 12093
rect 16485 12053 16497 12087
rect 16531 12084 16543 12087
rect 16850 12084 16856 12096
rect 16531 12056 16856 12084
rect 16531 12053 16543 12056
rect 16485 12047 16543 12053
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 17402 12084 17408 12096
rect 17363 12056 17408 12084
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 1857 11883 1915 11889
rect 1857 11849 1869 11883
rect 1903 11880 1915 11883
rect 2038 11880 2044 11892
rect 1903 11852 2044 11880
rect 1903 11849 1915 11852
rect 1857 11843 1915 11849
rect 2038 11840 2044 11852
rect 2096 11880 2102 11892
rect 2774 11880 2780 11892
rect 2096 11852 2780 11880
rect 2096 11840 2102 11852
rect 2774 11840 2780 11852
rect 2832 11840 2838 11892
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 4764 11852 5273 11880
rect 4764 11840 4770 11852
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 4890 11812 4896 11824
rect 4851 11784 4896 11812
rect 4890 11772 4896 11784
rect 4948 11772 4954 11824
rect 2406 11744 2412 11756
rect 2367 11716 2412 11744
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 2590 11744 2596 11756
rect 2551 11716 2596 11744
rect 2590 11704 2596 11716
rect 2648 11704 2654 11756
rect 5276 11744 5304 11843
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 11149 11883 11207 11889
rect 11149 11880 11161 11883
rect 10192 11852 11161 11880
rect 10192 11840 10198 11852
rect 11149 11849 11161 11852
rect 11195 11849 11207 11883
rect 13170 11880 13176 11892
rect 13131 11852 13176 11880
rect 11149 11843 11207 11849
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 13446 11880 13452 11892
rect 13407 11852 13452 11880
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 15286 11880 15292 11892
rect 13596 11852 15292 11880
rect 13596 11840 13602 11852
rect 10410 11772 10416 11824
rect 10468 11812 10474 11824
rect 10781 11815 10839 11821
rect 10781 11812 10793 11815
rect 10468 11784 10793 11812
rect 10468 11772 10474 11784
rect 10781 11781 10793 11784
rect 10827 11781 10839 11815
rect 10781 11775 10839 11781
rect 6822 11744 6828 11756
rect 5276 11716 6828 11744
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 10318 11744 10324 11756
rect 8864 11716 10324 11744
rect 2222 11636 2228 11688
rect 2280 11676 2286 11688
rect 2317 11679 2375 11685
rect 2317 11676 2329 11679
rect 2280 11648 2329 11676
rect 2280 11636 2286 11648
rect 2317 11645 2329 11648
rect 2363 11676 2375 11679
rect 3697 11679 3755 11685
rect 3697 11676 3709 11679
rect 2363 11648 3709 11676
rect 2363 11645 2375 11648
rect 2317 11639 2375 11645
rect 3697 11645 3709 11648
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 4614 11568 4620 11620
rect 4672 11608 4678 11620
rect 6270 11608 6276 11620
rect 4672 11580 6276 11608
rect 4672 11568 4678 11580
rect 6270 11568 6276 11580
rect 6328 11608 6334 11620
rect 6549 11611 6607 11617
rect 6549 11608 6561 11611
rect 6328 11580 6561 11608
rect 6328 11568 6334 11580
rect 6549 11577 6561 11580
rect 6595 11608 6607 11611
rect 7070 11611 7128 11617
rect 7070 11608 7082 11611
rect 6595 11580 7082 11608
rect 6595 11577 6607 11580
rect 6549 11571 6607 11577
rect 7070 11577 7082 11580
rect 7116 11577 7128 11611
rect 7070 11571 7128 11577
rect 1946 11540 1952 11552
rect 1907 11512 1952 11540
rect 1946 11500 1952 11512
rect 2004 11500 2010 11552
rect 3050 11540 3056 11552
rect 3011 11512 3056 11540
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 3421 11543 3479 11549
rect 3421 11509 3433 11543
rect 3467 11540 3479 11543
rect 3510 11540 3516 11552
rect 3467 11512 3516 11540
rect 3467 11509 3479 11512
rect 3421 11503 3479 11509
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 8864 11549 8892 11716
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 13648 11753 13676 11852
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 16301 11883 16359 11889
rect 16301 11849 16313 11883
rect 16347 11880 16359 11883
rect 16666 11880 16672 11892
rect 16347 11852 16672 11880
rect 16347 11849 16359 11852
rect 16301 11843 16359 11849
rect 16666 11840 16672 11852
rect 16724 11880 16730 11892
rect 16942 11880 16948 11892
rect 16724 11852 16948 11880
rect 16724 11840 16730 11852
rect 16942 11840 16948 11852
rect 17000 11840 17006 11892
rect 17678 11840 17684 11892
rect 17736 11880 17742 11892
rect 19058 11880 19064 11892
rect 17736 11852 19064 11880
rect 17736 11840 17742 11852
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11713 13691 11747
rect 16942 11744 16948 11756
rect 16903 11716 16948 11744
rect 13633 11707 13691 11713
rect 16942 11704 16948 11716
rect 17000 11704 17006 11756
rect 17678 11704 17684 11756
rect 17736 11744 17742 11756
rect 17773 11747 17831 11753
rect 17773 11744 17785 11747
rect 17736 11716 17785 11744
rect 17736 11704 17742 11716
rect 17773 11713 17785 11716
rect 17819 11713 17831 11747
rect 18598 11744 18604 11756
rect 18559 11716 18604 11744
rect 17773 11707 17831 11713
rect 10137 11679 10195 11685
rect 10137 11676 10149 11679
rect 9232 11648 10149 11676
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 7524 11512 8217 11540
rect 7524 11500 7530 11512
rect 8205 11509 8217 11512
rect 8251 11540 8263 11543
rect 8849 11543 8907 11549
rect 8849 11540 8861 11543
rect 8251 11512 8861 11540
rect 8251 11509 8263 11512
rect 8205 11503 8263 11509
rect 8849 11509 8861 11512
rect 8895 11509 8907 11543
rect 8849 11503 8907 11509
rect 9122 11500 9128 11552
rect 9180 11540 9186 11552
rect 9232 11549 9260 11648
rect 10137 11645 10149 11648
rect 10183 11676 10195 11679
rect 10226 11676 10232 11688
rect 10183 11648 10232 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11676 15991 11679
rect 16761 11679 16819 11685
rect 16761 11676 16773 11679
rect 15979 11648 16773 11676
rect 15979 11645 15991 11648
rect 15933 11639 15991 11645
rect 16761 11645 16773 11648
rect 16807 11676 16819 11679
rect 17402 11676 17408 11688
rect 16807 11648 17408 11676
rect 16807 11645 16819 11648
rect 16761 11639 16819 11645
rect 17402 11636 17408 11648
rect 17460 11636 17466 11688
rect 17788 11676 17816 11707
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 17788 11648 18521 11676
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 26418 11676 26424 11688
rect 26379 11648 26424 11676
rect 18509 11639 18567 11645
rect 26418 11636 26424 11648
rect 26476 11676 26482 11688
rect 26973 11679 27031 11685
rect 26973 11676 26985 11679
rect 26476 11648 26985 11676
rect 26476 11636 26482 11648
rect 26973 11645 26985 11648
rect 27019 11645 27031 11679
rect 26973 11639 27031 11645
rect 9674 11608 9680 11620
rect 9587 11580 9680 11608
rect 9674 11568 9680 11580
rect 9732 11608 9738 11620
rect 12805 11611 12863 11617
rect 9732 11580 10272 11608
rect 9732 11568 9738 11580
rect 10244 11552 10272 11580
rect 12805 11577 12817 11611
rect 12851 11608 12863 11611
rect 13900 11611 13958 11617
rect 13900 11608 13912 11611
rect 12851 11580 13912 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 13900 11577 13912 11580
rect 13946 11608 13958 11611
rect 14458 11608 14464 11620
rect 13946 11580 14464 11608
rect 13946 11577 13958 11580
rect 13900 11571 13958 11577
rect 14458 11568 14464 11580
rect 14516 11568 14522 11620
rect 16850 11608 16856 11620
rect 16811 11580 16856 11608
rect 16850 11568 16856 11580
rect 16908 11608 16914 11620
rect 16908 11580 18092 11608
rect 16908 11568 16914 11580
rect 9217 11543 9275 11549
rect 9217 11540 9229 11543
rect 9180 11512 9229 11540
rect 9180 11500 9186 11512
rect 9217 11509 9229 11512
rect 9263 11509 9275 11543
rect 9766 11540 9772 11552
rect 9727 11512 9772 11540
rect 9217 11503 9275 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 15013 11543 15071 11549
rect 10284 11512 10329 11540
rect 10284 11500 10290 11512
rect 15013 11509 15025 11543
rect 15059 11540 15071 11543
rect 15102 11540 15108 11552
rect 15059 11512 15108 11540
rect 15059 11509 15071 11512
rect 15013 11503 15071 11509
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 15654 11540 15660 11552
rect 15344 11512 15660 11540
rect 15344 11500 15350 11512
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 16390 11540 16396 11552
rect 16351 11512 16396 11540
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 17402 11540 17408 11552
rect 17363 11512 17408 11540
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 18064 11549 18092 11580
rect 18049 11543 18107 11549
rect 18049 11509 18061 11543
rect 18095 11509 18107 11543
rect 18414 11540 18420 11552
rect 18375 11512 18420 11540
rect 18049 11503 18107 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 26602 11540 26608 11552
rect 26563 11512 26608 11540
rect 26602 11500 26608 11512
rect 26660 11500 26666 11552
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 4430 11336 4436 11348
rect 2179 11308 4436 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 4430 11296 4436 11308
rect 4488 11336 4494 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4488 11308 4537 11336
rect 4488 11296 4494 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 6822 11336 6828 11348
rect 6783 11308 6828 11336
rect 4525 11299 4583 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 8294 11296 8300 11348
rect 8352 11336 8358 11348
rect 8757 11339 8815 11345
rect 8757 11336 8769 11339
rect 8352 11308 8769 11336
rect 8352 11296 8358 11308
rect 8757 11305 8769 11308
rect 8803 11305 8815 11339
rect 8757 11299 8815 11305
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 10042 11336 10048 11348
rect 9539 11308 10048 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10137 11339 10195 11345
rect 10137 11305 10149 11339
rect 10183 11336 10195 11339
rect 10778 11336 10784 11348
rect 10183 11308 10784 11336
rect 10183 11305 10195 11308
rect 10137 11299 10195 11305
rect 2041 11271 2099 11277
rect 2041 11237 2053 11271
rect 2087 11268 2099 11271
rect 2590 11268 2596 11280
rect 2087 11240 2596 11268
rect 2087 11237 2099 11240
rect 2041 11231 2099 11237
rect 2590 11228 2596 11240
rect 2648 11228 2654 11280
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11200 1731 11203
rect 2314 11200 2320 11212
rect 1719 11172 2320 11200
rect 1719 11169 1731 11172
rect 1673 11163 1731 11169
rect 2314 11160 2320 11172
rect 2372 11200 2378 11212
rect 2501 11203 2559 11209
rect 2501 11200 2513 11203
rect 2372 11172 2513 11200
rect 2372 11160 2378 11172
rect 2501 11169 2513 11172
rect 2547 11169 2559 11203
rect 2608 11200 2636 11228
rect 2608 11172 2728 11200
rect 2501 11163 2559 11169
rect 2700 11141 2728 11172
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4396 11172 4445 11200
rect 4396 11160 4402 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 6840 11200 6868 11296
rect 9950 11228 9956 11280
rect 10008 11268 10014 11280
rect 10502 11268 10508 11280
rect 10008 11240 10508 11268
rect 10008 11228 10014 11240
rect 10502 11228 10508 11240
rect 10560 11228 10566 11280
rect 7374 11200 7380 11212
rect 6840 11172 7380 11200
rect 4433 11163 4491 11169
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 7633 11203 7691 11209
rect 7633 11200 7645 11203
rect 7524 11172 7645 11200
rect 7524 11160 7530 11172
rect 7633 11169 7645 11172
rect 7679 11169 7691 11203
rect 10612 11200 10640 11308
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 13630 11336 13636 11348
rect 13311 11308 13636 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 13630 11296 13636 11308
rect 13688 11336 13694 11348
rect 13725 11339 13783 11345
rect 13725 11336 13737 11339
rect 13688 11308 13737 11336
rect 13688 11296 13694 11308
rect 13725 11305 13737 11308
rect 13771 11305 13783 11339
rect 13725 11299 13783 11305
rect 16209 11339 16267 11345
rect 16209 11305 16221 11339
rect 16255 11336 16267 11339
rect 16298 11336 16304 11348
rect 16255 11308 16304 11336
rect 16255 11305 16267 11308
rect 16209 11299 16267 11305
rect 16298 11296 16304 11308
rect 16356 11336 16362 11348
rect 17313 11339 17371 11345
rect 17313 11336 17325 11339
rect 16356 11308 17325 11336
rect 16356 11296 16362 11308
rect 17313 11305 17325 11308
rect 17359 11305 17371 11339
rect 17313 11299 17371 11305
rect 15470 11228 15476 11280
rect 15528 11268 15534 11280
rect 15654 11268 15660 11280
rect 15528 11240 15660 11268
rect 15528 11228 15534 11240
rect 15654 11228 15660 11240
rect 15712 11268 15718 11280
rect 16117 11271 16175 11277
rect 16117 11268 16129 11271
rect 15712 11240 16129 11268
rect 15712 11228 15718 11240
rect 16117 11237 16129 11240
rect 16163 11237 16175 11271
rect 16117 11231 16175 11237
rect 17954 11228 17960 11280
rect 18012 11268 18018 11280
rect 18325 11271 18383 11277
rect 18325 11268 18337 11271
rect 18012 11240 18337 11268
rect 18012 11228 18018 11240
rect 18325 11237 18337 11240
rect 18371 11268 18383 11271
rect 18414 11268 18420 11280
rect 18371 11240 18420 11268
rect 18371 11237 18383 11240
rect 18325 11231 18383 11237
rect 18414 11228 18420 11240
rect 18472 11228 18478 11280
rect 7633 11163 7691 11169
rect 9600 11172 10640 11200
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11101 2651 11135
rect 2593 11095 2651 11101
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11101 2743 11135
rect 4614 11132 4620 11144
rect 4575 11104 4620 11132
rect 2685 11095 2743 11101
rect 2608 10996 2636 11095
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 4065 11067 4123 11073
rect 4065 11064 4077 11067
rect 2832 11036 4077 11064
rect 2832 11024 2838 11036
rect 4065 11033 4077 11036
rect 4111 11033 4123 11067
rect 4065 11027 4123 11033
rect 2866 10996 2872 11008
rect 2608 10968 2872 10996
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 3237 10999 3295 11005
rect 3237 10965 3249 10999
rect 3283 10996 3295 10999
rect 3326 10996 3332 11008
rect 3283 10968 3332 10996
rect 3283 10965 3295 10968
rect 3237 10959 3295 10965
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 8938 10956 8944 11008
rect 8996 10996 9002 11008
rect 9398 10996 9404 11008
rect 8996 10968 9404 10996
rect 8996 10956 9002 10968
rect 9398 10956 9404 10968
rect 9456 10996 9462 11008
rect 9600 10996 9628 11172
rect 13722 11160 13728 11212
rect 13780 11200 13786 11212
rect 13817 11203 13875 11209
rect 13817 11200 13829 11203
rect 13780 11172 13829 11200
rect 13780 11160 13786 11172
rect 13817 11169 13829 11172
rect 13863 11169 13875 11203
rect 14458 11200 14464 11212
rect 14371 11172 14464 11200
rect 13817 11163 13875 11169
rect 14458 11160 14464 11172
rect 14516 11200 14522 11212
rect 17678 11200 17684 11212
rect 14516 11172 15884 11200
rect 17639 11172 17684 11200
rect 14516 11160 14522 11172
rect 15856 11144 15884 11172
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 21910 11160 21916 11212
rect 21968 11200 21974 11212
rect 26513 11203 26571 11209
rect 26513 11200 26525 11203
rect 21968 11172 26525 11200
rect 21968 11160 21974 11172
rect 26513 11169 26525 11172
rect 26559 11200 26571 11203
rect 27338 11200 27344 11212
rect 26559 11172 27344 11200
rect 26559 11169 26571 11172
rect 26513 11163 26571 11169
rect 27338 11160 27344 11172
rect 27396 11160 27402 11212
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 9732 11104 10241 11132
rect 9732 11092 9738 11104
rect 10229 11101 10241 11104
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 9769 11067 9827 11073
rect 9769 11033 9781 11067
rect 9815 11064 9827 11067
rect 10134 11064 10140 11076
rect 9815 11036 10140 11064
rect 9815 11033 9827 11036
rect 9769 11027 9827 11033
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 10244 11064 10272 11095
rect 10318 11092 10324 11144
rect 10376 11132 10382 11144
rect 10376 11104 10421 11132
rect 10376 11092 10382 11104
rect 13078 11092 13084 11144
rect 13136 11132 13142 11144
rect 13909 11135 13967 11141
rect 13909 11132 13921 11135
rect 13136 11104 13921 11132
rect 13136 11092 13142 11104
rect 13909 11101 13921 11104
rect 13955 11132 13967 11135
rect 15102 11132 15108 11144
rect 13955 11104 15108 11132
rect 13955 11101 13967 11104
rect 13909 11095 13967 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 16393 11135 16451 11141
rect 16393 11132 16405 11135
rect 15896 11104 16405 11132
rect 15896 11092 15902 11104
rect 16393 11101 16405 11104
rect 16439 11132 16451 11135
rect 16666 11132 16672 11144
rect 16439 11104 16672 11132
rect 16439 11101 16451 11104
rect 16393 11095 16451 11101
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 17494 11092 17500 11144
rect 17552 11132 17558 11144
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 17552 11104 17785 11132
rect 17552 11092 17558 11104
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 17862 11092 17868 11144
rect 17920 11132 17926 11144
rect 17957 11135 18015 11141
rect 17957 11132 17969 11135
rect 17920 11104 17969 11132
rect 17920 11092 17926 11104
rect 17957 11101 17969 11104
rect 18003 11132 18015 11135
rect 18598 11132 18604 11144
rect 18003 11104 18604 11132
rect 18003 11101 18015 11104
rect 17957 11095 18015 11101
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 10502 11064 10508 11076
rect 10244 11036 10508 11064
rect 10502 11024 10508 11036
rect 10560 11024 10566 11076
rect 11514 11024 11520 11076
rect 11572 11064 11578 11076
rect 16574 11064 16580 11076
rect 11572 11036 16580 11064
rect 11572 11024 11578 11036
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 26694 11064 26700 11076
rect 26655 11036 26700 11064
rect 26694 11024 26700 11036
rect 26752 11024 26758 11076
rect 9456 10968 9628 10996
rect 13357 10999 13415 11005
rect 9456 10956 9462 10968
rect 13357 10965 13369 10999
rect 13403 10996 13415 10999
rect 13722 10996 13728 11008
rect 13403 10968 13728 10996
rect 13403 10965 13415 10968
rect 13357 10959 13415 10965
rect 13722 10956 13728 10968
rect 13780 10956 13786 11008
rect 15746 10996 15752 11008
rect 15707 10968 15752 10996
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 2409 10795 2467 10801
rect 2409 10761 2421 10795
rect 2455 10792 2467 10795
rect 2590 10792 2596 10804
rect 2455 10764 2596 10792
rect 2455 10761 2467 10764
rect 2409 10755 2467 10761
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 2866 10792 2872 10804
rect 2827 10764 2872 10792
rect 2866 10752 2872 10764
rect 2924 10752 2930 10804
rect 4157 10795 4215 10801
rect 4157 10761 4169 10795
rect 4203 10792 4215 10795
rect 4614 10792 4620 10804
rect 4203 10764 4620 10792
rect 4203 10761 4215 10764
rect 4157 10755 4215 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 7466 10792 7472 10804
rect 7427 10764 7472 10792
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 8938 10792 8944 10804
rect 8899 10764 8944 10792
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9674 10792 9680 10804
rect 9635 10764 9680 10792
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 9769 10795 9827 10801
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 10042 10792 10048 10804
rect 9815 10764 10048 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 13872 10764 14381 10792
rect 13872 10752 13878 10764
rect 14369 10761 14381 10764
rect 14415 10761 14427 10795
rect 15194 10792 15200 10804
rect 15155 10764 15200 10792
rect 14369 10755 14427 10761
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 17037 10795 17095 10801
rect 17037 10761 17049 10795
rect 17083 10792 17095 10795
rect 17862 10792 17868 10804
rect 17083 10764 17868 10792
rect 17083 10761 17095 10764
rect 17037 10755 17095 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 27338 10792 27344 10804
rect 27299 10764 27344 10792
rect 27338 10752 27344 10764
rect 27396 10752 27402 10804
rect 4430 10724 4436 10736
rect 4391 10696 4436 10724
rect 4430 10684 4436 10696
rect 4488 10684 4494 10736
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 7745 10727 7803 10733
rect 7745 10724 7757 10727
rect 7432 10696 7757 10724
rect 7432 10684 7438 10696
rect 7745 10693 7757 10696
rect 7791 10693 7803 10727
rect 15212 10724 15240 10752
rect 15212 10696 16252 10724
rect 7745 10687 7803 10693
rect 2038 10656 2044 10668
rect 1412 10628 2044 10656
rect 1412 10597 1440 10628
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 3510 10656 3516 10668
rect 2823 10628 3516 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4396 10628 4813 10656
rect 4396 10616 4402 10628
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 10318 10656 10324 10668
rect 10279 10628 10324 10656
rect 4801 10619 4859 10625
rect 10318 10616 10324 10628
rect 10376 10656 10382 10668
rect 11149 10659 11207 10665
rect 11149 10656 11161 10659
rect 10376 10628 11161 10656
rect 10376 10616 10382 10628
rect 11149 10625 11161 10628
rect 11195 10656 11207 10659
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11195 10628 11529 10656
rect 11195 10625 11207 10628
rect 11149 10619 11207 10625
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 13265 10659 13323 10665
rect 13265 10625 13277 10659
rect 13311 10656 13323 10659
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 13311 10628 13921 10656
rect 13311 10625 13323 10628
rect 13265 10619 13323 10625
rect 13909 10625 13921 10628
rect 13955 10656 13967 10659
rect 14366 10656 14372 10668
rect 13955 10628 14372 10656
rect 13955 10625 13967 10628
rect 13909 10619 13967 10625
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 16224 10665 16252 10696
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10656 14887 10659
rect 16209 10659 16267 10665
rect 14875 10628 16160 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10557 1455 10591
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 1397 10551 1455 10557
rect 9232 10560 10241 10588
rect 3237 10523 3295 10529
rect 3237 10489 3249 10523
rect 3283 10520 3295 10523
rect 3418 10520 3424 10532
rect 3283 10492 3424 10520
rect 3283 10489 3295 10492
rect 3237 10483 3295 10489
rect 3418 10480 3424 10492
rect 3476 10480 3482 10532
rect 3326 10452 3332 10464
rect 3287 10424 3332 10452
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 9122 10412 9128 10464
rect 9180 10452 9186 10464
rect 9232 10461 9260 10560
rect 10229 10557 10241 10560
rect 10275 10588 10287 10591
rect 11330 10588 11336 10600
rect 10275 10560 11336 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 11330 10548 11336 10560
rect 11388 10548 11394 10600
rect 15565 10591 15623 10597
rect 15565 10557 15577 10591
rect 15611 10588 15623 10591
rect 15654 10588 15660 10600
rect 15611 10560 15660 10588
rect 15611 10557 15623 10560
rect 15565 10551 15623 10557
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 15746 10548 15752 10600
rect 15804 10588 15810 10600
rect 16132 10597 16160 10628
rect 16209 10625 16221 10659
rect 16255 10625 16267 10659
rect 16209 10619 16267 10625
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15804 10560 16037 10588
rect 15804 10548 15810 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 16390 10588 16396 10600
rect 16163 10560 16396 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 16390 10548 16396 10560
rect 16448 10548 16454 10600
rect 26418 10588 26424 10600
rect 26331 10560 26424 10588
rect 26418 10548 26424 10560
rect 26476 10588 26482 10600
rect 26973 10591 27031 10597
rect 26973 10588 26985 10591
rect 26476 10560 26985 10588
rect 26476 10548 26482 10560
rect 26973 10557 26985 10560
rect 27019 10557 27031 10591
rect 26973 10551 27031 10557
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 10152 10492 10793 10520
rect 10152 10464 10180 10492
rect 10781 10489 10793 10492
rect 10827 10489 10839 10523
rect 10781 10483 10839 10489
rect 13446 10480 13452 10532
rect 13504 10520 13510 10532
rect 13817 10523 13875 10529
rect 13817 10520 13829 10523
rect 13504 10492 13829 10520
rect 13504 10480 13510 10492
rect 13817 10489 13829 10492
rect 13863 10520 13875 10523
rect 13863 10492 15700 10520
rect 13863 10489 13875 10492
rect 13817 10483 13875 10489
rect 9217 10455 9275 10461
rect 9217 10452 9229 10455
rect 9180 10424 9229 10452
rect 9180 10412 9186 10424
rect 9217 10421 9229 10424
rect 9263 10421 9275 10455
rect 10134 10452 10140 10464
rect 10095 10424 10140 10452
rect 9217 10415 9275 10421
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13078 10452 13084 10464
rect 12943 10424 13084 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13078 10412 13084 10424
rect 13136 10412 13142 10464
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 13357 10455 13415 10461
rect 13357 10452 13369 10455
rect 13228 10424 13369 10452
rect 13228 10412 13234 10424
rect 13357 10421 13369 10424
rect 13403 10421 13415 10455
rect 13722 10452 13728 10464
rect 13683 10424 13728 10452
rect 13357 10415 13415 10421
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 15672 10461 15700 10492
rect 15657 10455 15715 10461
rect 15657 10421 15669 10455
rect 15703 10421 15715 10455
rect 15657 10415 15715 10421
rect 17405 10455 17463 10461
rect 17405 10421 17417 10455
rect 17451 10452 17463 10455
rect 17494 10452 17500 10464
rect 17451 10424 17500 10452
rect 17451 10421 17463 10424
rect 17405 10415 17463 10421
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 17678 10452 17684 10464
rect 17639 10424 17684 10452
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 26602 10452 26608 10464
rect 26563 10424 26608 10452
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 6086 10248 6092 10260
rect 6047 10220 6092 10248
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 6880 10220 6929 10248
rect 6880 10208 6886 10220
rect 6917 10217 6929 10220
rect 6963 10248 6975 10251
rect 7374 10248 7380 10260
rect 6963 10220 7380 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7374 10208 7380 10220
rect 7432 10248 7438 10260
rect 7834 10248 7840 10260
rect 7432 10220 7840 10248
rect 7432 10208 7438 10220
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 9674 10248 9680 10260
rect 9635 10220 9680 10248
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 9766 10208 9772 10260
rect 9824 10248 9830 10260
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 9824 10220 10149 10248
rect 9824 10208 9830 10220
rect 10137 10217 10149 10220
rect 10183 10248 10195 10251
rect 10410 10248 10416 10260
rect 10183 10220 10416 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10410 10208 10416 10220
rect 10468 10208 10474 10260
rect 12897 10251 12955 10257
rect 12897 10217 12909 10251
rect 12943 10248 12955 10251
rect 13722 10248 13728 10260
rect 12943 10220 13728 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 14366 10248 14372 10260
rect 14327 10220 14372 10248
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 16485 10251 16543 10257
rect 16485 10248 16497 10251
rect 15804 10220 16497 10248
rect 15804 10208 15810 10220
rect 16485 10217 16497 10220
rect 16531 10217 16543 10251
rect 16485 10211 16543 10217
rect 1857 10183 1915 10189
rect 1857 10149 1869 10183
rect 1903 10180 1915 10183
rect 2866 10180 2872 10192
rect 1903 10152 2872 10180
rect 1903 10149 1915 10152
rect 1857 10143 1915 10149
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 2958 10140 2964 10192
rect 3016 10140 3022 10192
rect 15838 10180 15844 10192
rect 15799 10152 15844 10180
rect 15838 10140 15844 10152
rect 15896 10140 15902 10192
rect 16209 10183 16267 10189
rect 16209 10149 16221 10183
rect 16255 10180 16267 10183
rect 16298 10180 16304 10192
rect 16255 10152 16304 10180
rect 16255 10149 16267 10152
rect 16209 10143 16267 10149
rect 16298 10140 16304 10152
rect 16356 10140 16362 10192
rect 2498 10072 2504 10124
rect 2556 10112 2562 10124
rect 2685 10115 2743 10121
rect 2685 10112 2697 10115
rect 2556 10084 2697 10112
rect 2556 10072 2562 10084
rect 2685 10081 2697 10084
rect 2731 10112 2743 10115
rect 2976 10112 3004 10140
rect 2731 10084 3004 10112
rect 4976 10115 5034 10121
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 4976 10081 4988 10115
rect 5022 10112 5034 10115
rect 5442 10112 5448 10124
rect 5022 10084 5448 10112
rect 5022 10081 5034 10084
rect 4976 10075 5034 10081
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 6972 10084 7113 10112
rect 6972 10072 6978 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 9858 10072 9864 10124
rect 9916 10112 9922 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9916 10084 10057 10112
rect 9916 10072 9922 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 12894 10072 12900 10124
rect 12952 10112 12958 10124
rect 12989 10115 13047 10121
rect 12989 10112 13001 10115
rect 12952 10084 13001 10112
rect 12952 10072 12958 10084
rect 12989 10081 13001 10084
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 13245 10115 13303 10121
rect 13245 10112 13257 10115
rect 13136 10084 13257 10112
rect 13136 10072 13142 10084
rect 13245 10081 13257 10084
rect 13291 10081 13303 10115
rect 13245 10075 13303 10081
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2774 10044 2780 10056
rect 2271 10016 2780 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 2774 10004 2780 10016
rect 2832 10044 2838 10056
rect 2961 10047 3019 10053
rect 2832 10016 2925 10044
rect 2832 10004 2838 10016
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3510 10044 3516 10056
rect 3007 10016 3516 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 2406 9936 2412 9988
rect 2464 9976 2470 9988
rect 2976 9976 3004 10007
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 2464 9948 3004 9976
rect 2464 9936 2470 9948
rect 3418 9908 3424 9920
rect 3379 9880 3424 9908
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 4617 9911 4675 9917
rect 4617 9877 4629 9911
rect 4663 9908 4675 9911
rect 4890 9908 4896 9920
rect 4663 9880 4896 9908
rect 4663 9877 4675 9880
rect 4617 9871 4675 9877
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 8352 9880 8585 9908
rect 8352 9868 8358 9880
rect 8573 9877 8585 9880
rect 8619 9908 8631 9911
rect 9306 9908 9312 9920
rect 8619 9880 9312 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 3476 9676 4108 9704
rect 3476 9664 3482 9676
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 2041 9639 2099 9645
rect 2041 9605 2053 9639
rect 2087 9636 2099 9639
rect 2130 9636 2136 9648
rect 2087 9608 2136 9636
rect 2087 9605 2099 9608
rect 2041 9599 2099 9605
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 2056 9500 2084 9599
rect 2130 9596 2136 9608
rect 2188 9596 2194 9648
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 2961 9639 3019 9645
rect 2961 9636 2973 9639
rect 2832 9608 2973 9636
rect 2832 9596 2838 9608
rect 2961 9605 2973 9608
rect 3007 9605 3019 9639
rect 4080 9636 4108 9676
rect 4706 9664 4712 9716
rect 4764 9704 4770 9716
rect 4764 9676 5580 9704
rect 4764 9664 4770 9676
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 4080 9608 4537 9636
rect 2961 9599 3019 9605
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 5552 9636 5580 9676
rect 6822 9664 6828 9716
rect 6880 9664 6886 9716
rect 10410 9704 10416 9716
rect 10371 9676 10416 9704
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 13078 9704 13084 9716
rect 13039 9676 13084 9704
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 13446 9704 13452 9716
rect 13407 9676 13452 9704
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 14093 9707 14151 9713
rect 14093 9673 14105 9707
rect 14139 9704 14151 9707
rect 14366 9704 14372 9716
rect 14139 9676 14372 9704
rect 14139 9673 14151 9676
rect 14093 9667 14151 9673
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 5997 9639 6055 9645
rect 5997 9636 6009 9639
rect 5552 9608 6009 9636
rect 4525 9599 4583 9605
rect 5997 9605 6009 9608
rect 6043 9636 6055 9639
rect 6840 9636 6868 9664
rect 6043 9608 6868 9636
rect 10137 9639 10195 9645
rect 6043 9605 6055 9608
rect 5997 9599 6055 9605
rect 10137 9605 10149 9639
rect 10183 9636 10195 9639
rect 10318 9636 10324 9648
rect 10183 9608 10324 9636
rect 10183 9605 10195 9608
rect 10137 9599 10195 9605
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 3786 9568 3792 9580
rect 3651 9540 3792 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 3786 9528 3792 9540
rect 3844 9568 3850 9580
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 3844 9540 4077 9568
rect 3844 9528 3850 9540
rect 4065 9537 4077 9540
rect 4111 9568 4123 9571
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 4111 9540 5181 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 5169 9537 5181 9540
rect 5215 9568 5227 9571
rect 5442 9568 5448 9580
rect 5215 9540 5448 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 9033 9571 9091 9577
rect 9033 9568 9045 9571
rect 8352 9540 9045 9568
rect 8352 9528 8358 9540
rect 9033 9537 9045 9540
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 1443 9472 2084 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4212 9472 4445 9500
rect 4212 9460 4218 9472
rect 4433 9469 4445 9472
rect 4479 9500 4491 9503
rect 4982 9500 4988 9512
rect 4479 9472 4988 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9500 8171 9503
rect 9232 9500 9260 9531
rect 12066 9528 12072 9580
rect 12124 9568 12130 9580
rect 12894 9568 12900 9580
rect 12124 9540 12900 9568
rect 12124 9528 12130 9540
rect 12894 9528 12900 9540
rect 12952 9568 12958 9580
rect 13446 9568 13452 9580
rect 12952 9540 13452 9568
rect 12952 9528 12958 9540
rect 13446 9528 13452 9540
rect 13504 9568 13510 9580
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 13504 9540 14197 9568
rect 13504 9528 13510 9540
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 10318 9500 10324 9512
rect 8159 9472 10324 9500
rect 8159 9469 8171 9472
rect 8113 9463 8171 9469
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 11790 9460 11796 9512
rect 11848 9500 11854 9512
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 11848 9472 12265 9500
rect 11848 9460 11854 9472
rect 12253 9469 12265 9472
rect 12299 9500 12311 9503
rect 12621 9503 12679 9509
rect 12621 9500 12633 9503
rect 12299 9472 12633 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12621 9469 12633 9472
rect 12667 9469 12679 9503
rect 12621 9463 12679 9469
rect 2869 9435 2927 9441
rect 2869 9401 2881 9435
rect 2915 9432 2927 9435
rect 3694 9432 3700 9444
rect 2915 9404 3700 9432
rect 2915 9401 2927 9404
rect 2869 9395 2927 9401
rect 3436 9376 3464 9404
rect 3694 9392 3700 9404
rect 3752 9392 3758 9444
rect 8386 9432 8392 9444
rect 8299 9404 8392 9432
rect 8386 9392 8392 9404
rect 8444 9432 8450 9444
rect 8444 9404 8984 9432
rect 8444 9392 8450 9404
rect 8956 9376 8984 9404
rect 14366 9392 14372 9444
rect 14424 9441 14430 9444
rect 14424 9435 14488 9441
rect 14424 9401 14442 9435
rect 14476 9401 14488 9435
rect 14424 9395 14488 9401
rect 14424 9392 14430 9395
rect 2409 9367 2467 9373
rect 2409 9333 2421 9367
rect 2455 9364 2467 9367
rect 2498 9364 2504 9376
rect 2455 9336 2504 9364
rect 2455 9333 2467 9336
rect 2409 9327 2467 9333
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 3329 9367 3387 9373
rect 3329 9364 3341 9367
rect 3108 9336 3341 9364
rect 3108 9324 3114 9336
rect 3329 9333 3341 9336
rect 3375 9333 3387 9367
rect 3329 9327 3387 9333
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 4893 9367 4951 9373
rect 3476 9336 3521 9364
rect 3476 9324 3482 9336
rect 4893 9333 4905 9367
rect 4939 9364 4951 9367
rect 4982 9364 4988 9376
rect 4939 9336 4988 9364
rect 4939 9333 4951 9336
rect 4893 9327 4951 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5500 9336 5549 9364
rect 5500 9324 5506 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 5537 9327 5595 9333
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 6972 9336 7021 9364
rect 6972 9324 6978 9336
rect 7009 9333 7021 9336
rect 7055 9333 7067 9367
rect 7009 9327 7067 9333
rect 8478 9324 8484 9376
rect 8536 9364 8542 9376
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 8536 9336 8585 9364
rect 8536 9324 8542 9336
rect 8573 9333 8585 9336
rect 8619 9333 8631 9367
rect 8938 9364 8944 9376
rect 8899 9336 8944 9364
rect 8573 9327 8631 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 9858 9364 9864 9376
rect 9815 9336 9864 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 12066 9364 12072 9376
rect 12027 9336 12072 9364
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 15562 9364 15568 9376
rect 15523 9336 15568 9364
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1452 9132 1593 9160
rect 1452 9120 1458 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 1581 9123 1639 9129
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 3326 9120 3332 9172
rect 3384 9160 3390 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3384 9132 4077 9160
rect 3384 9120 3390 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4522 9160 4528 9172
rect 4483 9132 4528 9160
rect 4065 9123 4123 9129
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 8478 9160 8484 9172
rect 8439 9132 8484 9160
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9129 9735 9163
rect 13446 9160 13452 9172
rect 13407 9132 13452 9160
rect 9677 9123 9735 9129
rect 3421 9095 3479 9101
rect 3421 9061 3433 9095
rect 3467 9092 3479 9095
rect 3786 9092 3792 9104
rect 3467 9064 3792 9092
rect 3467 9061 3479 9064
rect 3421 9055 3479 9061
rect 3786 9052 3792 9064
rect 3844 9052 3850 9104
rect 7466 9052 7472 9104
rect 7524 9092 7530 9104
rect 8389 9095 8447 9101
rect 8389 9092 8401 9095
rect 7524 9064 8401 9092
rect 7524 9052 7530 9064
rect 8389 9061 8401 9064
rect 8435 9092 8447 9095
rect 9692 9092 9720 9123
rect 13446 9120 13452 9132
rect 13504 9160 13510 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 13504 9132 14197 9160
rect 13504 9120 13510 9132
rect 14185 9129 14197 9132
rect 14231 9129 14243 9163
rect 26694 9160 26700 9172
rect 26655 9132 26700 9160
rect 14185 9123 14243 9129
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 12066 9092 12072 9104
rect 8435 9064 9720 9092
rect 11348 9064 12072 9092
rect 8435 9061 8447 9064
rect 8389 9055 8447 9061
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2314 9024 2320 9036
rect 1443 8996 2320 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 4430 9024 4436 9036
rect 4391 8996 4436 9024
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 10042 9024 10048 9036
rect 10003 8996 10048 9024
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 11348 9033 11376 9064
rect 12066 9052 12072 9064
rect 12124 9052 12130 9104
rect 11606 9033 11612 9036
rect 11333 9027 11391 9033
rect 11333 8993 11345 9027
rect 11379 8993 11391 9027
rect 11600 9024 11612 9033
rect 11567 8996 11612 9024
rect 11333 8987 11391 8993
rect 11600 8987 11612 8996
rect 11606 8984 11612 8987
rect 11664 8984 11670 9036
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 5442 8956 5448 8968
rect 4755 8928 5448 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 5626 8956 5632 8968
rect 5587 8928 5632 8956
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 8570 8956 8576 8968
rect 8168 8928 8576 8956
rect 8168 8916 8174 8928
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9950 8956 9956 8968
rect 9088 8928 9956 8956
rect 9088 8916 9094 8928
rect 9950 8916 9956 8928
rect 10008 8956 10014 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 10008 8928 10149 8956
rect 10008 8916 10014 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10318 8956 10324 8968
rect 10279 8928 10324 8956
rect 10137 8919 10195 8925
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 13078 8888 13084 8900
rect 13039 8860 13084 8888
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 3050 8820 3056 8832
rect 3011 8792 3056 8820
rect 3050 8780 3056 8792
rect 3108 8780 3114 8832
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 5169 8823 5227 8829
rect 5169 8820 5181 8823
rect 4948 8792 5181 8820
rect 4948 8780 4954 8792
rect 5169 8789 5181 8792
rect 5215 8820 5227 8823
rect 5534 8820 5540 8832
rect 5215 8792 5540 8820
rect 5215 8789 5227 8792
rect 5169 8783 5227 8789
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 8018 8820 8024 8832
rect 7979 8792 8024 8820
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 9214 8820 9220 8832
rect 9175 8792 9220 8820
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 12710 8820 12716 8832
rect 12671 8792 12716 8820
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1544 8588 1593 8616
rect 1544 8576 1550 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 2314 8616 2320 8628
rect 2275 8588 2320 8616
rect 1581 8579 1639 8585
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 3142 8616 3148 8628
rect 3103 8588 3148 8616
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 3786 8616 3792 8628
rect 3747 8588 3792 8616
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4522 8616 4528 8628
rect 4203 8588 4528 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4522 8576 4528 8588
rect 4580 8576 4586 8628
rect 7466 8616 7472 8628
rect 7427 8588 7472 8616
rect 7466 8576 7472 8588
rect 7524 8576 7530 8628
rect 8110 8616 8116 8628
rect 8071 8588 8116 8616
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8478 8616 8484 8628
rect 8439 8588 8484 8616
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11388 8588 12081 8616
rect 11388 8576 11394 8588
rect 12069 8585 12081 8588
rect 12115 8616 12127 8619
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 12115 8588 12173 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27341 8619 27399 8625
rect 27341 8616 27353 8619
rect 26568 8588 27353 8616
rect 26568 8576 26574 8588
rect 27341 8585 27353 8588
rect 27387 8585 27399 8619
rect 27341 8579 27399 8585
rect 2682 8548 2688 8560
rect 2643 8520 2688 8548
rect 2682 8508 2688 8520
rect 2740 8508 2746 8560
rect 3896 8520 6408 8548
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 3896 8480 3924 8520
rect 2087 8452 3924 8480
rect 5813 8483 5871 8489
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6380 8480 6408 8520
rect 6914 8508 6920 8560
rect 6972 8548 6978 8560
rect 7561 8551 7619 8557
rect 7561 8548 7573 8551
rect 6972 8520 7573 8548
rect 6972 8508 6978 8520
rect 7561 8517 7573 8520
rect 7607 8517 7619 8551
rect 26602 8548 26608 8560
rect 26563 8520 26608 8548
rect 7561 8511 7619 8517
rect 26602 8508 26608 8520
rect 26660 8508 26666 8560
rect 27706 8548 27712 8560
rect 27667 8520 27712 8548
rect 27706 8508 27712 8520
rect 27764 8508 27770 8560
rect 8202 8480 8208 8492
rect 5859 8452 6316 8480
rect 6380 8452 8208 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 2056 8412 2084 8443
rect 1443 8384 2084 8412
rect 2501 8415 2559 8421
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2501 8381 2513 8415
rect 2547 8412 2559 8415
rect 3142 8412 3148 8424
rect 2547 8384 3148 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5123 8384 5549 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 5537 8381 5549 8384
rect 5583 8412 5595 8415
rect 5718 8412 5724 8424
rect 5583 8384 5724 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 4430 8344 4436 8356
rect 4391 8316 4436 8344
rect 4430 8304 4436 8316
rect 4488 8304 4494 8356
rect 4890 8304 4896 8356
rect 4948 8344 4954 8356
rect 5629 8347 5687 8353
rect 5629 8344 5641 8347
rect 4948 8316 5641 8344
rect 4948 8304 4954 8316
rect 5629 8313 5641 8316
rect 5675 8313 5687 8347
rect 5629 8307 5687 8313
rect 5166 8276 5172 8288
rect 5127 8248 5172 8276
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 6288 8285 6316 8452
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 9030 8480 9036 8492
rect 8991 8452 9036 8480
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 13354 8480 13360 8492
rect 11664 8452 13360 8480
rect 11664 8440 11670 8452
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 7745 8415 7803 8421
rect 7745 8412 7757 8415
rect 7708 8384 7757 8412
rect 7708 8372 7714 8384
rect 7745 8381 7757 8384
rect 7791 8412 7803 8415
rect 13078 8412 13084 8424
rect 7791 8384 11008 8412
rect 13039 8384 13084 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 8662 8304 8668 8356
rect 8720 8344 8726 8356
rect 9214 8344 9220 8356
rect 8720 8316 9220 8344
rect 8720 8304 8726 8316
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 10980 8353 11008 8384
rect 13078 8372 13084 8384
rect 13136 8372 13142 8424
rect 26418 8412 26424 8424
rect 26379 8384 26424 8412
rect 26418 8372 26424 8384
rect 26476 8412 26482 8424
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26476 8384 26985 8412
rect 26476 8372 26482 8384
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 27522 8412 27528 8424
rect 27483 8384 27528 8412
rect 26973 8375 27031 8381
rect 27522 8372 27528 8384
rect 27580 8412 27586 8424
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 27580 8384 28089 8412
rect 27580 8372 27586 8384
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 10965 8347 11023 8353
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 12069 8347 12127 8353
rect 11011 8316 11100 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 6273 8279 6331 8285
rect 6273 8245 6285 8279
rect 6319 8276 6331 8279
rect 6914 8276 6920 8288
rect 6319 8248 6920 8276
rect 6319 8245 6331 8248
rect 6273 8239 6331 8245
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 11072 8276 11100 8316
rect 12069 8313 12081 8347
rect 12115 8344 12127 8347
rect 12342 8344 12348 8356
rect 12115 8316 12348 8344
rect 12115 8313 12127 8316
rect 12069 8307 12127 8313
rect 12342 8304 12348 8316
rect 12400 8344 12406 8356
rect 13173 8347 13231 8353
rect 13173 8344 13185 8347
rect 12400 8316 13185 8344
rect 12400 8304 12406 8316
rect 13173 8313 13185 8316
rect 13219 8313 13231 8347
rect 13173 8307 13231 8313
rect 11330 8276 11336 8288
rect 11072 8248 11336 8276
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11425 8279 11483 8285
rect 11425 8245 11437 8279
rect 11471 8276 11483 8279
rect 11606 8276 11612 8288
rect 11471 8248 11612 8276
rect 11471 8245 11483 8248
rect 11425 8239 11483 8245
rect 11606 8236 11612 8248
rect 11664 8276 11670 8288
rect 11793 8279 11851 8285
rect 11793 8276 11805 8279
rect 11664 8248 11805 8276
rect 11664 8236 11670 8248
rect 11793 8245 11805 8248
rect 11839 8245 11851 8279
rect 11793 8239 11851 8245
rect 12713 8279 12771 8285
rect 12713 8245 12725 8279
rect 12759 8276 12771 8279
rect 12802 8276 12808 8288
rect 12759 8248 12808 8276
rect 12759 8245 12771 8248
rect 12713 8239 12771 8245
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 16117 8279 16175 8285
rect 16117 8245 16129 8279
rect 16163 8276 16175 8279
rect 16298 8276 16304 8288
rect 16163 8248 16304 8276
rect 16163 8245 16175 8248
rect 16117 8239 16175 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 5442 8072 5448 8084
rect 5403 8044 5448 8072
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 5684 8044 6653 8072
rect 5684 8032 5690 8044
rect 6641 8041 6653 8044
rect 6687 8072 6699 8075
rect 7006 8072 7012 8084
rect 6687 8044 7012 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 7650 8072 7656 8084
rect 7611 8044 7656 8072
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 7837 8075 7895 8081
rect 7837 8041 7849 8075
rect 7883 8072 7895 8075
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 7883 8044 9873 8072
rect 7883 8041 7895 8044
rect 7837 8035 7895 8041
rect 9861 8041 9873 8044
rect 9907 8072 9919 8075
rect 10042 8072 10048 8084
rect 9907 8044 10048 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 11425 8075 11483 8081
rect 11425 8041 11437 8075
rect 11471 8072 11483 8075
rect 11514 8072 11520 8084
rect 11471 8044 11520 8072
rect 11471 8041 11483 8044
rect 11425 8035 11483 8041
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 12066 8072 12072 8084
rect 12027 8044 12072 8072
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12529 8075 12587 8081
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 12710 8072 12716 8084
rect 12575 8044 12716 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 6362 7964 6368 8016
rect 6420 8004 6426 8016
rect 6733 8007 6791 8013
rect 6733 8004 6745 8007
rect 6420 7976 6745 8004
rect 6420 7964 6426 7976
rect 6733 7973 6745 7976
rect 6779 7973 6791 8007
rect 6733 7967 6791 7973
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 2406 7936 2412 7948
rect 1443 7908 2412 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4321 7939 4379 7945
rect 4321 7936 4333 7939
rect 4212 7908 4333 7936
rect 4212 7896 4218 7908
rect 4321 7905 4333 7908
rect 4367 7905 4379 7939
rect 4321 7899 4379 7905
rect 8380 7939 8438 7945
rect 8380 7905 8392 7939
rect 8426 7936 8438 7939
rect 8754 7936 8760 7948
rect 8426 7908 8760 7936
rect 8426 7905 8438 7908
rect 8380 7899 8438 7905
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 3970 7868 3976 7880
rect 2976 7840 3976 7868
rect 2976 7744 3004 7840
rect 3970 7828 3976 7840
rect 4028 7868 4034 7880
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 4028 7840 4077 7868
rect 4028 7828 4034 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 6914 7868 6920 7880
rect 6875 7840 6920 7868
rect 4065 7831 4123 7837
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 7892 7840 8125 7868
rect 7892 7828 7898 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 11514 7868 11520 7880
rect 11475 7840 11520 7868
rect 8113 7831 8171 7837
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 11606 7828 11612 7880
rect 11664 7868 11670 7880
rect 11664 7840 11709 7868
rect 11664 7828 11670 7840
rect 10318 7800 10324 7812
rect 10231 7772 10324 7800
rect 10318 7760 10324 7772
rect 10376 7800 10382 7812
rect 10870 7800 10876 7812
rect 10376 7772 10876 7800
rect 10376 7760 10382 7772
rect 10870 7760 10876 7772
rect 10928 7800 10934 7812
rect 12544 7800 12572 8035
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 13081 8075 13139 8081
rect 13081 8072 13093 8075
rect 13044 8044 13093 8072
rect 13044 8032 13050 8044
rect 13081 8041 13093 8044
rect 13127 8041 13139 8075
rect 13081 8035 13139 8041
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 15562 8072 15568 8084
rect 15436 8044 15568 8072
rect 15436 8032 15442 8044
rect 15562 8032 15568 8044
rect 15620 8072 15626 8084
rect 16209 8075 16267 8081
rect 16209 8072 16221 8075
rect 15620 8044 16221 8072
rect 15620 8032 15626 8044
rect 16209 8041 16221 8044
rect 16255 8072 16267 8075
rect 16390 8072 16396 8084
rect 16255 8044 16396 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 26694 8072 26700 8084
rect 26655 8044 26700 8072
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 13078 7896 13084 7948
rect 13136 7936 13142 7948
rect 13173 7939 13231 7945
rect 13173 7936 13185 7939
rect 13136 7908 13185 7936
rect 13136 7896 13142 7908
rect 13173 7905 13185 7908
rect 13219 7936 13231 7939
rect 13446 7936 13452 7948
rect 13219 7908 13452 7936
rect 13219 7905 13231 7908
rect 13173 7899 13231 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 26510 7936 26516 7948
rect 26471 7908 26516 7936
rect 26510 7896 26516 7908
rect 26568 7896 26574 7948
rect 13354 7868 13360 7880
rect 13315 7840 13360 7868
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 15838 7828 15844 7880
rect 15896 7868 15902 7880
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 15896 7840 16313 7868
rect 15896 7828 15902 7840
rect 16301 7837 16313 7840
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7868 16543 7871
rect 16666 7868 16672 7880
rect 16531 7840 16672 7868
rect 16531 7837 16543 7840
rect 16485 7831 16543 7837
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 12986 7800 12992 7812
rect 10928 7772 12992 7800
rect 10928 7760 10934 7772
rect 12986 7760 12992 7772
rect 13044 7760 13050 7812
rect 2958 7732 2964 7744
rect 2919 7704 2964 7732
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 6270 7732 6276 7744
rect 6231 7704 6276 7732
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 9490 7732 9496 7744
rect 9451 7704 9496 7732
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 10686 7732 10692 7744
rect 10599 7704 10692 7732
rect 10686 7692 10692 7704
rect 10744 7732 10750 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10744 7704 11069 7732
rect 10744 7692 10750 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 12710 7732 12716 7744
rect 12671 7704 12716 7732
rect 11057 7695 11115 7701
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 15841 7735 15899 7741
rect 15841 7732 15853 7735
rect 15804 7704 15853 7732
rect 15804 7692 15810 7704
rect 15841 7701 15853 7704
rect 15887 7701 15899 7735
rect 15841 7695 15899 7701
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 2406 7528 2412 7540
rect 2367 7500 2412 7528
rect 2406 7488 2412 7500
rect 2464 7488 2470 7540
rect 6362 7528 6368 7540
rect 6323 7500 6368 7528
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 7006 7528 7012 7540
rect 6967 7500 7012 7528
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7834 7528 7840 7540
rect 7795 7500 7840 7528
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 8570 7528 8576 7540
rect 8531 7500 8576 7528
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 11609 7531 11667 7537
rect 11609 7528 11621 7531
rect 11480 7500 11621 7528
rect 11480 7488 11486 7500
rect 11609 7497 11621 7500
rect 11655 7497 11667 7531
rect 11790 7528 11796 7540
rect 11751 7500 11796 7528
rect 11609 7491 11667 7497
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 15102 7528 15108 7540
rect 15015 7500 15108 7528
rect 15102 7488 15108 7500
rect 15160 7528 15166 7540
rect 15838 7528 15844 7540
rect 15160 7500 15844 7528
rect 15160 7488 15166 7500
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 26510 7488 26516 7540
rect 26568 7528 26574 7540
rect 27341 7531 27399 7537
rect 27341 7528 27353 7531
rect 26568 7500 27353 7528
rect 26568 7488 26574 7500
rect 27341 7497 27353 7500
rect 27387 7497 27399 7531
rect 27341 7491 27399 7497
rect 1578 7460 1584 7472
rect 1539 7432 1584 7460
rect 1578 7420 1584 7432
rect 1636 7420 1642 7472
rect 2958 7392 2964 7404
rect 2919 7364 2964 7392
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 4706 7352 4712 7404
rect 4764 7392 4770 7404
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4764 7364 5089 7392
rect 4764 7352 4770 7364
rect 5077 7361 5089 7364
rect 5123 7392 5135 7395
rect 5810 7392 5816 7404
rect 5123 7364 5816 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 8588 7392 8616 7488
rect 8754 7420 8760 7472
rect 8812 7460 8818 7472
rect 9769 7463 9827 7469
rect 9769 7460 9781 7463
rect 8812 7432 9781 7460
rect 8812 7420 8818 7432
rect 9769 7429 9781 7432
rect 9815 7460 9827 7463
rect 9815 7432 10916 7460
rect 9815 7429 9827 7432
rect 9769 7423 9827 7429
rect 10888 7404 10916 7432
rect 12250 7420 12256 7472
rect 12308 7460 12314 7472
rect 15381 7463 15439 7469
rect 15381 7460 15393 7463
rect 12308 7432 15393 7460
rect 12308 7420 12314 7432
rect 15381 7429 15393 7432
rect 15427 7429 15439 7463
rect 15381 7423 15439 7429
rect 9217 7395 9275 7401
rect 9217 7392 9229 7395
rect 8588 7364 9229 7392
rect 9217 7361 9229 7364
rect 9263 7392 9275 7395
rect 9490 7392 9496 7404
rect 9263 7364 9496 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 10686 7392 10692 7404
rect 10647 7364 10692 7392
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 10870 7392 10876 7404
rect 10831 7364 10876 7392
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12768 7364 12909 7392
rect 12768 7352 12774 7364
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 3228 7327 3286 7333
rect 3228 7324 3240 7327
rect 1443 7296 2084 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 2056 7200 2084 7296
rect 3160 7296 3240 7324
rect 2869 7259 2927 7265
rect 2869 7225 2881 7259
rect 2915 7256 2927 7259
rect 3160 7256 3188 7296
rect 3228 7293 3240 7296
rect 3274 7324 3286 7327
rect 4724 7324 4752 7352
rect 3274 7296 4752 7324
rect 5537 7327 5595 7333
rect 3274 7293 3286 7296
rect 3228 7287 3286 7293
rect 5537 7293 5549 7327
rect 5583 7324 5595 7327
rect 5626 7324 5632 7336
rect 5583 7296 5632 7324
rect 5583 7293 5595 7296
rect 5537 7287 5595 7293
rect 5626 7284 5632 7296
rect 5684 7324 5690 7336
rect 6270 7324 6276 7336
rect 5684 7296 6276 7324
rect 5684 7284 5690 7296
rect 6270 7284 6276 7296
rect 6328 7284 6334 7336
rect 8205 7327 8263 7333
rect 8205 7293 8217 7327
rect 8251 7324 8263 7327
rect 8754 7324 8760 7336
rect 8251 7296 8760 7324
rect 8251 7293 8263 7296
rect 8205 7287 8263 7293
rect 8754 7284 8760 7296
rect 8812 7284 8818 7336
rect 9122 7324 9128 7336
rect 9083 7296 9128 7324
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 10137 7327 10195 7333
rect 10137 7293 10149 7327
rect 10183 7324 10195 7327
rect 10594 7324 10600 7336
rect 10183 7296 10600 7324
rect 10183 7293 10195 7296
rect 10137 7287 10195 7293
rect 10594 7284 10600 7296
rect 10652 7284 10658 7336
rect 11330 7284 11336 7336
rect 11388 7324 11394 7336
rect 11882 7324 11888 7336
rect 11388 7296 11888 7324
rect 11388 7284 11394 7296
rect 11882 7284 11888 7296
rect 11940 7324 11946 7336
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11940 7296 11989 7324
rect 11940 7284 11946 7296
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 12802 7324 12808 7336
rect 12763 7296 12808 7324
rect 11977 7287 12035 7293
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 12912 7324 12940 7355
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 15396 7392 15424 7423
rect 15562 7420 15568 7472
rect 15620 7460 15626 7472
rect 15749 7463 15807 7469
rect 15749 7460 15761 7463
rect 15620 7432 15761 7460
rect 15620 7420 15626 7432
rect 15749 7429 15761 7432
rect 15795 7429 15807 7463
rect 18138 7460 18144 7472
rect 15749 7423 15807 7429
rect 16408 7432 18144 7460
rect 16408 7401 16436 7432
rect 18138 7420 18144 7432
rect 18196 7420 18202 7472
rect 16393 7395 16451 7401
rect 16393 7392 16405 7395
rect 13044 7364 13089 7392
rect 15396 7364 16405 7392
rect 13044 7352 13050 7364
rect 16393 7361 16405 7364
rect 16439 7361 16451 7395
rect 16393 7355 16451 7361
rect 16577 7395 16635 7401
rect 16577 7361 16589 7395
rect 16623 7392 16635 7395
rect 16666 7392 16672 7404
rect 16623 7364 16672 7392
rect 16623 7361 16635 7364
rect 16577 7355 16635 7361
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 13817 7327 13875 7333
rect 13817 7324 13829 7327
rect 12912 7296 13829 7324
rect 13817 7293 13829 7296
rect 13863 7293 13875 7327
rect 16298 7324 16304 7336
rect 16259 7296 16304 7324
rect 13817 7287 13875 7293
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 26418 7324 26424 7336
rect 26379 7296 26424 7324
rect 26418 7284 26424 7296
rect 26476 7324 26482 7336
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26476 7296 26985 7324
rect 26476 7284 26482 7296
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 26973 7287 27031 7293
rect 9030 7256 9036 7268
rect 2915 7228 3188 7256
rect 8943 7228 9036 7256
rect 2915 7225 2927 7228
rect 2869 7219 2927 7225
rect 9030 7216 9036 7228
rect 9088 7256 9094 7268
rect 12820 7256 12848 7284
rect 14185 7259 14243 7265
rect 14185 7256 14197 7259
rect 9088 7228 10272 7256
rect 12820 7228 14197 7256
rect 9088 7216 9094 7228
rect 2038 7188 2044 7200
rect 1999 7160 2044 7188
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 4341 7191 4399 7197
rect 4341 7188 4353 7191
rect 4212 7160 4353 7188
rect 4212 7148 4218 7160
rect 4341 7157 4353 7160
rect 4387 7188 4399 7191
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 4387 7160 4629 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4617 7157 4629 7160
rect 4663 7157 4675 7191
rect 4617 7151 4675 7157
rect 5074 7148 5080 7200
rect 5132 7188 5138 7200
rect 5169 7191 5227 7197
rect 5169 7188 5181 7191
rect 5132 7160 5181 7188
rect 5132 7148 5138 7160
rect 5169 7157 5181 7160
rect 5215 7157 5227 7191
rect 5169 7151 5227 7157
rect 5258 7148 5264 7200
rect 5316 7188 5322 7200
rect 5629 7191 5687 7197
rect 5629 7188 5641 7191
rect 5316 7160 5641 7188
rect 5316 7148 5322 7160
rect 5629 7157 5641 7160
rect 5675 7157 5687 7191
rect 5629 7151 5687 7157
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 6914 7188 6920 7200
rect 6512 7160 6920 7188
rect 6512 7148 6518 7160
rect 6914 7148 6920 7160
rect 6972 7188 6978 7200
rect 7377 7191 7435 7197
rect 7377 7188 7389 7191
rect 6972 7160 7389 7188
rect 6972 7148 6978 7160
rect 7377 7157 7389 7160
rect 7423 7157 7435 7191
rect 7377 7151 7435 7157
rect 8665 7191 8723 7197
rect 8665 7157 8677 7191
rect 8711 7188 8723 7191
rect 8938 7188 8944 7200
rect 8711 7160 8944 7188
rect 8711 7157 8723 7160
rect 8665 7151 8723 7157
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 10244 7197 10272 7228
rect 14185 7225 14197 7228
rect 14231 7225 14243 7259
rect 14185 7219 14243 7225
rect 10229 7191 10287 7197
rect 10229 7157 10241 7191
rect 10275 7157 10287 7191
rect 11330 7188 11336 7200
rect 11291 7160 11336 7188
rect 10229 7151 10287 7157
rect 11330 7148 11336 7160
rect 11388 7188 11394 7200
rect 11514 7188 11520 7200
rect 11388 7160 11520 7188
rect 11388 7148 11394 7160
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 13446 7188 13452 7200
rect 12492 7160 12537 7188
rect 13407 7160 13452 7188
rect 12492 7148 12498 7160
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 15930 7188 15936 7200
rect 15891 7160 15936 7188
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 16724 7160 16957 7188
rect 16724 7148 16730 7160
rect 16945 7157 16957 7160
rect 16991 7157 17003 7191
rect 26602 7188 26608 7200
rect 26563 7160 26608 7188
rect 16945 7151 17003 7157
rect 26602 7148 26608 7160
rect 26660 7148 26666 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 4157 6987 4215 6993
rect 4157 6984 4169 6987
rect 4028 6956 4169 6984
rect 4028 6944 4034 6956
rect 4157 6953 4169 6956
rect 4203 6984 4215 6987
rect 4249 6987 4307 6993
rect 4249 6984 4261 6987
rect 4203 6956 4261 6984
rect 4203 6953 4215 6956
rect 4157 6947 4215 6953
rect 4249 6953 4261 6956
rect 4295 6953 4307 6987
rect 5626 6984 5632 6996
rect 5587 6956 5632 6984
rect 4249 6947 4307 6953
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 9030 6984 9036 6996
rect 8991 6956 9036 6984
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 10045 6987 10103 6993
rect 10045 6953 10057 6987
rect 10091 6984 10103 6987
rect 10134 6984 10140 6996
rect 10091 6956 10140 6984
rect 10091 6953 10103 6956
rect 10045 6947 10103 6953
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 11149 6987 11207 6993
rect 11149 6953 11161 6987
rect 11195 6984 11207 6987
rect 11606 6984 11612 6996
rect 11195 6956 11612 6984
rect 11195 6953 11207 6956
rect 11149 6947 11207 6953
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 11882 6984 11888 6996
rect 11843 6956 11888 6984
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12805 6987 12863 6993
rect 12805 6953 12817 6987
rect 12851 6984 12863 6987
rect 12894 6984 12900 6996
rect 12851 6956 12900 6984
rect 12851 6953 12863 6956
rect 12805 6947 12863 6953
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 13173 6987 13231 6993
rect 13173 6953 13185 6987
rect 13219 6984 13231 6987
rect 13354 6984 13360 6996
rect 13219 6956 13360 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 15105 6987 15163 6993
rect 15105 6953 15117 6987
rect 15151 6984 15163 6987
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 15151 6956 15669 6984
rect 15151 6953 15163 6956
rect 15105 6947 15163 6953
rect 15657 6953 15669 6956
rect 15703 6984 15715 6987
rect 15930 6984 15936 6996
rect 15703 6956 15936 6984
rect 15703 6953 15715 6956
rect 15657 6947 15715 6953
rect 15930 6944 15936 6956
rect 15988 6944 15994 6996
rect 16298 6984 16304 6996
rect 16259 6956 16304 6984
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 2590 6876 2596 6928
rect 2648 6916 2654 6928
rect 3234 6916 3240 6928
rect 2648 6888 3240 6916
rect 2648 6876 2654 6888
rect 3234 6876 3240 6888
rect 3292 6876 3298 6928
rect 5074 6916 5080 6928
rect 4080 6888 5080 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1946 6848 1952 6860
rect 1443 6820 1952 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2498 6848 2504 6860
rect 2459 6820 2504 6848
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 3145 6851 3203 6857
rect 3145 6817 3157 6851
rect 3191 6848 3203 6851
rect 3418 6848 3424 6860
rect 3191 6820 3424 6848
rect 3191 6817 3203 6820
rect 3145 6811 3203 6817
rect 3418 6808 3424 6820
rect 3476 6848 3482 6860
rect 4080 6848 4108 6888
rect 5074 6876 5080 6888
rect 5132 6876 5138 6928
rect 5810 6876 5816 6928
rect 5868 6916 5874 6928
rect 5868 6888 6868 6916
rect 5868 6876 5874 6888
rect 5166 6848 5172 6860
rect 3476 6820 4108 6848
rect 5127 6820 5172 6848
rect 3476 6808 3482 6820
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 6181 6851 6239 6857
rect 6181 6817 6193 6851
rect 6227 6848 6239 6851
rect 6270 6848 6276 6860
rect 6227 6820 6276 6848
rect 6227 6817 6239 6820
rect 6181 6811 6239 6817
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 6454 6808 6460 6860
rect 6512 6848 6518 6860
rect 6621 6851 6679 6857
rect 6621 6848 6633 6851
rect 6512 6820 6633 6848
rect 6512 6808 6518 6820
rect 6621 6817 6633 6820
rect 6667 6817 6679 6851
rect 6840 6848 6868 6888
rect 8938 6876 8944 6928
rect 8996 6916 9002 6928
rect 15746 6916 15752 6928
rect 8996 6888 9628 6916
rect 15707 6888 15752 6916
rect 8996 6876 9002 6888
rect 8757 6851 8815 6857
rect 6840 6820 7788 6848
rect 6621 6811 6679 6817
rect 6362 6780 6368 6792
rect 6012 6752 6368 6780
rect 1578 6712 1584 6724
rect 1539 6684 1584 6712
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 6012 6721 6040 6752
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 7760 6721 7788 6820
rect 8757 6817 8769 6851
rect 8803 6848 8815 6851
rect 9122 6848 9128 6860
rect 8803 6820 9128 6848
rect 8803 6817 8815 6820
rect 8757 6811 8815 6817
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 9600 6848 9628 6888
rect 15746 6876 15752 6888
rect 15804 6876 15810 6928
rect 26510 6848 26516 6860
rect 9600 6820 9812 6848
rect 26471 6820 26516 6848
rect 9784 6780 9812 6820
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 10134 6780 10140 6792
rect 9784 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10318 6780 10324 6792
rect 10279 6752 10324 6780
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15528 6752 15853 6780
rect 15528 6740 15534 6752
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 4157 6715 4215 6721
rect 4157 6681 4169 6715
rect 4203 6712 4215 6715
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 4203 6684 6009 6712
rect 4203 6681 4215 6684
rect 4157 6675 4215 6681
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 7745 6715 7803 6721
rect 7745 6681 7757 6715
rect 7791 6681 7803 6715
rect 26694 6712 26700 6724
rect 26655 6684 26700 6712
rect 7745 6675 7803 6681
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 2682 6644 2688 6656
rect 2643 6616 2688 6644
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 9674 6644 9680 6656
rect 9635 6616 9680 6644
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 13630 6604 13636 6656
rect 13688 6644 13694 6656
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 13688 6616 13737 6644
rect 13688 6604 13694 6616
rect 13725 6613 13737 6616
rect 13771 6613 13783 6647
rect 13725 6607 13783 6613
rect 15194 6604 15200 6656
rect 15252 6644 15258 6656
rect 15289 6647 15347 6653
rect 15289 6644 15301 6647
rect 15252 6616 15301 6644
rect 15252 6604 15258 6616
rect 15289 6613 15301 6616
rect 15335 6613 15347 6647
rect 16666 6644 16672 6656
rect 16627 6616 16672 6644
rect 15289 6607 15347 6613
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 17034 6644 17040 6656
rect 16995 6616 17040 6644
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1946 6440 1952 6452
rect 1907 6412 1952 6440
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 2498 6440 2504 6452
rect 2459 6412 2504 6440
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 6089 6443 6147 6449
rect 6089 6409 6101 6443
rect 6135 6440 6147 6443
rect 6270 6440 6276 6452
rect 6135 6412 6276 6440
rect 6135 6409 6147 6412
rect 6089 6403 6147 6409
rect 6270 6400 6276 6412
rect 6328 6440 6334 6452
rect 6822 6440 6828 6452
rect 6328 6412 6828 6440
rect 6328 6400 6334 6412
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 8628 6412 8769 6440
rect 8628 6400 8634 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 10318 6440 10324 6452
rect 10279 6412 10324 6440
rect 8757 6403 8815 6409
rect 6362 6332 6368 6384
rect 6420 6372 6426 6384
rect 7009 6375 7067 6381
rect 7009 6372 7021 6375
rect 6420 6344 7021 6372
rect 6420 6332 6426 6344
rect 7009 6341 7021 6344
rect 7055 6341 7067 6375
rect 7009 6335 7067 6341
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6304 3019 6307
rect 3605 6307 3663 6313
rect 3605 6304 3617 6307
rect 3007 6276 3617 6304
rect 3007 6273 3019 6276
rect 2961 6267 3019 6273
rect 3605 6273 3617 6276
rect 3651 6304 3663 6307
rect 4062 6304 4068 6316
rect 3651 6276 4068 6304
rect 3651 6273 3663 6276
rect 3605 6267 3663 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2130 6236 2136 6248
rect 1443 6208 2136 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2130 6196 2136 6208
rect 2188 6196 2194 6248
rect 3418 6236 3424 6248
rect 3379 6208 3424 6236
rect 3418 6196 3424 6208
rect 3476 6196 3482 6248
rect 7024 6236 7052 6335
rect 8772 6304 8800 6403
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 15105 6443 15163 6449
rect 15105 6409 15117 6443
rect 15151 6440 15163 6443
rect 15470 6440 15476 6452
rect 15151 6412 15476 6440
rect 15151 6409 15163 6412
rect 15105 6403 15163 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 10134 6332 10140 6384
rect 10192 6372 10198 6384
rect 10597 6375 10655 6381
rect 10597 6372 10609 6375
rect 10192 6344 10609 6372
rect 10192 6332 10198 6344
rect 10597 6341 10609 6344
rect 10643 6341 10655 6375
rect 10597 6335 10655 6341
rect 8772 6276 9076 6304
rect 8938 6236 8944 6248
rect 7024 6208 8944 6236
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 9048 6236 9076 6276
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 10284 6276 10977 6304
rect 10284 6264 10290 6276
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 13630 6264 13636 6316
rect 13688 6304 13694 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 13688 6276 13737 6304
rect 13688 6264 13694 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 16022 6264 16028 6316
rect 16080 6304 16086 6316
rect 16666 6304 16672 6316
rect 16080 6276 16672 6304
rect 16080 6264 16086 6276
rect 16666 6264 16672 6276
rect 16724 6304 16730 6316
rect 16761 6307 16819 6313
rect 16761 6304 16773 6307
rect 16724 6276 16773 6304
rect 16724 6264 16730 6276
rect 16761 6273 16773 6276
rect 16807 6273 16819 6307
rect 16761 6267 16819 6273
rect 9197 6239 9255 6245
rect 9197 6236 9209 6239
rect 9048 6208 9209 6236
rect 9197 6205 9209 6208
rect 9243 6205 9255 6239
rect 9197 6199 9255 6205
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 12253 6239 12311 6245
rect 12253 6236 12265 6239
rect 11848 6208 12265 6236
rect 11848 6196 11854 6208
rect 12253 6205 12265 6208
rect 12299 6236 12311 6239
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12299 6208 12633 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 12621 6199 12679 6205
rect 16482 6196 16488 6248
rect 16540 6236 16546 6248
rect 16577 6239 16635 6245
rect 16577 6236 16589 6239
rect 16540 6208 16589 6236
rect 16540 6196 16546 6208
rect 16577 6205 16589 6208
rect 16623 6236 16635 6239
rect 17034 6236 17040 6248
rect 16623 6208 17040 6236
rect 16623 6205 16635 6208
rect 16577 6199 16635 6205
rect 17034 6196 17040 6208
rect 17092 6196 17098 6248
rect 26510 6236 26516 6248
rect 26471 6208 26516 6236
rect 26510 6196 26516 6208
rect 26568 6196 26574 6248
rect 13633 6171 13691 6177
rect 13633 6137 13645 6171
rect 13679 6168 13691 6171
rect 13906 6168 13912 6180
rect 13679 6140 13912 6168
rect 13679 6137 13691 6140
rect 13633 6131 13691 6137
rect 13906 6128 13912 6140
rect 13964 6177 13970 6180
rect 13964 6171 14028 6177
rect 13964 6137 13982 6171
rect 14016 6137 14028 6171
rect 13964 6131 14028 6137
rect 13964 6128 13970 6131
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 3053 6103 3111 6109
rect 3053 6100 3065 6103
rect 2740 6072 3065 6100
rect 2740 6060 2746 6072
rect 3053 6069 3065 6072
rect 3099 6069 3111 6103
rect 3053 6063 3111 6069
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 3568 6072 3613 6100
rect 3568 6060 3574 6072
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 6365 6103 6423 6109
rect 6365 6100 6377 6103
rect 5592 6072 6377 6100
rect 5592 6060 5598 6072
rect 6365 6069 6377 6072
rect 6411 6100 6423 6103
rect 6454 6100 6460 6112
rect 6411 6072 6460 6100
rect 6411 6069 6423 6072
rect 6365 6063 6423 6069
rect 6454 6060 6460 6072
rect 6512 6100 6518 6112
rect 6822 6100 6828 6112
rect 6512 6072 6828 6100
rect 6512 6060 6518 6072
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 12069 6103 12127 6109
rect 12069 6069 12081 6103
rect 12115 6100 12127 6103
rect 12434 6100 12440 6112
rect 12115 6072 12440 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 16022 6100 16028 6112
rect 15983 6072 16028 6100
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 16209 6103 16267 6109
rect 16209 6069 16221 6103
rect 16255 6100 16267 6103
rect 16298 6100 16304 6112
rect 16255 6072 16304 6100
rect 16255 6069 16267 6072
rect 16209 6063 16267 6069
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 16669 6103 16727 6109
rect 16669 6069 16681 6103
rect 16715 6100 16727 6103
rect 16850 6100 16856 6112
rect 16715 6072 16856 6100
rect 16715 6069 16727 6072
rect 16669 6063 16727 6069
rect 16850 6060 16856 6072
rect 16908 6100 16914 6112
rect 17221 6103 17279 6109
rect 17221 6100 17233 6103
rect 16908 6072 17233 6100
rect 16908 6060 16914 6072
rect 17221 6069 17233 6072
rect 17267 6069 17279 6103
rect 17221 6063 17279 6069
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 2041 5899 2099 5905
rect 2041 5865 2053 5899
rect 2087 5896 2099 5899
rect 2130 5896 2136 5908
rect 2087 5868 2136 5896
rect 2087 5865 2099 5868
rect 2041 5859 2099 5865
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 3145 5899 3203 5905
rect 3145 5865 3157 5899
rect 3191 5896 3203 5899
rect 3510 5896 3516 5908
rect 3191 5868 3516 5896
rect 3191 5865 3203 5868
rect 3145 5859 3203 5865
rect 3510 5856 3516 5868
rect 3568 5896 3574 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3568 5868 4077 5896
rect 3568 5856 3574 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 6086 5896 6092 5908
rect 6047 5868 6092 5896
rect 4065 5859 4123 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 8938 5896 8944 5908
rect 8899 5868 8944 5896
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 9953 5899 10011 5905
rect 9953 5865 9965 5899
rect 9999 5896 10011 5899
rect 10318 5896 10324 5908
rect 9999 5868 10324 5896
rect 9999 5865 10011 5868
rect 9953 5859 10011 5865
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 13906 5896 13912 5908
rect 13867 5868 13912 5896
rect 13906 5856 13912 5868
rect 13964 5856 13970 5908
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 15746 5896 15752 5908
rect 15151 5868 15752 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 16850 5896 16856 5908
rect 16811 5868 16856 5896
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17313 5899 17371 5905
rect 17313 5865 17325 5899
rect 17359 5896 17371 5899
rect 17586 5896 17592 5908
rect 17359 5868 17592 5896
rect 17359 5865 17371 5868
rect 17313 5859 17371 5865
rect 17586 5856 17592 5868
rect 17644 5856 17650 5908
rect 26694 5896 26700 5908
rect 26655 5868 26700 5896
rect 26694 5856 26700 5868
rect 26752 5856 26758 5908
rect 5994 5828 6000 5840
rect 5907 5800 6000 5828
rect 5994 5788 6000 5800
rect 6052 5828 6058 5840
rect 6546 5828 6552 5840
rect 6052 5800 6552 5828
rect 6052 5788 6058 5800
rect 6546 5788 6552 5800
rect 6604 5788 6610 5840
rect 10336 5828 10364 5856
rect 10566 5831 10624 5837
rect 10566 5828 10578 5831
rect 10336 5800 10578 5828
rect 10566 5797 10578 5800
rect 10612 5797 10624 5831
rect 10566 5791 10624 5797
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 12774 5831 12832 5837
rect 12774 5828 12786 5831
rect 12584 5800 12786 5828
rect 12584 5788 12590 5800
rect 12774 5797 12786 5800
rect 12820 5797 12832 5831
rect 13924 5828 13952 5856
rect 16022 5828 16028 5840
rect 13924 5800 16028 5828
rect 12774 5791 12832 5797
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 2406 5760 2412 5772
rect 1443 5732 2412 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 2406 5720 2412 5732
rect 2464 5720 2470 5772
rect 3881 5763 3939 5769
rect 3881 5729 3893 5763
rect 3927 5760 3939 5763
rect 4338 5760 4344 5772
rect 3927 5732 4344 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 4338 5720 4344 5732
rect 4396 5760 4402 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4396 5732 4445 5760
rect 4396 5720 4402 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10410 5760 10416 5772
rect 10367 5732 10416 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 13078 5760 13084 5772
rect 12492 5732 13084 5760
rect 12492 5720 12498 5732
rect 4522 5692 4528 5704
rect 4483 5664 4528 5692
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 4706 5692 4712 5704
rect 4667 5664 4712 5692
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 6270 5692 6276 5704
rect 6231 5664 6276 5692
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 12544 5701 12572 5732
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 15378 5720 15384 5772
rect 15436 5760 15442 5772
rect 15657 5763 15715 5769
rect 15657 5760 15669 5763
rect 15436 5732 15669 5760
rect 15436 5720 15442 5732
rect 15657 5729 15669 5732
rect 15703 5729 15715 5763
rect 15657 5723 15715 5729
rect 15856 5704 15884 5800
rect 16022 5788 16028 5800
rect 16080 5788 16086 5840
rect 17218 5760 17224 5772
rect 17179 5732 17224 5760
rect 17218 5720 17224 5732
rect 17276 5720 17282 5772
rect 26510 5760 26516 5772
rect 26471 5732 26516 5760
rect 26510 5720 26516 5732
rect 26568 5720 26574 5772
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5661 12587 5695
rect 15746 5692 15752 5704
rect 15707 5664 15752 5692
rect 12529 5655 12587 5661
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 15838 5652 15844 5704
rect 15896 5692 15902 5704
rect 17405 5695 17463 5701
rect 15896 5664 15989 5692
rect 15896 5652 15902 5664
rect 17405 5661 17417 5695
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 4724 5624 4752 5652
rect 4120 5596 4752 5624
rect 4120 5584 4126 5596
rect 16206 5584 16212 5636
rect 16264 5624 16270 5636
rect 16393 5627 16451 5633
rect 16393 5624 16405 5627
rect 16264 5596 16405 5624
rect 16264 5584 16270 5596
rect 16393 5593 16405 5596
rect 16439 5624 16451 5627
rect 16942 5624 16948 5636
rect 16439 5596 16948 5624
rect 16439 5593 16451 5596
rect 16393 5587 16451 5593
rect 16942 5584 16948 5596
rect 17000 5624 17006 5636
rect 17420 5624 17448 5655
rect 17000 5596 17448 5624
rect 17000 5584 17006 5596
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 5169 5559 5227 5565
rect 5169 5556 5181 5559
rect 4856 5528 5181 5556
rect 4856 5516 4862 5528
rect 5169 5525 5181 5528
rect 5215 5556 5227 5559
rect 5629 5559 5687 5565
rect 5629 5556 5641 5559
rect 5215 5528 5641 5556
rect 5215 5525 5227 5528
rect 5169 5519 5227 5525
rect 5629 5525 5641 5528
rect 5675 5525 5687 5559
rect 5629 5519 5687 5525
rect 11701 5559 11759 5565
rect 11701 5525 11713 5559
rect 11747 5556 11759 5559
rect 12526 5556 12532 5568
rect 11747 5528 12532 5556
rect 11747 5525 11759 5528
rect 11701 5519 11759 5525
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 13630 5516 13636 5568
rect 13688 5556 13694 5568
rect 14185 5559 14243 5565
rect 14185 5556 14197 5559
rect 13688 5528 14197 5556
rect 13688 5516 13694 5528
rect 14185 5525 14197 5528
rect 14231 5525 14243 5559
rect 15286 5556 15292 5568
rect 15247 5528 15292 5556
rect 14185 5519 14243 5525
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 2406 5352 2412 5364
rect 2367 5324 2412 5352
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 3513 5355 3571 5361
rect 3513 5321 3525 5355
rect 3559 5352 3571 5355
rect 4062 5352 4068 5364
rect 3559 5324 4068 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4338 5352 4344 5364
rect 4299 5324 4344 5352
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 5718 5352 5724 5364
rect 5679 5324 5724 5352
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 6328 5324 6377 5352
rect 6328 5312 6334 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 10318 5352 10324 5364
rect 10279 5324 10324 5352
rect 6365 5315 6423 5321
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 10689 5355 10747 5361
rect 10689 5352 10701 5355
rect 10468 5324 10701 5352
rect 10468 5312 10474 5324
rect 10689 5321 10701 5324
rect 10735 5321 10747 5355
rect 10689 5315 10747 5321
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 12621 5355 12679 5361
rect 12621 5352 12633 5355
rect 12584 5324 12633 5352
rect 12584 5312 12590 5324
rect 12621 5321 12633 5324
rect 12667 5321 12679 5355
rect 12621 5315 12679 5321
rect 15749 5355 15807 5361
rect 15749 5321 15761 5355
rect 15795 5352 15807 5355
rect 15838 5352 15844 5364
rect 15795 5324 15844 5352
rect 15795 5321 15807 5324
rect 15749 5315 15807 5321
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 16393 5355 16451 5361
rect 16393 5321 16405 5355
rect 16439 5352 16451 5355
rect 16482 5352 16488 5364
rect 16439 5324 16488 5352
rect 16439 5321 16451 5324
rect 16393 5315 16451 5321
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 17218 5312 17224 5364
rect 17276 5352 17282 5364
rect 17773 5355 17831 5361
rect 17773 5352 17785 5355
rect 17276 5324 17785 5352
rect 17276 5312 17282 5324
rect 17773 5321 17785 5324
rect 17819 5352 17831 5355
rect 17862 5352 17868 5364
rect 17819 5324 17868 5352
rect 17819 5321 17831 5324
rect 17773 5315 17831 5321
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 26602 5352 26608 5364
rect 26563 5324 26608 5352
rect 26602 5312 26608 5324
rect 26660 5312 26666 5364
rect 3881 5287 3939 5293
rect 3881 5253 3893 5287
rect 3927 5284 3939 5287
rect 5534 5284 5540 5296
rect 3927 5256 5540 5284
rect 3927 5253 3939 5256
rect 3881 5247 3939 5253
rect 4908 5228 4936 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 6089 5287 6147 5293
rect 6089 5253 6101 5287
rect 6135 5284 6147 5287
rect 6546 5284 6552 5296
rect 6135 5256 6552 5284
rect 6135 5253 6147 5256
rect 6089 5247 6147 5253
rect 6546 5244 6552 5256
rect 6604 5244 6610 5296
rect 16301 5287 16359 5293
rect 16301 5253 16313 5287
rect 16347 5284 16359 5287
rect 16574 5284 16580 5296
rect 16347 5256 16580 5284
rect 16347 5253 16359 5256
rect 16301 5247 16359 5253
rect 16574 5244 16580 5256
rect 16632 5244 16638 5296
rect 17497 5287 17555 5293
rect 17497 5253 17509 5287
rect 17543 5284 17555 5287
rect 17586 5284 17592 5296
rect 17543 5256 17592 5284
rect 17543 5253 17555 5256
rect 17497 5247 17555 5253
rect 17586 5244 17592 5256
rect 17644 5244 17650 5296
rect 4798 5216 4804 5228
rect 4759 5188 4804 5216
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 4890 5176 4896 5228
rect 4948 5216 4954 5228
rect 13541 5219 13599 5225
rect 4948 5188 4993 5216
rect 4948 5176 4954 5188
rect 13541 5185 13553 5219
rect 13587 5216 13599 5219
rect 16942 5216 16948 5228
rect 13587 5188 13768 5216
rect 16903 5188 16948 5216
rect 13587 5185 13599 5188
rect 13541 5179 13599 5185
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 4249 5151 4307 5157
rect 1443 5120 2084 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 2056 5024 2084 5120
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 4706 5148 4712 5160
rect 4295 5120 4712 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 13630 5148 13636 5160
rect 13096 5120 13636 5148
rect 13096 5024 13124 5120
rect 13630 5108 13636 5120
rect 13688 5108 13694 5160
rect 13740 5148 13768 5188
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 13900 5151 13958 5157
rect 13900 5148 13912 5151
rect 13740 5120 13912 5148
rect 13900 5117 13912 5120
rect 13946 5148 13958 5151
rect 15470 5148 15476 5160
rect 13946 5120 15476 5148
rect 13946 5117 13958 5120
rect 13900 5111 13958 5117
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 16206 5108 16212 5160
rect 16264 5148 16270 5160
rect 16758 5148 16764 5160
rect 16264 5120 16764 5148
rect 16264 5108 16270 5120
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 26421 5151 26479 5157
rect 26421 5148 26433 5151
rect 26344 5120 26433 5148
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 16853 5083 16911 5089
rect 16853 5080 16865 5083
rect 16632 5052 16865 5080
rect 16632 5040 16638 5052
rect 16853 5049 16865 5052
rect 16899 5080 16911 5083
rect 18138 5080 18144 5092
rect 16899 5052 18144 5080
rect 16899 5049 16911 5052
rect 16853 5043 16911 5049
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 26344 5024 26372 5120
rect 26421 5117 26433 5120
rect 26467 5117 26479 5151
rect 26421 5111 26479 5117
rect 26510 5108 26516 5160
rect 26568 5148 26574 5160
rect 26973 5151 27031 5157
rect 26973 5148 26985 5151
rect 26568 5120 26985 5148
rect 26568 5108 26574 5120
rect 26973 5117 26985 5120
rect 27019 5117 27031 5151
rect 26973 5111 27031 5117
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 1581 5015 1639 5021
rect 1581 5012 1593 5015
rect 1452 4984 1593 5012
rect 1452 4972 1458 4984
rect 1581 4981 1593 4984
rect 1627 4981 1639 5015
rect 2038 5012 2044 5024
rect 1999 4984 2044 5012
rect 1581 4975 1639 4981
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 13078 5012 13084 5024
rect 13039 4984 13084 5012
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 15013 5015 15071 5021
rect 15013 5012 15025 5015
rect 14332 4984 15025 5012
rect 14332 4972 14338 4984
rect 15013 4981 15025 4984
rect 15059 4981 15071 5015
rect 15378 5012 15384 5024
rect 15339 4984 15384 5012
rect 15013 4975 15071 4981
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 26326 5012 26332 5024
rect 26287 4984 26332 5012
rect 26326 4972 26332 4984
rect 26384 4972 26390 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4808 2099 4811
rect 2314 4808 2320 4820
rect 2087 4780 2320 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 2056 4672 2084 4771
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 3881 4811 3939 4817
rect 3881 4777 3893 4811
rect 3927 4808 3939 4811
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 3927 4780 4261 4808
rect 3927 4777 3939 4780
rect 3881 4771 3939 4777
rect 4249 4777 4261 4780
rect 4295 4808 4307 4811
rect 4522 4808 4528 4820
rect 4295 4780 4528 4808
rect 4295 4777 4307 4780
rect 4249 4771 4307 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 6972 4780 7389 4808
rect 6972 4768 6978 4780
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 10226 4808 10232 4820
rect 10139 4780 10232 4808
rect 7377 4771 7435 4777
rect 10226 4768 10232 4780
rect 10284 4808 10290 4820
rect 10410 4808 10416 4820
rect 10284 4780 10416 4808
rect 10284 4768 10290 4780
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 13722 4768 13728 4820
rect 13780 4808 13786 4820
rect 14001 4811 14059 4817
rect 14001 4808 14013 4811
rect 13780 4780 14013 4808
rect 13780 4768 13786 4780
rect 14001 4777 14013 4780
rect 14047 4808 14059 4811
rect 15102 4808 15108 4820
rect 14047 4780 15108 4808
rect 14047 4777 14059 4780
rect 14001 4771 14059 4777
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 15565 4811 15623 4817
rect 15565 4777 15577 4811
rect 15611 4808 15623 4811
rect 15746 4808 15752 4820
rect 15611 4780 15752 4808
rect 15611 4777 15623 4780
rect 15565 4771 15623 4777
rect 15746 4768 15752 4780
rect 15804 4808 15810 4820
rect 16669 4811 16727 4817
rect 16669 4808 16681 4811
rect 15804 4780 16681 4808
rect 15804 4768 15810 4780
rect 16669 4777 16681 4780
rect 16715 4777 16727 4811
rect 17126 4808 17132 4820
rect 17087 4780 17132 4808
rect 16669 4771 16727 4777
rect 17126 4768 17132 4780
rect 17184 4768 17190 4820
rect 19886 4768 19892 4820
rect 19944 4808 19950 4820
rect 20070 4808 20076 4820
rect 19944 4780 20076 4808
rect 19944 4768 19950 4780
rect 20070 4768 20076 4780
rect 20128 4768 20134 4820
rect 26694 4808 26700 4820
rect 26655 4780 26700 4808
rect 26694 4768 26700 4780
rect 26752 4768 26758 4820
rect 4617 4743 4675 4749
rect 4617 4709 4629 4743
rect 4663 4740 4675 4743
rect 4706 4740 4712 4752
rect 4663 4712 4712 4740
rect 4663 4709 4675 4712
rect 4617 4703 4675 4709
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 6270 4749 6276 4752
rect 5353 4743 5411 4749
rect 5353 4709 5365 4743
rect 5399 4740 5411 4743
rect 6264 4740 6276 4749
rect 5399 4712 6276 4740
rect 5399 4709 5411 4712
rect 5353 4703 5411 4709
rect 6264 4703 6276 4712
rect 6270 4700 6276 4703
rect 6328 4700 6334 4752
rect 6362 4700 6368 4752
rect 6420 4700 6426 4752
rect 16206 4700 16212 4752
rect 16264 4740 16270 4752
rect 16393 4743 16451 4749
rect 16393 4740 16405 4743
rect 16264 4712 16405 4740
rect 16264 4700 16270 4712
rect 16393 4709 16405 4712
rect 16439 4709 16451 4743
rect 17034 4740 17040 4752
rect 16995 4712 17040 4740
rect 16393 4703 16451 4709
rect 17034 4700 17040 4712
rect 17092 4700 17098 4752
rect 1443 4644 2084 4672
rect 2501 4675 2559 4681
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 2501 4641 2513 4675
rect 2547 4672 2559 4675
rect 2774 4672 2780 4684
rect 2547 4644 2780 4672
rect 2547 4641 2559 4644
rect 2501 4635 2559 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 5997 4675 6055 4681
rect 5997 4672 6009 4675
rect 5592 4644 6009 4672
rect 5592 4632 5598 4644
rect 5997 4641 6009 4644
rect 6043 4672 6055 4675
rect 6380 4672 6408 4700
rect 6043 4644 6408 4672
rect 10505 4675 10563 4681
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 10505 4641 10517 4675
rect 10551 4672 10563 4675
rect 10594 4672 10600 4684
rect 10551 4644 10600 4672
rect 10551 4641 10563 4644
rect 10505 4635 10563 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17402 4672 17408 4684
rect 17000 4644 17408 4672
rect 17000 4632 17006 4644
rect 4614 4564 4620 4616
rect 4672 4604 4678 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4672 4576 4721 4604
rect 4672 4564 4678 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 4890 4604 4896 4616
rect 4851 4576 4896 4604
rect 4709 4567 4767 4573
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 14090 4604 14096 4616
rect 14051 4576 14096 4604
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 17236 4613 17264 4644
rect 17402 4632 17408 4644
rect 17460 4672 17466 4684
rect 17681 4675 17739 4681
rect 17681 4672 17693 4675
rect 17460 4644 17693 4672
rect 17460 4632 17466 4644
rect 17681 4641 17693 4644
rect 17727 4641 17739 4675
rect 17681 4635 17739 4641
rect 26418 4632 26424 4684
rect 26476 4672 26482 4684
rect 26513 4675 26571 4681
rect 26513 4672 26525 4675
rect 26476 4644 26525 4672
rect 26476 4632 26482 4644
rect 26513 4641 26525 4644
rect 26559 4641 26571 4675
rect 26513 4635 26571 4641
rect 17221 4607 17279 4613
rect 17221 4573 17233 4607
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 1670 4496 1676 4548
rect 1728 4536 1734 4548
rect 2685 4539 2743 4545
rect 2685 4536 2697 4539
rect 1728 4508 2697 4536
rect 1728 4496 1734 4508
rect 2685 4505 2697 4508
rect 2731 4505 2743 4539
rect 2685 4499 2743 4505
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 10689 4471 10747 4477
rect 10689 4437 10701 4471
rect 10735 4468 10747 4471
rect 11698 4468 11704 4480
rect 10735 4440 11704 4468
rect 10735 4437 10747 4440
rect 10689 4431 10747 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 13630 4468 13636 4480
rect 13591 4440 13636 4468
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 6181 4267 6239 4273
rect 6181 4233 6193 4267
rect 6227 4264 6239 4267
rect 6270 4264 6276 4276
rect 6227 4236 6276 4264
rect 6227 4233 6239 4236
rect 6181 4227 6239 4233
rect 2406 4128 2412 4140
rect 2367 4100 2412 4128
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2832 4100 3065 4128
rect 2832 4088 2838 4100
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 3053 4091 3111 4097
rect 3620 4100 4261 4128
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 2424 4060 2452 4088
rect 3620 4069 3648 4100
rect 4249 4097 4261 4100
rect 4295 4128 4307 4131
rect 4982 4128 4988 4140
rect 4295 4100 4988 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5350 4128 5356 4140
rect 5263 4100 5356 4128
rect 5350 4088 5356 4100
rect 5408 4128 5414 4140
rect 6196 4128 6224 4227
rect 6270 4224 6276 4236
rect 6328 4224 6334 4276
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 6420 4236 6469 4264
rect 6420 4224 6426 4236
rect 6457 4233 6469 4236
rect 6503 4233 6515 4267
rect 14090 4264 14096 4276
rect 14051 4236 14096 4264
rect 6457 4227 6515 4233
rect 14090 4224 14096 4236
rect 14148 4264 14154 4276
rect 15197 4267 15255 4273
rect 15197 4264 15209 4267
rect 14148 4236 15209 4264
rect 14148 4224 14154 4236
rect 15197 4233 15209 4236
rect 15243 4233 15255 4267
rect 17034 4264 17040 4276
rect 16995 4236 17040 4264
rect 15197 4227 15255 4233
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 17402 4264 17408 4276
rect 17363 4236 17408 4264
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 26418 4224 26424 4276
rect 26476 4264 26482 4276
rect 27341 4267 27399 4273
rect 27341 4264 27353 4267
rect 26476 4236 27353 4264
rect 26476 4224 26482 4236
rect 27341 4233 27353 4236
rect 27387 4233 27399 4267
rect 27341 4227 27399 4233
rect 14274 4196 14280 4208
rect 13832 4168 14280 4196
rect 5408 4100 6224 4128
rect 13725 4131 13783 4137
rect 5408 4088 5414 4100
rect 13725 4097 13737 4131
rect 13771 4128 13783 4131
rect 13832 4128 13860 4168
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 15105 4199 15163 4205
rect 15105 4165 15117 4199
rect 15151 4196 15163 4199
rect 15470 4196 15476 4208
rect 15151 4168 15476 4196
rect 15151 4165 15163 4168
rect 15105 4159 15163 4165
rect 15470 4156 15476 4168
rect 15528 4196 15534 4208
rect 16761 4199 16819 4205
rect 15528 4168 15792 4196
rect 15528 4156 15534 4168
rect 15764 4137 15792 4168
rect 16761 4165 16773 4199
rect 16807 4196 16819 4199
rect 17126 4196 17132 4208
rect 16807 4168 17132 4196
rect 16807 4165 16819 4168
rect 16761 4159 16819 4165
rect 17126 4156 17132 4168
rect 17184 4156 17190 4208
rect 13771 4100 13860 4128
rect 14737 4131 14795 4137
rect 13771 4097 13783 4100
rect 13725 4091 13783 4097
rect 14737 4097 14749 4131
rect 14783 4128 14795 4131
rect 15749 4131 15807 4137
rect 14783 4100 15700 4128
rect 14783 4097 14795 4100
rect 14737 4091 14795 4097
rect 2501 4063 2559 4069
rect 2501 4060 2513 4063
rect 1443 4032 2084 4060
rect 2424 4032 2513 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 2056 4001 2084 4032
rect 2501 4029 2513 4032
rect 2547 4029 2559 4063
rect 2501 4023 2559 4029
rect 3605 4063 3663 4069
rect 3605 4029 3617 4063
rect 3651 4029 3663 4063
rect 4522 4060 4528 4072
rect 4483 4032 4528 4060
rect 3605 4023 3663 4029
rect 4522 4020 4528 4032
rect 4580 4060 4586 4072
rect 5074 4060 5080 4072
rect 4580 4032 4936 4060
rect 5035 4032 5080 4060
rect 4580 4020 4586 4032
rect 2041 3995 2099 4001
rect 2041 3961 2053 3995
rect 2087 3992 2099 3995
rect 2590 3992 2596 4004
rect 2087 3964 2596 3992
rect 2087 3961 2099 3964
rect 2041 3955 2099 3961
rect 2590 3952 2596 3964
rect 2648 3952 2654 4004
rect 3513 3995 3571 4001
rect 3513 3961 3525 3995
rect 3559 3992 3571 3995
rect 4614 3992 4620 4004
rect 3559 3964 4620 3992
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 4908 3992 4936 4032
rect 5074 4020 5080 4032
rect 5132 4060 5138 4072
rect 5721 4063 5779 4069
rect 5721 4060 5733 4063
rect 5132 4032 5733 4060
rect 5132 4020 5138 4032
rect 5721 4029 5733 4032
rect 5767 4029 5779 4063
rect 5721 4023 5779 4029
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4060 10195 4063
rect 10226 4060 10232 4072
rect 10183 4032 10232 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10226 4020 10232 4032
rect 10284 4020 10290 4072
rect 10404 4063 10462 4069
rect 10404 4060 10416 4063
rect 10397 4029 10416 4060
rect 10450 4060 10462 4063
rect 13740 4060 13768 4091
rect 10450 4032 13768 4060
rect 10450 4029 10462 4032
rect 10397 4023 10462 4029
rect 5169 3995 5227 4001
rect 5169 3992 5181 3995
rect 4908 3964 5181 3992
rect 5169 3961 5181 3964
rect 5215 3961 5227 3995
rect 5169 3955 5227 3961
rect 10045 3995 10103 4001
rect 10045 3961 10057 3995
rect 10091 3992 10103 3995
rect 10397 3992 10425 4023
rect 15286 4020 15292 4072
rect 15344 4060 15350 4072
rect 15672 4069 15700 4100
rect 15749 4097 15761 4131
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 15565 4063 15623 4069
rect 15565 4060 15577 4063
rect 15344 4032 15577 4060
rect 15344 4020 15350 4032
rect 15565 4029 15577 4032
rect 15611 4029 15623 4063
rect 15565 4023 15623 4029
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4060 15715 4063
rect 16298 4060 16304 4072
rect 15703 4032 16304 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 26418 4060 26424 4072
rect 26331 4032 26424 4060
rect 26418 4020 26424 4032
rect 26476 4060 26482 4072
rect 26973 4063 27031 4069
rect 26973 4060 26985 4063
rect 26476 4032 26985 4060
rect 26476 4020 26482 4032
rect 26973 4029 26985 4032
rect 27019 4029 27031 4063
rect 26973 4023 27031 4029
rect 10091 3964 10425 3992
rect 13357 3995 13415 4001
rect 10091 3961 10103 3964
rect 10045 3955 10103 3961
rect 13357 3961 13369 3995
rect 13403 3992 13415 3995
rect 13722 3992 13728 4004
rect 13403 3964 13728 3992
rect 13403 3961 13415 3964
rect 13357 3955 13415 3961
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 2774 3924 2780 3936
rect 2731 3896 2780 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 3786 3924 3792 3936
rect 3747 3896 3792 3924
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4706 3924 4712 3936
rect 4667 3896 4712 3924
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 10652 3896 11529 3924
rect 10652 3884 10658 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 26602 3924 26608 3936
rect 26563 3896 26608 3924
rect 11517 3887 11575 3893
rect 26602 3884 26608 3896
rect 26660 3884 26666 3936
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 4706 3720 4712 3732
rect 3927 3692 4712 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 5074 3720 5080 3732
rect 5035 3692 5080 3720
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 10594 3720 10600 3732
rect 10555 3692 10600 3720
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 15344 3692 15485 3720
rect 15344 3680 15350 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 26694 3720 26700 3732
rect 26655 3692 26700 3720
rect 15473 3683 15531 3689
rect 26694 3680 26700 3692
rect 26752 3680 26758 3732
rect 4341 3655 4399 3661
rect 4341 3621 4353 3655
rect 4387 3652 4399 3655
rect 4890 3652 4896 3664
rect 4387 3624 4896 3652
rect 4387 3621 4399 3624
rect 4341 3615 4399 3621
rect 4890 3612 4896 3624
rect 4948 3612 4954 3664
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3584 1455 3587
rect 1762 3584 1768 3596
rect 1443 3556 1768 3584
rect 1443 3553 1455 3556
rect 1397 3547 1455 3553
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3584 2743 3587
rect 2958 3584 2964 3596
rect 2731 3556 2964 3584
rect 2731 3553 2743 3556
rect 2685 3547 2743 3553
rect 2958 3544 2964 3556
rect 3016 3584 3022 3596
rect 4062 3584 4068 3596
rect 3016 3556 4068 3584
rect 3016 3544 3022 3556
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 11517 3587 11575 3593
rect 11517 3584 11529 3587
rect 10284 3556 11529 3584
rect 10284 3544 10290 3556
rect 11517 3553 11529 3556
rect 11563 3584 11575 3587
rect 11606 3584 11612 3596
rect 11563 3556 11612 3584
rect 11563 3553 11575 3556
rect 11517 3547 11575 3553
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 11790 3593 11796 3596
rect 11784 3584 11796 3593
rect 11751 3556 11796 3584
rect 11784 3547 11796 3556
rect 11790 3544 11796 3547
rect 11848 3544 11854 3596
rect 15194 3544 15200 3596
rect 15252 3584 15258 3596
rect 15841 3587 15899 3593
rect 15841 3584 15853 3587
rect 15252 3556 15853 3584
rect 15252 3544 15258 3556
rect 15841 3553 15853 3556
rect 15887 3553 15899 3587
rect 25314 3584 25320 3596
rect 25275 3556 25320 3584
rect 15841 3547 15899 3553
rect 25314 3544 25320 3556
rect 25372 3544 25378 3596
rect 26513 3587 26571 3593
rect 26513 3553 26525 3587
rect 26559 3584 26571 3587
rect 26786 3584 26792 3596
rect 26559 3556 26792 3584
rect 26559 3553 26571 3556
rect 26513 3547 26571 3553
rect 26786 3544 26792 3556
rect 26844 3544 26850 3596
rect 1486 3476 1492 3528
rect 1544 3516 1550 3528
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 1544 3488 1593 3516
rect 1544 3476 1550 3488
rect 1581 3485 1593 3488
rect 1627 3485 1639 3519
rect 5166 3516 5172 3528
rect 5127 3488 5172 3516
rect 1581 3479 1639 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5350 3516 5356 3528
rect 5311 3488 5356 3516
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 22094 3476 22100 3528
rect 22152 3516 22158 3528
rect 23198 3516 23204 3528
rect 22152 3488 23204 3516
rect 22152 3476 22158 3488
rect 23198 3476 23204 3488
rect 23256 3476 23262 3528
rect 4614 3408 4620 3460
rect 4672 3448 4678 3460
rect 4709 3451 4767 3457
rect 4709 3448 4721 3451
rect 4672 3420 4721 3448
rect 4672 3408 4678 3420
rect 4709 3417 4721 3420
rect 4755 3417 4767 3451
rect 4709 3411 4767 3417
rect 9861 3451 9919 3457
rect 9861 3417 9873 3451
rect 9907 3448 9919 3451
rect 10778 3448 10784 3460
rect 9907 3420 10784 3448
rect 9907 3417 9919 3420
rect 9861 3411 9919 3417
rect 10778 3408 10784 3420
rect 10836 3408 10842 3460
rect 2866 3380 2872 3392
rect 2827 3352 2872 3380
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 12894 3380 12900 3392
rect 12855 3352 12900 3380
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13078 3340 13084 3392
rect 13136 3380 13142 3392
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 13136 3352 13185 3380
rect 13136 3340 13142 3352
rect 13173 3349 13185 3352
rect 13219 3349 13231 3383
rect 13173 3343 13231 3349
rect 16025 3383 16083 3389
rect 16025 3349 16037 3383
rect 16071 3380 16083 3383
rect 16942 3380 16948 3392
rect 16071 3352 16948 3380
rect 16071 3349 16083 3352
rect 16025 3343 16083 3349
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 25501 3383 25559 3389
rect 25501 3349 25513 3383
rect 25547 3380 25559 3383
rect 25866 3380 25872 3392
rect 25547 3352 25872 3380
rect 25547 3349 25559 3352
rect 25501 3343 25559 3349
rect 25866 3340 25872 3352
rect 25924 3340 25930 3392
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 1765 3179 1823 3185
rect 1765 3145 1777 3179
rect 1811 3176 1823 3179
rect 2682 3176 2688 3188
rect 1811 3148 2688 3176
rect 1811 3145 1823 3148
rect 1765 3139 1823 3145
rect 1872 2981 1900 3148
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 2958 3176 2964 3188
rect 2823 3148 2964 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3789 3179 3847 3185
rect 3789 3145 3801 3179
rect 3835 3176 3847 3179
rect 3878 3176 3884 3188
rect 3835 3148 3884 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2972 3203 2975
rect 3804 2972 3832 3139
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4798 3176 4804 3188
rect 4711 3148 4804 3176
rect 4798 3136 4804 3148
rect 4856 3176 4862 3188
rect 5166 3176 5172 3188
rect 4856 3148 5172 3176
rect 4856 3136 4862 3148
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 5810 3176 5816 3188
rect 5408 3148 5816 3176
rect 5408 3136 5414 3148
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 8846 3176 8852 3188
rect 8807 3148 8852 3176
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 25130 3176 25136 3188
rect 25091 3148 25136 3176
rect 25130 3136 25136 3148
rect 25188 3136 25194 3188
rect 25314 3136 25320 3188
rect 25372 3176 25378 3188
rect 25869 3179 25927 3185
rect 25869 3176 25881 3179
rect 25372 3148 25881 3176
rect 25372 3136 25378 3148
rect 25869 3145 25881 3148
rect 25915 3145 25927 3179
rect 26602 3176 26608 3188
rect 26563 3148 26608 3176
rect 25869 3139 25927 3145
rect 26602 3136 26608 3148
rect 26660 3136 26666 3188
rect 26786 3136 26792 3188
rect 26844 3176 26850 3188
rect 27341 3179 27399 3185
rect 27341 3176 27353 3179
rect 26844 3148 27353 3176
rect 26844 3136 26850 3148
rect 27341 3145 27353 3148
rect 27387 3145 27399 3179
rect 27341 3139 27399 3145
rect 4433 3111 4491 3117
rect 4433 3077 4445 3111
rect 4479 3108 4491 3111
rect 4982 3108 4988 3120
rect 4479 3080 4988 3108
rect 4479 3077 4491 3080
rect 4433 3071 4491 3077
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 11606 3068 11612 3120
rect 11664 3108 11670 3120
rect 12161 3111 12219 3117
rect 12161 3108 12173 3111
rect 11664 3080 12173 3108
rect 11664 3068 11670 3080
rect 12161 3077 12173 3080
rect 12207 3077 12219 3111
rect 12161 3071 12219 3077
rect 6270 3040 6276 3052
rect 6231 3012 6276 3040
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 3191 2944 3832 2972
rect 5077 2975 5135 2981
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 5077 2941 5089 2975
rect 5123 2972 5135 2975
rect 6288 2972 6316 3000
rect 5123 2944 6316 2972
rect 8021 2975 8079 2981
rect 5123 2941 5135 2944
rect 5077 2935 5135 2941
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8846 2972 8852 2984
rect 8067 2944 8852 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 10137 2975 10195 2981
rect 10137 2941 10149 2975
rect 10183 2972 10195 2975
rect 10226 2972 10232 2984
rect 10183 2944 10232 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 10226 2932 10232 2944
rect 10284 2932 10290 2984
rect 12176 2972 12204 3071
rect 14108 3012 15332 3040
rect 13078 2972 13084 2984
rect 12176 2944 13084 2972
rect 13078 2932 13084 2944
rect 13136 2972 13142 2984
rect 14108 2972 14136 3012
rect 15194 2972 15200 2984
rect 13136 2944 14136 2972
rect 15155 2944 15200 2972
rect 13136 2932 13142 2944
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 15304 2981 15332 3012
rect 15289 2975 15347 2981
rect 15289 2941 15301 2975
rect 15335 2972 15347 2975
rect 15378 2972 15384 2984
rect 15335 2944 15384 2972
rect 15335 2941 15347 2944
rect 15289 2935 15347 2941
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 18233 2975 18291 2981
rect 18233 2972 18245 2975
rect 17644 2944 18245 2972
rect 17644 2932 17650 2944
rect 18233 2941 18245 2944
rect 18279 2972 18291 2975
rect 18785 2975 18843 2981
rect 18785 2972 18797 2975
rect 18279 2944 18797 2972
rect 18279 2941 18291 2944
rect 18233 2935 18291 2941
rect 18785 2941 18797 2944
rect 18831 2941 18843 2975
rect 18785 2935 18843 2941
rect 25130 2932 25136 2984
rect 25188 2972 25194 2984
rect 25317 2975 25375 2981
rect 25317 2972 25329 2975
rect 25188 2944 25329 2972
rect 25188 2932 25194 2944
rect 25317 2941 25329 2944
rect 25363 2941 25375 2975
rect 26418 2972 26424 2984
rect 26379 2944 26424 2972
rect 25317 2935 25375 2941
rect 26418 2932 26424 2944
rect 26476 2972 26482 2984
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26476 2944 26985 2972
rect 26476 2932 26482 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 27522 2972 27528 2984
rect 27483 2944 27528 2972
rect 26973 2935 27031 2941
rect 27522 2932 27528 2944
rect 27580 2972 27586 2984
rect 28077 2975 28135 2981
rect 28077 2972 28089 2975
rect 27580 2944 28089 2972
rect 27580 2932 27586 2944
rect 28077 2941 28089 2944
rect 28123 2941 28135 2975
rect 28077 2935 28135 2941
rect 474 2864 480 2916
rect 532 2904 538 2916
rect 2133 2907 2191 2913
rect 2133 2904 2145 2907
rect 532 2876 2145 2904
rect 532 2864 538 2876
rect 2133 2873 2145 2876
rect 2179 2873 2191 2907
rect 2133 2867 2191 2873
rect 5353 2907 5411 2913
rect 5353 2873 5365 2907
rect 5399 2904 5411 2907
rect 5626 2904 5632 2916
rect 5399 2876 5632 2904
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 5626 2864 5632 2876
rect 5684 2864 5690 2916
rect 8294 2904 8300 2916
rect 8255 2876 8300 2904
rect 8294 2864 8300 2876
rect 8352 2864 8358 2916
rect 10045 2907 10103 2913
rect 10045 2873 10057 2907
rect 10091 2904 10103 2907
rect 10404 2907 10462 2913
rect 10404 2904 10416 2907
rect 10091 2876 10416 2904
rect 10091 2873 10103 2876
rect 10045 2867 10103 2873
rect 10404 2873 10416 2876
rect 10450 2904 10462 2907
rect 10594 2904 10600 2916
rect 10450 2876 10600 2904
rect 10450 2873 10462 2876
rect 10404 2867 10462 2873
rect 10594 2864 10600 2876
rect 10652 2864 10658 2916
rect 12894 2904 12900 2916
rect 12855 2876 12900 2904
rect 12894 2864 12900 2876
rect 12952 2904 12958 2916
rect 13326 2907 13384 2913
rect 13326 2904 13338 2907
rect 12952 2876 13338 2904
rect 12952 2864 12958 2876
rect 13326 2873 13338 2876
rect 13372 2873 13384 2907
rect 15534 2907 15592 2913
rect 15534 2904 15546 2907
rect 13326 2867 13384 2873
rect 14752 2876 15546 2904
rect 3326 2836 3332 2848
rect 3287 2808 3332 2836
rect 3326 2796 3332 2808
rect 3384 2796 3390 2848
rect 10870 2796 10876 2848
rect 10928 2836 10934 2848
rect 11517 2839 11575 2845
rect 11517 2836 11529 2839
rect 10928 2808 11529 2836
rect 10928 2796 10934 2808
rect 11517 2805 11529 2808
rect 11563 2836 11575 2839
rect 11790 2836 11796 2848
rect 11563 2808 11796 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 13814 2796 13820 2848
rect 13872 2836 13878 2848
rect 14752 2845 14780 2876
rect 15534 2873 15546 2876
rect 15580 2873 15592 2907
rect 15534 2867 15592 2873
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 13872 2808 14473 2836
rect 13872 2796 13878 2808
rect 14461 2805 14473 2808
rect 14507 2836 14519 2839
rect 14737 2839 14795 2845
rect 14737 2836 14749 2839
rect 14507 2808 14749 2836
rect 14507 2805 14519 2808
rect 14461 2799 14519 2805
rect 14737 2805 14749 2808
rect 14783 2805 14795 2839
rect 14737 2799 14795 2805
rect 16574 2796 16580 2848
rect 16632 2836 16638 2848
rect 16669 2839 16727 2845
rect 16669 2836 16681 2839
rect 16632 2808 16681 2836
rect 16632 2796 16638 2808
rect 16669 2805 16681 2808
rect 16715 2805 16727 2839
rect 17034 2836 17040 2848
rect 16995 2808 17040 2836
rect 16669 2799 16727 2805
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 18414 2836 18420 2848
rect 18375 2808 18420 2836
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 25498 2836 25504 2848
rect 25459 2808 25504 2836
rect 25498 2796 25504 2808
rect 25556 2796 25562 2848
rect 27706 2836 27712 2848
rect 27667 2808 27712 2836
rect 27706 2796 27712 2808
rect 27764 2796 27770 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 1673 2635 1731 2641
rect 1673 2601 1685 2635
rect 1719 2632 1731 2635
rect 1762 2632 1768 2644
rect 1719 2604 1768 2632
rect 1719 2601 1731 2604
rect 1673 2595 1731 2601
rect 1762 2592 1768 2604
rect 1820 2592 1826 2644
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 3510 2632 3516 2644
rect 2823 2604 3516 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2792 2496 2820 2595
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5868 2604 6009 2632
rect 5868 2592 5874 2604
rect 5997 2601 6009 2604
rect 6043 2601 6055 2635
rect 5997 2595 6055 2601
rect 8297 2635 8355 2641
rect 8297 2601 8309 2635
rect 8343 2632 8355 2635
rect 9582 2632 9588 2644
rect 8343 2604 9588 2632
rect 8343 2601 8355 2604
rect 8297 2595 8355 2601
rect 5442 2564 5448 2576
rect 1995 2468 2820 2496
rect 4448 2536 5448 2564
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2498 2428 2504 2440
rect 2271 2400 2504 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 4448 2428 4476 2536
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 7742 2564 7748 2576
rect 7703 2536 7748 2564
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 4884 2499 4942 2505
rect 4884 2496 4896 2499
rect 4571 2468 4896 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4884 2465 4896 2468
rect 4930 2496 4942 2499
rect 6638 2496 6644 2508
rect 4930 2468 6644 2496
rect 4930 2465 4942 2468
rect 4884 2459 4942 2465
rect 6638 2456 6644 2468
rect 6696 2456 6702 2508
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 8312 2496 8340 2595
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10226 2632 10232 2644
rect 10187 2604 10232 2632
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11606 2632 11612 2644
rect 11567 2604 11612 2632
rect 11606 2592 11612 2604
rect 11664 2592 11670 2644
rect 13814 2632 13820 2644
rect 13775 2604 13820 2632
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17034 2592 17040 2644
rect 17092 2632 17098 2644
rect 17129 2635 17187 2641
rect 17129 2632 17141 2635
rect 17092 2604 17141 2632
rect 17092 2592 17098 2604
rect 17129 2601 17141 2604
rect 17175 2601 17187 2635
rect 19610 2632 19616 2644
rect 19571 2604 19616 2632
rect 17129 2595 17187 2601
rect 19610 2592 19616 2604
rect 19668 2592 19674 2644
rect 23014 2632 23020 2644
rect 22975 2604 23020 2632
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 7515 2468 8340 2496
rect 10321 2499 10379 2505
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 10888 2496 10916 2592
rect 10367 2468 10916 2496
rect 11425 2499 11483 2505
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11471 2468 11989 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11977 2465 11989 2468
rect 12023 2496 12035 2499
rect 12894 2496 12900 2508
rect 12023 2468 12900 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 12894 2456 12900 2468
rect 12952 2456 12958 2508
rect 13173 2499 13231 2505
rect 13173 2465 13185 2499
rect 13219 2496 13231 2499
rect 13832 2496 13860 2592
rect 14921 2567 14979 2573
rect 14921 2533 14933 2567
rect 14967 2564 14979 2567
rect 15289 2567 15347 2573
rect 15289 2564 15301 2567
rect 14967 2536 15301 2564
rect 14967 2533 14979 2536
rect 14921 2527 14979 2533
rect 15289 2533 15301 2536
rect 15335 2564 15347 2567
rect 15740 2567 15798 2573
rect 15740 2564 15752 2567
rect 15335 2536 15752 2564
rect 15335 2533 15347 2536
rect 15289 2527 15347 2533
rect 15740 2533 15752 2536
rect 15786 2564 15798 2567
rect 16482 2564 16488 2576
rect 15786 2536 16488 2564
rect 15786 2533 15798 2536
rect 15740 2527 15798 2533
rect 13219 2468 13860 2496
rect 14277 2499 14335 2505
rect 13219 2465 13231 2468
rect 13173 2459 13231 2465
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14936 2496 14964 2527
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 14323 2468 14964 2496
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15436 2468 15485 2496
rect 15436 2456 15442 2468
rect 15473 2465 15485 2468
rect 15519 2496 15531 2499
rect 17052 2496 17080 2592
rect 15519 2468 17080 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 18138 2456 18144 2508
rect 18196 2496 18202 2508
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18196 2468 18337 2496
rect 18196 2456 18202 2468
rect 18325 2465 18337 2468
rect 18371 2496 18383 2499
rect 18877 2499 18935 2505
rect 18877 2496 18889 2499
rect 18371 2468 18889 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18877 2465 18889 2468
rect 18923 2465 18935 2499
rect 19426 2496 19432 2508
rect 19387 2468 19432 2496
rect 18877 2459 18935 2465
rect 19426 2456 19432 2468
rect 19484 2496 19490 2508
rect 19981 2499 20039 2505
rect 19981 2496 19993 2499
rect 19484 2468 19993 2496
rect 19484 2456 19490 2468
rect 19981 2465 19993 2468
rect 20027 2465 20039 2499
rect 22830 2496 22836 2508
rect 22791 2468 22836 2496
rect 19981 2459 20039 2465
rect 22830 2456 22836 2468
rect 22888 2496 22894 2508
rect 23385 2499 23443 2505
rect 23385 2496 23397 2499
rect 22888 2468 23397 2496
rect 22888 2456 22894 2468
rect 23385 2465 23397 2468
rect 23431 2465 23443 2499
rect 24578 2496 24584 2508
rect 24539 2468 24584 2496
rect 23385 2459 23443 2465
rect 24578 2456 24584 2468
rect 24636 2496 24642 2508
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24636 2468 25145 2496
rect 24636 2456 24642 2468
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25682 2496 25688 2508
rect 25643 2468 25688 2496
rect 25133 2459 25191 2465
rect 25682 2456 25688 2468
rect 25740 2496 25746 2508
rect 26237 2499 26295 2505
rect 26237 2496 26249 2499
rect 25740 2468 26249 2496
rect 25740 2456 25746 2468
rect 26237 2465 26249 2468
rect 26283 2465 26295 2499
rect 26878 2496 26884 2508
rect 26839 2468 26884 2496
rect 26237 2459 26295 2465
rect 26878 2456 26884 2468
rect 26936 2496 26942 2508
rect 27433 2499 27491 2505
rect 27433 2496 27445 2499
rect 26936 2468 27445 2496
rect 26936 2456 26942 2468
rect 27433 2465 27445 2468
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 3927 2400 4629 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 10505 2363 10563 2369
rect 10505 2329 10517 2363
rect 10551 2360 10563 2363
rect 12802 2360 12808 2372
rect 10551 2332 12808 2360
rect 10551 2329 10563 2332
rect 10505 2323 10563 2329
rect 12802 2320 12808 2332
rect 12860 2320 12866 2372
rect 14461 2363 14519 2369
rect 14461 2329 14473 2363
rect 14507 2360 14519 2363
rect 18506 2360 18512 2372
rect 14507 2332 15516 2360
rect 18467 2332 18512 2360
rect 14507 2329 14519 2332
rect 14461 2323 14519 2329
rect 13357 2295 13415 2301
rect 13357 2261 13369 2295
rect 13403 2292 13415 2295
rect 14734 2292 14740 2304
rect 13403 2264 14740 2292
rect 13403 2261 13415 2264
rect 13357 2255 13415 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 15488 2292 15516 2332
rect 18506 2320 18512 2332
rect 18564 2320 18570 2372
rect 15838 2292 15844 2304
rect 15488 2264 15844 2292
rect 15838 2252 15844 2264
rect 15896 2252 15902 2304
rect 24762 2292 24768 2304
rect 24723 2264 24768 2292
rect 24762 2252 24768 2264
rect 24820 2252 24826 2304
rect 25866 2292 25872 2304
rect 25827 2264 25872 2292
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 27062 2292 27068 2304
rect 27023 2264 27068 2292
rect 27062 2252 27068 2264
rect 27120 2252 27126 2304
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 3332 22516 3384 22568
rect 7656 22516 7708 22568
rect 4068 22108 4120 22160
rect 13452 22108 13504 22160
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 3700 21088 3752 21140
rect 6368 21020 6420 21072
rect 25596 21020 25648 21072
rect 3884 20952 3936 21004
rect 15844 20952 15896 21004
rect 19064 20952 19116 21004
rect 19524 20952 19576 21004
rect 21640 20995 21692 21004
rect 21640 20961 21649 20995
rect 21649 20961 21683 20995
rect 21683 20961 21692 20995
rect 21640 20952 21692 20961
rect 8208 20884 8260 20936
rect 5172 20816 5224 20868
rect 3332 20748 3384 20800
rect 5080 20748 5132 20800
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 9588 20544 9640 20596
rect 11336 20544 11388 20596
rect 12716 20544 12768 20596
rect 19432 20544 19484 20596
rect 21640 20587 21692 20596
rect 21640 20553 21649 20587
rect 21649 20553 21683 20587
rect 21683 20553 21692 20587
rect 21640 20544 21692 20553
rect 20536 20519 20588 20528
rect 20536 20485 20545 20519
rect 20545 20485 20579 20519
rect 20579 20485 20588 20519
rect 20536 20476 20588 20485
rect 23848 20519 23900 20528
rect 23848 20485 23857 20519
rect 23857 20485 23891 20519
rect 23891 20485 23900 20519
rect 23848 20476 23900 20485
rect 25136 20408 25188 20460
rect 25872 20408 25924 20460
rect 12716 20340 12768 20392
rect 18052 20383 18104 20392
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 19156 20383 19208 20392
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 23664 20383 23716 20392
rect 19524 20272 19576 20324
rect 20720 20272 20772 20324
rect 21640 20272 21692 20324
rect 22100 20272 22152 20324
rect 23664 20349 23673 20383
rect 23673 20349 23707 20383
rect 23707 20349 23716 20383
rect 23664 20340 23716 20349
rect 9220 20247 9272 20256
rect 9220 20213 9229 20247
rect 9229 20213 9263 20247
rect 9263 20213 9272 20247
rect 9220 20204 9272 20213
rect 13084 20204 13136 20256
rect 16488 20247 16540 20256
rect 16488 20213 16497 20247
rect 16497 20213 16531 20247
rect 16531 20213 16540 20247
rect 16488 20204 16540 20213
rect 18236 20247 18288 20256
rect 18236 20213 18245 20247
rect 18245 20213 18279 20247
rect 18279 20213 18288 20247
rect 18236 20204 18288 20213
rect 19064 20247 19116 20256
rect 19064 20213 19073 20247
rect 19073 20213 19107 20247
rect 19107 20213 19116 20247
rect 19064 20204 19116 20213
rect 19432 20204 19484 20256
rect 22008 20247 22060 20256
rect 22008 20213 22017 20247
rect 22017 20213 22051 20247
rect 22051 20213 22060 20247
rect 22008 20204 22060 20213
rect 22376 20247 22428 20256
rect 22376 20213 22385 20247
rect 22385 20213 22419 20247
rect 22419 20213 22428 20247
rect 22376 20204 22428 20213
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 21548 20000 21600 20052
rect 17316 19907 17368 19916
rect 17316 19873 17325 19907
rect 17325 19873 17359 19907
rect 17359 19873 17368 19907
rect 17316 19864 17368 19873
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 20720 19864 20772 19916
rect 17500 19771 17552 19780
rect 17500 19737 17509 19771
rect 17509 19737 17543 19771
rect 17543 19737 17552 19771
rect 17500 19728 17552 19737
rect 19616 19771 19668 19780
rect 19616 19737 19625 19771
rect 19625 19737 19659 19771
rect 19659 19737 19668 19771
rect 19616 19728 19668 19737
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 17316 19388 17368 19440
rect 19156 19388 19208 19440
rect 15752 19320 15804 19372
rect 16488 19320 16540 19372
rect 17224 19320 17276 19372
rect 17868 19320 17920 19372
rect 18696 19320 18748 19372
rect 19248 19320 19300 19372
rect 19432 19159 19484 19168
rect 19432 19125 19441 19159
rect 19441 19125 19475 19159
rect 19475 19125 19484 19159
rect 19432 19116 19484 19125
rect 19708 19116 19760 19168
rect 20720 19116 20772 19168
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 19340 18708 19392 18760
rect 29368 18708 29420 18760
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 8024 14424 8076 14476
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 7932 14288 7984 14340
rect 7748 14263 7800 14272
rect 7748 14229 7757 14263
rect 7757 14229 7791 14263
rect 7791 14229 7800 14263
rect 7748 14220 7800 14229
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 8024 14059 8076 14068
rect 8024 14025 8033 14059
rect 8033 14025 8067 14059
rect 8067 14025 8076 14059
rect 8024 14016 8076 14025
rect 8208 14016 8260 14068
rect 8300 13880 8352 13932
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 8484 13855 8536 13864
rect 7840 13812 7892 13821
rect 8484 13821 8493 13855
rect 8493 13821 8527 13855
rect 8527 13821 8536 13855
rect 8484 13812 8536 13821
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 7380 13472 7432 13524
rect 7748 13472 7800 13524
rect 7932 13472 7984 13524
rect 8208 13472 8260 13524
rect 8760 13472 8812 13524
rect 8576 13404 8628 13456
rect 1676 13336 1728 13388
rect 2688 13336 2740 13388
rect 7656 13336 7708 13388
rect 8116 13336 8168 13388
rect 9496 13336 9548 13388
rect 10140 13336 10192 13388
rect 11336 13404 11388 13456
rect 11060 13379 11112 13388
rect 11060 13345 11094 13379
rect 11094 13345 11112 13379
rect 11060 13336 11112 13345
rect 12164 13336 12216 13388
rect 2596 13268 2648 13320
rect 8300 13200 8352 13252
rect 12900 13268 12952 13320
rect 1400 13132 1452 13184
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 12164 13175 12216 13184
rect 12164 13141 12173 13175
rect 12173 13141 12207 13175
rect 12207 13141 12216 13175
rect 12164 13132 12216 13141
rect 15108 13132 15160 13184
rect 15292 13132 15344 13184
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 1676 12971 1728 12980
rect 1676 12937 1685 12971
rect 1685 12937 1719 12971
rect 1719 12937 1728 12971
rect 1676 12928 1728 12937
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 8760 12928 8812 12980
rect 12164 12928 12216 12980
rect 15108 12971 15160 12980
rect 15108 12937 15117 12971
rect 15117 12937 15151 12971
rect 15151 12937 15160 12971
rect 15108 12928 15160 12937
rect 3516 12792 3568 12844
rect 7104 12792 7156 12844
rect 7564 12835 7616 12844
rect 7564 12801 7573 12835
rect 7573 12801 7607 12835
rect 7607 12801 7616 12835
rect 7564 12792 7616 12801
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 7380 12767 7432 12776
rect 7380 12733 7389 12767
rect 7389 12733 7423 12767
rect 7423 12733 7432 12767
rect 7380 12724 7432 12733
rect 2136 12699 2188 12708
rect 2136 12665 2145 12699
rect 2145 12665 2179 12699
rect 2179 12665 2188 12699
rect 2688 12699 2740 12708
rect 2136 12656 2188 12665
rect 2688 12665 2697 12699
rect 2697 12665 2731 12699
rect 2731 12665 2740 12699
rect 2688 12656 2740 12665
rect 10140 12835 10192 12844
rect 10140 12801 10149 12835
rect 10149 12801 10183 12835
rect 10183 12801 10192 12835
rect 10140 12792 10192 12801
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 14464 12792 14516 12844
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 8576 12724 8628 12776
rect 15200 12724 15252 12776
rect 16396 12724 16448 12776
rect 9128 12656 9180 12708
rect 9588 12656 9640 12708
rect 10324 12656 10376 12708
rect 11060 12656 11112 12708
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 5540 12631 5592 12640
rect 5540 12597 5549 12631
rect 5549 12597 5583 12631
rect 5583 12597 5592 12631
rect 5540 12588 5592 12597
rect 7196 12588 7248 12640
rect 9036 12631 9088 12640
rect 9036 12597 9045 12631
rect 9045 12597 9079 12631
rect 9079 12597 9088 12631
rect 9036 12588 9088 12597
rect 10876 12588 10928 12640
rect 13636 12631 13688 12640
rect 13636 12597 13645 12631
rect 13645 12597 13679 12631
rect 13679 12597 13688 12631
rect 13636 12588 13688 12597
rect 15200 12588 15252 12640
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 2780 12427 2832 12436
rect 2780 12393 2789 12427
rect 2789 12393 2823 12427
rect 2823 12393 2832 12427
rect 2780 12384 2832 12393
rect 6276 12384 6328 12436
rect 7104 12427 7156 12436
rect 7104 12393 7113 12427
rect 7113 12393 7147 12427
rect 7147 12393 7156 12427
rect 7104 12384 7156 12393
rect 8300 12384 8352 12436
rect 8576 12384 8628 12436
rect 10876 12427 10928 12436
rect 10876 12393 10885 12427
rect 10885 12393 10919 12427
rect 10919 12393 10928 12427
rect 10876 12384 10928 12393
rect 11336 12384 11388 12436
rect 15200 12384 15252 12436
rect 16396 12384 16448 12436
rect 4896 12316 4948 12368
rect 5540 12316 5592 12368
rect 2872 12248 2924 12300
rect 3056 12248 3108 12300
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 13452 12316 13504 12368
rect 3516 12180 3568 12232
rect 4160 12180 4212 12232
rect 4712 12180 4764 12232
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 10324 12248 10376 12300
rect 16764 12248 16816 12300
rect 17684 12248 17736 12300
rect 13176 12180 13228 12232
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 14464 12180 14516 12232
rect 17500 12180 17552 12232
rect 18604 12180 18656 12232
rect 9036 12155 9088 12164
rect 9036 12121 9045 12155
rect 9045 12121 9079 12155
rect 9079 12121 9088 12155
rect 9036 12112 9088 12121
rect 2412 12044 2464 12096
rect 6276 12087 6328 12096
rect 6276 12053 6285 12087
rect 6285 12053 6319 12087
rect 6319 12053 6328 12087
rect 6276 12044 6328 12053
rect 11336 12044 11388 12096
rect 12900 12044 12952 12096
rect 13544 12044 13596 12096
rect 13728 12044 13780 12096
rect 16856 12044 16908 12096
rect 17408 12087 17460 12096
rect 17408 12053 17417 12087
rect 17417 12053 17451 12087
rect 17451 12053 17460 12087
rect 17408 12044 17460 12053
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 2044 11840 2096 11892
rect 2780 11840 2832 11892
rect 4712 11840 4764 11892
rect 4896 11815 4948 11824
rect 4896 11781 4905 11815
rect 4905 11781 4939 11815
rect 4939 11781 4948 11815
rect 4896 11772 4948 11781
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 2596 11747 2648 11756
rect 2596 11713 2605 11747
rect 2605 11713 2639 11747
rect 2639 11713 2648 11747
rect 2596 11704 2648 11713
rect 10140 11840 10192 11892
rect 13176 11883 13228 11892
rect 13176 11849 13185 11883
rect 13185 11849 13219 11883
rect 13219 11849 13228 11883
rect 13176 11840 13228 11849
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 13544 11840 13596 11892
rect 15292 11883 15344 11892
rect 10416 11772 10468 11824
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 10324 11747 10376 11756
rect 2228 11636 2280 11688
rect 4620 11568 4672 11620
rect 6276 11568 6328 11620
rect 1952 11543 2004 11552
rect 1952 11509 1961 11543
rect 1961 11509 1995 11543
rect 1995 11509 2004 11543
rect 1952 11500 2004 11509
rect 3056 11543 3108 11552
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3056 11500 3108 11509
rect 3516 11500 3568 11552
rect 7472 11500 7524 11552
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 15292 11849 15301 11883
rect 15301 11849 15335 11883
rect 15335 11849 15344 11883
rect 15292 11840 15344 11849
rect 16672 11840 16724 11892
rect 16948 11840 17000 11892
rect 17684 11840 17736 11892
rect 19064 11883 19116 11892
rect 19064 11849 19073 11883
rect 19073 11849 19107 11883
rect 19107 11849 19116 11883
rect 19064 11840 19116 11849
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 17684 11704 17736 11756
rect 18604 11747 18656 11756
rect 9128 11500 9180 11552
rect 10232 11636 10284 11688
rect 17408 11636 17460 11688
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 26424 11679 26476 11688
rect 26424 11645 26433 11679
rect 26433 11645 26467 11679
rect 26467 11645 26476 11679
rect 26424 11636 26476 11645
rect 9680 11611 9732 11620
rect 9680 11577 9689 11611
rect 9689 11577 9723 11611
rect 9723 11577 9732 11611
rect 9680 11568 9732 11577
rect 14464 11568 14516 11620
rect 16856 11611 16908 11620
rect 16856 11577 16865 11611
rect 16865 11577 16899 11611
rect 16899 11577 16908 11611
rect 16856 11568 16908 11577
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 10232 11543 10284 11552
rect 10232 11509 10241 11543
rect 10241 11509 10275 11543
rect 10275 11509 10284 11543
rect 10232 11500 10284 11509
rect 15108 11500 15160 11552
rect 15292 11500 15344 11552
rect 15660 11500 15712 11552
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 18420 11543 18472 11552
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 18420 11500 18472 11509
rect 26608 11543 26660 11552
rect 26608 11509 26617 11543
rect 26617 11509 26651 11543
rect 26651 11509 26660 11543
rect 26608 11500 26660 11509
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 4436 11296 4488 11348
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 8300 11296 8352 11348
rect 10048 11296 10100 11348
rect 2596 11228 2648 11280
rect 2320 11160 2372 11212
rect 4344 11160 4396 11212
rect 9956 11228 10008 11280
rect 10508 11228 10560 11280
rect 7380 11203 7432 11212
rect 7380 11169 7389 11203
rect 7389 11169 7423 11203
rect 7423 11169 7432 11203
rect 7380 11160 7432 11169
rect 7472 11160 7524 11212
rect 10784 11296 10836 11348
rect 13636 11296 13688 11348
rect 16304 11296 16356 11348
rect 15476 11228 15528 11280
rect 15660 11228 15712 11280
rect 17960 11228 18012 11280
rect 18420 11228 18472 11280
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 2780 11024 2832 11076
rect 2872 10956 2924 11008
rect 3332 10956 3384 11008
rect 8944 10956 8996 11008
rect 9404 10956 9456 11008
rect 13728 11160 13780 11212
rect 14464 11203 14516 11212
rect 14464 11169 14473 11203
rect 14473 11169 14507 11203
rect 14507 11169 14516 11203
rect 17684 11203 17736 11212
rect 14464 11160 14516 11169
rect 17684 11169 17693 11203
rect 17693 11169 17727 11203
rect 17727 11169 17736 11203
rect 17684 11160 17736 11169
rect 21916 11160 21968 11212
rect 27344 11160 27396 11212
rect 9680 11092 9732 11144
rect 10140 11024 10192 11076
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 13084 11092 13136 11144
rect 15108 11092 15160 11144
rect 15844 11092 15896 11144
rect 16672 11092 16724 11144
rect 17500 11092 17552 11144
rect 17868 11092 17920 11144
rect 18604 11092 18656 11144
rect 10508 11024 10560 11076
rect 11520 11024 11572 11076
rect 16580 11024 16632 11076
rect 26700 11067 26752 11076
rect 26700 11033 26709 11067
rect 26709 11033 26743 11067
rect 26743 11033 26752 11067
rect 26700 11024 26752 11033
rect 13728 10956 13780 11008
rect 15752 10999 15804 11008
rect 15752 10965 15761 10999
rect 15761 10965 15795 10999
rect 15795 10965 15804 10999
rect 15752 10956 15804 10965
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 2596 10752 2648 10804
rect 2872 10795 2924 10804
rect 2872 10761 2881 10795
rect 2881 10761 2915 10795
rect 2915 10761 2924 10795
rect 2872 10752 2924 10761
rect 4620 10752 4672 10804
rect 7472 10795 7524 10804
rect 7472 10761 7481 10795
rect 7481 10761 7515 10795
rect 7515 10761 7524 10795
rect 7472 10752 7524 10761
rect 8944 10795 8996 10804
rect 8944 10761 8953 10795
rect 8953 10761 8987 10795
rect 8987 10761 8996 10795
rect 8944 10752 8996 10761
rect 9680 10795 9732 10804
rect 9680 10761 9689 10795
rect 9689 10761 9723 10795
rect 9723 10761 9732 10795
rect 9680 10752 9732 10761
rect 10048 10752 10100 10804
rect 13820 10752 13872 10804
rect 15200 10795 15252 10804
rect 15200 10761 15209 10795
rect 15209 10761 15243 10795
rect 15243 10761 15252 10795
rect 15200 10752 15252 10761
rect 17868 10752 17920 10804
rect 27344 10795 27396 10804
rect 27344 10761 27353 10795
rect 27353 10761 27387 10795
rect 27387 10761 27396 10795
rect 27344 10752 27396 10761
rect 4436 10727 4488 10736
rect 4436 10693 4445 10727
rect 4445 10693 4479 10727
rect 4479 10693 4488 10727
rect 4436 10684 4488 10693
rect 7380 10684 7432 10736
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 3516 10659 3568 10668
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 4344 10616 4396 10668
rect 10324 10659 10376 10668
rect 10324 10625 10333 10659
rect 10333 10625 10367 10659
rect 10367 10625 10376 10659
rect 10324 10616 10376 10625
rect 14372 10616 14424 10668
rect 3424 10480 3476 10532
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 9128 10412 9180 10464
rect 11336 10548 11388 10600
rect 15660 10548 15712 10600
rect 15752 10548 15804 10600
rect 16396 10548 16448 10600
rect 26424 10591 26476 10600
rect 26424 10557 26433 10591
rect 26433 10557 26467 10591
rect 26467 10557 26476 10591
rect 26424 10548 26476 10557
rect 13452 10480 13504 10532
rect 10140 10455 10192 10464
rect 10140 10421 10149 10455
rect 10149 10421 10183 10455
rect 10183 10421 10192 10455
rect 10140 10412 10192 10421
rect 13084 10412 13136 10464
rect 13176 10412 13228 10464
rect 13728 10455 13780 10464
rect 13728 10421 13737 10455
rect 13737 10421 13771 10455
rect 13771 10421 13780 10455
rect 13728 10412 13780 10421
rect 17500 10412 17552 10464
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 26608 10455 26660 10464
rect 26608 10421 26617 10455
rect 26617 10421 26651 10455
rect 26651 10421 26660 10455
rect 26608 10412 26660 10421
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 6092 10251 6144 10260
rect 6092 10217 6101 10251
rect 6101 10217 6135 10251
rect 6135 10217 6144 10251
rect 6092 10208 6144 10217
rect 6828 10208 6880 10260
rect 7380 10208 7432 10260
rect 7840 10208 7892 10260
rect 9680 10251 9732 10260
rect 9680 10217 9689 10251
rect 9689 10217 9723 10251
rect 9723 10217 9732 10251
rect 9680 10208 9732 10217
rect 9772 10208 9824 10260
rect 10416 10208 10468 10260
rect 13728 10208 13780 10260
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 15752 10208 15804 10260
rect 2872 10140 2924 10192
rect 2964 10140 3016 10192
rect 15844 10183 15896 10192
rect 15844 10149 15853 10183
rect 15853 10149 15887 10183
rect 15887 10149 15896 10183
rect 15844 10140 15896 10149
rect 16304 10140 16356 10192
rect 2504 10072 2556 10124
rect 5448 10072 5500 10124
rect 6920 10072 6972 10124
rect 9864 10072 9916 10124
rect 12900 10072 12952 10124
rect 13084 10072 13136 10124
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 2780 10004 2832 10013
rect 2412 9936 2464 9988
rect 3516 10004 3568 10056
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 4896 9868 4948 9920
rect 8300 9868 8352 9920
rect 9312 9868 9364 9920
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 3424 9664 3476 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 2136 9596 2188 9648
rect 2780 9596 2832 9648
rect 4712 9664 4764 9716
rect 6828 9664 6880 9716
rect 10416 9707 10468 9716
rect 10416 9673 10425 9707
rect 10425 9673 10459 9707
rect 10459 9673 10468 9707
rect 10416 9664 10468 9673
rect 13084 9707 13136 9716
rect 13084 9673 13093 9707
rect 13093 9673 13127 9707
rect 13127 9673 13136 9707
rect 13084 9664 13136 9673
rect 13452 9707 13504 9716
rect 13452 9673 13461 9707
rect 13461 9673 13495 9707
rect 13495 9673 13504 9707
rect 13452 9664 13504 9673
rect 14372 9664 14424 9716
rect 10324 9596 10376 9648
rect 3792 9528 3844 9580
rect 5448 9528 5500 9580
rect 8300 9528 8352 9580
rect 4160 9460 4212 9512
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 12072 9528 12124 9580
rect 12900 9528 12952 9580
rect 13452 9528 13504 9580
rect 10324 9460 10376 9512
rect 11796 9460 11848 9512
rect 3700 9392 3752 9444
rect 8392 9435 8444 9444
rect 8392 9401 8401 9435
rect 8401 9401 8435 9435
rect 8435 9401 8444 9435
rect 8392 9392 8444 9401
rect 14372 9392 14424 9444
rect 2504 9324 2556 9376
rect 3056 9324 3108 9376
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 4988 9324 5040 9376
rect 5448 9324 5500 9376
rect 6920 9324 6972 9376
rect 8484 9324 8536 9376
rect 8944 9367 8996 9376
rect 8944 9333 8953 9367
rect 8953 9333 8987 9367
rect 8987 9333 8996 9367
rect 8944 9324 8996 9333
rect 9864 9324 9916 9376
rect 12072 9367 12124 9376
rect 12072 9333 12081 9367
rect 12081 9333 12115 9367
rect 12115 9333 12124 9367
rect 12072 9324 12124 9333
rect 15568 9367 15620 9376
rect 15568 9333 15577 9367
rect 15577 9333 15611 9367
rect 15611 9333 15620 9367
rect 15568 9324 15620 9333
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 1400 9120 1452 9172
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 3332 9120 3384 9172
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 8484 9163 8536 9172
rect 8484 9129 8493 9163
rect 8493 9129 8527 9163
rect 8527 9129 8536 9163
rect 8484 9120 8536 9129
rect 13452 9163 13504 9172
rect 3792 9052 3844 9104
rect 7472 9052 7524 9104
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 26700 9163 26752 9172
rect 26700 9129 26709 9163
rect 26709 9129 26743 9163
rect 26743 9129 26752 9163
rect 26700 9120 26752 9129
rect 2320 8984 2372 9036
rect 4436 9027 4488 9036
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 12072 9052 12124 9104
rect 11612 9027 11664 9036
rect 11612 8993 11646 9027
rect 11646 8993 11664 9027
rect 11612 8984 11664 8993
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 5448 8916 5500 8968
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 8116 8916 8168 8968
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 9036 8916 9088 8968
rect 9956 8916 10008 8968
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 13084 8891 13136 8900
rect 13084 8857 13093 8891
rect 13093 8857 13127 8891
rect 13127 8857 13136 8891
rect 13084 8848 13136 8857
rect 3056 8823 3108 8832
rect 3056 8789 3065 8823
rect 3065 8789 3099 8823
rect 3099 8789 3108 8823
rect 3056 8780 3108 8789
rect 4896 8780 4948 8832
rect 5540 8780 5592 8832
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 9220 8823 9272 8832
rect 9220 8789 9229 8823
rect 9229 8789 9263 8823
rect 9263 8789 9272 8823
rect 9220 8780 9272 8789
rect 12716 8823 12768 8832
rect 12716 8789 12725 8823
rect 12725 8789 12759 8823
rect 12759 8789 12768 8823
rect 12716 8780 12768 8789
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 1492 8576 1544 8628
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 3148 8619 3200 8628
rect 3148 8585 3157 8619
rect 3157 8585 3191 8619
rect 3191 8585 3200 8619
rect 3148 8576 3200 8585
rect 3792 8619 3844 8628
rect 3792 8585 3801 8619
rect 3801 8585 3835 8619
rect 3835 8585 3844 8619
rect 3792 8576 3844 8585
rect 4528 8576 4580 8628
rect 7472 8619 7524 8628
rect 7472 8585 7481 8619
rect 7481 8585 7515 8619
rect 7515 8585 7524 8619
rect 7472 8576 7524 8585
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 8484 8619 8536 8628
rect 8484 8585 8493 8619
rect 8493 8585 8527 8619
rect 8527 8585 8536 8619
rect 8484 8576 8536 8585
rect 11336 8576 11388 8628
rect 26516 8576 26568 8628
rect 2688 8551 2740 8560
rect 2688 8517 2697 8551
rect 2697 8517 2731 8551
rect 2731 8517 2740 8551
rect 2688 8508 2740 8517
rect 6920 8508 6972 8560
rect 26608 8551 26660 8560
rect 26608 8517 26617 8551
rect 26617 8517 26651 8551
rect 26651 8517 26660 8551
rect 26608 8508 26660 8517
rect 27712 8551 27764 8560
rect 27712 8517 27721 8551
rect 27721 8517 27755 8551
rect 27755 8517 27764 8551
rect 27712 8508 27764 8517
rect 3148 8372 3200 8424
rect 5724 8372 5776 8424
rect 4436 8347 4488 8356
rect 4436 8313 4445 8347
rect 4445 8313 4479 8347
rect 4479 8313 4488 8347
rect 4436 8304 4488 8313
rect 4896 8304 4948 8356
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 8208 8440 8260 8492
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 11612 8440 11664 8492
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 7656 8372 7708 8424
rect 13084 8415 13136 8424
rect 8668 8304 8720 8356
rect 9220 8347 9272 8356
rect 9220 8313 9229 8347
rect 9229 8313 9263 8347
rect 9263 8313 9272 8347
rect 9220 8304 9272 8313
rect 13084 8381 13093 8415
rect 13093 8381 13127 8415
rect 13127 8381 13136 8415
rect 13084 8372 13136 8381
rect 26424 8415 26476 8424
rect 26424 8381 26433 8415
rect 26433 8381 26467 8415
rect 26467 8381 26476 8415
rect 26424 8372 26476 8381
rect 27528 8415 27580 8424
rect 27528 8381 27537 8415
rect 27537 8381 27571 8415
rect 27571 8381 27580 8415
rect 27528 8372 27580 8381
rect 6920 8236 6972 8288
rect 12348 8304 12400 8356
rect 11336 8236 11388 8288
rect 11612 8236 11664 8288
rect 12808 8236 12860 8288
rect 16304 8236 16356 8288
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 5448 8075 5500 8084
rect 5448 8041 5457 8075
rect 5457 8041 5491 8075
rect 5491 8041 5500 8075
rect 5448 8032 5500 8041
rect 5632 8032 5684 8084
rect 7012 8032 7064 8084
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 10048 8032 10100 8084
rect 11520 8032 11572 8084
rect 12072 8075 12124 8084
rect 12072 8041 12081 8075
rect 12081 8041 12115 8075
rect 12115 8041 12124 8075
rect 12072 8032 12124 8041
rect 6368 7964 6420 8016
rect 2412 7896 2464 7948
rect 4160 7896 4212 7948
rect 8760 7896 8812 7948
rect 3976 7828 4028 7880
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 7840 7828 7892 7880
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 11612 7871 11664 7880
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 10324 7803 10376 7812
rect 10324 7769 10333 7803
rect 10333 7769 10367 7803
rect 10367 7769 10376 7803
rect 10324 7760 10376 7769
rect 10876 7760 10928 7812
rect 12716 8032 12768 8084
rect 12992 8032 13044 8084
rect 15384 8032 15436 8084
rect 15568 8032 15620 8084
rect 16396 8032 16448 8084
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 13084 7896 13136 7948
rect 13452 7896 13504 7948
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 15844 7828 15896 7880
rect 16672 7828 16724 7880
rect 12992 7760 13044 7812
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 12716 7735 12768 7744
rect 12716 7701 12725 7735
rect 12725 7701 12759 7735
rect 12759 7701 12768 7735
rect 12716 7692 12768 7701
rect 15752 7692 15804 7744
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 2412 7531 2464 7540
rect 2412 7497 2421 7531
rect 2421 7497 2455 7531
rect 2455 7497 2464 7531
rect 2412 7488 2464 7497
rect 6368 7531 6420 7540
rect 6368 7497 6377 7531
rect 6377 7497 6411 7531
rect 6411 7497 6420 7531
rect 6368 7488 6420 7497
rect 7012 7531 7064 7540
rect 7012 7497 7021 7531
rect 7021 7497 7055 7531
rect 7055 7497 7064 7531
rect 7012 7488 7064 7497
rect 7840 7531 7892 7540
rect 7840 7497 7849 7531
rect 7849 7497 7883 7531
rect 7883 7497 7892 7531
rect 7840 7488 7892 7497
rect 8576 7531 8628 7540
rect 8576 7497 8585 7531
rect 8585 7497 8619 7531
rect 8619 7497 8628 7531
rect 8576 7488 8628 7497
rect 11428 7488 11480 7540
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 15108 7531 15160 7540
rect 15108 7497 15117 7531
rect 15117 7497 15151 7531
rect 15151 7497 15160 7531
rect 15108 7488 15160 7497
rect 15844 7488 15896 7540
rect 26516 7488 26568 7540
rect 1584 7463 1636 7472
rect 1584 7429 1593 7463
rect 1593 7429 1627 7463
rect 1627 7429 1636 7463
rect 1584 7420 1636 7429
rect 2964 7395 3016 7404
rect 2964 7361 2973 7395
rect 2973 7361 3007 7395
rect 3007 7361 3016 7395
rect 2964 7352 3016 7361
rect 4712 7352 4764 7404
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 8760 7420 8812 7472
rect 12256 7420 12308 7472
rect 9496 7352 9548 7404
rect 10692 7395 10744 7404
rect 10692 7361 10701 7395
rect 10701 7361 10735 7395
rect 10735 7361 10744 7395
rect 10692 7352 10744 7361
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 12716 7352 12768 7404
rect 5632 7284 5684 7336
rect 6276 7284 6328 7336
rect 8760 7284 8812 7336
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 10600 7327 10652 7336
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 10600 7284 10652 7293
rect 11336 7284 11388 7336
rect 11888 7284 11940 7336
rect 12808 7327 12860 7336
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 15568 7420 15620 7472
rect 18144 7420 18196 7472
rect 12992 7352 13044 7361
rect 16672 7352 16724 7404
rect 16304 7327 16356 7336
rect 16304 7293 16313 7327
rect 16313 7293 16347 7327
rect 16347 7293 16356 7327
rect 16304 7284 16356 7293
rect 26424 7327 26476 7336
rect 26424 7293 26433 7327
rect 26433 7293 26467 7327
rect 26467 7293 26476 7327
rect 26424 7284 26476 7293
rect 9036 7259 9088 7268
rect 9036 7225 9045 7259
rect 9045 7225 9079 7259
rect 9079 7225 9088 7259
rect 9036 7216 9088 7225
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 4160 7148 4212 7200
rect 5080 7148 5132 7200
rect 5264 7148 5316 7200
rect 6460 7148 6512 7200
rect 6920 7148 6972 7200
rect 8944 7148 8996 7200
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 11520 7148 11572 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 13452 7191 13504 7200
rect 12440 7148 12492 7157
rect 13452 7157 13461 7191
rect 13461 7157 13495 7191
rect 13495 7157 13504 7191
rect 13452 7148 13504 7157
rect 15936 7191 15988 7200
rect 15936 7157 15945 7191
rect 15945 7157 15979 7191
rect 15979 7157 15988 7191
rect 15936 7148 15988 7157
rect 16672 7148 16724 7200
rect 26608 7191 26660 7200
rect 26608 7157 26617 7191
rect 26617 7157 26651 7191
rect 26651 7157 26660 7191
rect 26608 7148 26660 7157
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 3976 6944 4028 6996
rect 5632 6987 5684 6996
rect 5632 6953 5641 6987
rect 5641 6953 5675 6987
rect 5675 6953 5684 6987
rect 5632 6944 5684 6953
rect 9036 6987 9088 6996
rect 9036 6953 9045 6987
rect 9045 6953 9079 6987
rect 9079 6953 9088 6987
rect 9036 6944 9088 6953
rect 10140 6944 10192 6996
rect 11612 6944 11664 6996
rect 11888 6987 11940 6996
rect 11888 6953 11897 6987
rect 11897 6953 11931 6987
rect 11931 6953 11940 6987
rect 11888 6944 11940 6953
rect 12900 6944 12952 6996
rect 13360 6944 13412 6996
rect 15936 6944 15988 6996
rect 16304 6987 16356 6996
rect 16304 6953 16313 6987
rect 16313 6953 16347 6987
rect 16347 6953 16356 6987
rect 16304 6944 16356 6953
rect 2596 6876 2648 6928
rect 3240 6876 3292 6928
rect 1952 6808 2004 6860
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2504 6808 2556 6817
rect 3424 6808 3476 6860
rect 5080 6876 5132 6928
rect 5816 6876 5868 6928
rect 5172 6851 5224 6860
rect 5172 6817 5181 6851
rect 5181 6817 5215 6851
rect 5215 6817 5224 6851
rect 5172 6808 5224 6817
rect 6276 6808 6328 6860
rect 6460 6808 6512 6860
rect 8944 6876 8996 6928
rect 15752 6919 15804 6928
rect 6368 6783 6420 6792
rect 1584 6715 1636 6724
rect 1584 6681 1593 6715
rect 1593 6681 1627 6715
rect 1627 6681 1636 6715
rect 1584 6672 1636 6681
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 9128 6808 9180 6860
rect 15752 6885 15761 6919
rect 15761 6885 15795 6919
rect 15795 6885 15804 6919
rect 15752 6876 15804 6885
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 15476 6740 15528 6792
rect 26700 6715 26752 6724
rect 26700 6681 26709 6715
rect 26709 6681 26743 6715
rect 26743 6681 26752 6715
rect 26700 6672 26752 6681
rect 2688 6647 2740 6656
rect 2688 6613 2697 6647
rect 2697 6613 2731 6647
rect 2731 6613 2740 6647
rect 2688 6604 2740 6613
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 13636 6604 13688 6656
rect 15200 6604 15252 6656
rect 16672 6647 16724 6656
rect 16672 6613 16681 6647
rect 16681 6613 16715 6647
rect 16715 6613 16724 6647
rect 16672 6604 16724 6613
rect 17040 6647 17092 6656
rect 17040 6613 17049 6647
rect 17049 6613 17083 6647
rect 17083 6613 17092 6647
rect 17040 6604 17092 6613
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 1952 6443 2004 6452
rect 1952 6409 1961 6443
rect 1961 6409 1995 6443
rect 1995 6409 2004 6443
rect 1952 6400 2004 6409
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 6276 6400 6328 6452
rect 6828 6400 6880 6452
rect 8576 6400 8628 6452
rect 10324 6443 10376 6452
rect 6368 6332 6420 6384
rect 4068 6264 4120 6316
rect 2136 6196 2188 6248
rect 3424 6239 3476 6248
rect 3424 6205 3433 6239
rect 3433 6205 3467 6239
rect 3467 6205 3476 6239
rect 3424 6196 3476 6205
rect 10324 6409 10333 6443
rect 10333 6409 10367 6443
rect 10367 6409 10376 6443
rect 10324 6400 10376 6409
rect 15476 6443 15528 6452
rect 15476 6409 15485 6443
rect 15485 6409 15519 6443
rect 15519 6409 15528 6443
rect 15476 6400 15528 6409
rect 10140 6332 10192 6384
rect 8944 6239 8996 6248
rect 8944 6205 8953 6239
rect 8953 6205 8987 6239
rect 8987 6205 8996 6239
rect 8944 6196 8996 6205
rect 10232 6264 10284 6316
rect 13636 6264 13688 6316
rect 16028 6264 16080 6316
rect 16672 6264 16724 6316
rect 11796 6196 11848 6248
rect 16488 6196 16540 6248
rect 17040 6196 17092 6248
rect 26516 6239 26568 6248
rect 26516 6205 26525 6239
rect 26525 6205 26559 6239
rect 26559 6205 26568 6239
rect 26516 6196 26568 6205
rect 13912 6128 13964 6180
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 2688 6060 2740 6112
rect 3516 6103 3568 6112
rect 3516 6069 3525 6103
rect 3525 6069 3559 6103
rect 3559 6069 3568 6103
rect 3516 6060 3568 6069
rect 5540 6060 5592 6112
rect 6460 6060 6512 6112
rect 6828 6060 6880 6112
rect 12440 6060 12492 6112
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 16304 6060 16356 6112
rect 16856 6060 16908 6112
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 2136 5856 2188 5908
rect 3516 5856 3568 5908
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 10324 5856 10376 5908
rect 13912 5899 13964 5908
rect 13912 5865 13921 5899
rect 13921 5865 13955 5899
rect 13955 5865 13964 5899
rect 13912 5856 13964 5865
rect 15752 5856 15804 5908
rect 16856 5899 16908 5908
rect 16856 5865 16865 5899
rect 16865 5865 16899 5899
rect 16899 5865 16908 5899
rect 16856 5856 16908 5865
rect 17592 5856 17644 5908
rect 26700 5899 26752 5908
rect 26700 5865 26709 5899
rect 26709 5865 26743 5899
rect 26743 5865 26752 5899
rect 26700 5856 26752 5865
rect 6000 5831 6052 5840
rect 6000 5797 6009 5831
rect 6009 5797 6043 5831
rect 6043 5797 6052 5831
rect 6000 5788 6052 5797
rect 6552 5788 6604 5840
rect 12532 5788 12584 5840
rect 2412 5720 2464 5772
rect 4344 5720 4396 5772
rect 10416 5720 10468 5772
rect 12440 5720 12492 5772
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4528 5652 4580 5661
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 13084 5720 13136 5772
rect 15384 5720 15436 5772
rect 16028 5788 16080 5840
rect 17224 5763 17276 5772
rect 17224 5729 17233 5763
rect 17233 5729 17267 5763
rect 17267 5729 17276 5763
rect 17224 5720 17276 5729
rect 26516 5763 26568 5772
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 4068 5584 4120 5636
rect 16212 5584 16264 5636
rect 16948 5584 17000 5636
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 4804 5516 4856 5568
rect 12532 5516 12584 5568
rect 13636 5516 13688 5568
rect 15292 5559 15344 5568
rect 15292 5525 15301 5559
rect 15301 5525 15335 5559
rect 15335 5525 15344 5559
rect 15292 5516 15344 5525
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 2412 5355 2464 5364
rect 2412 5321 2421 5355
rect 2421 5321 2455 5355
rect 2455 5321 2464 5355
rect 2412 5312 2464 5321
rect 4068 5312 4120 5364
rect 4344 5355 4396 5364
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 5724 5355 5776 5364
rect 5724 5321 5733 5355
rect 5733 5321 5767 5355
rect 5767 5321 5776 5355
rect 5724 5312 5776 5321
rect 6276 5312 6328 5364
rect 10324 5355 10376 5364
rect 10324 5321 10333 5355
rect 10333 5321 10367 5355
rect 10367 5321 10376 5355
rect 10324 5312 10376 5321
rect 10416 5312 10468 5364
rect 12532 5312 12584 5364
rect 15844 5312 15896 5364
rect 16488 5312 16540 5364
rect 17224 5312 17276 5364
rect 17868 5312 17920 5364
rect 26608 5355 26660 5364
rect 26608 5321 26617 5355
rect 26617 5321 26651 5355
rect 26651 5321 26660 5355
rect 26608 5312 26660 5321
rect 5540 5244 5592 5296
rect 6552 5244 6604 5296
rect 16580 5244 16632 5296
rect 17592 5244 17644 5296
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 16948 5219 17000 5228
rect 4712 5151 4764 5160
rect 4712 5117 4721 5151
rect 4721 5117 4755 5151
rect 4755 5117 4764 5151
rect 4712 5108 4764 5117
rect 13636 5151 13688 5160
rect 13636 5117 13645 5151
rect 13645 5117 13679 5151
rect 13679 5117 13688 5151
rect 13636 5108 13688 5117
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 15476 5108 15528 5160
rect 16212 5108 16264 5160
rect 16764 5151 16816 5160
rect 16764 5117 16773 5151
rect 16773 5117 16807 5151
rect 16807 5117 16816 5151
rect 16764 5108 16816 5117
rect 16580 5040 16632 5092
rect 18144 5040 18196 5092
rect 26516 5108 26568 5160
rect 1400 4972 1452 5024
rect 2044 5015 2096 5024
rect 2044 4981 2053 5015
rect 2053 4981 2087 5015
rect 2087 4981 2096 5015
rect 2044 4972 2096 4981
rect 13084 5015 13136 5024
rect 13084 4981 13093 5015
rect 13093 4981 13127 5015
rect 13127 4981 13136 5015
rect 13084 4972 13136 4981
rect 14280 4972 14332 5024
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 15384 4972 15436 4981
rect 26332 5015 26384 5024
rect 26332 4981 26341 5015
rect 26341 4981 26375 5015
rect 26375 4981 26384 5015
rect 26332 4972 26384 4981
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 2320 4768 2372 4820
rect 4528 4768 4580 4820
rect 6920 4768 6972 4820
rect 10232 4811 10284 4820
rect 10232 4777 10241 4811
rect 10241 4777 10275 4811
rect 10275 4777 10284 4811
rect 10232 4768 10284 4777
rect 10416 4768 10468 4820
rect 13728 4768 13780 4820
rect 15108 4768 15160 4820
rect 15752 4768 15804 4820
rect 17132 4811 17184 4820
rect 17132 4777 17141 4811
rect 17141 4777 17175 4811
rect 17175 4777 17184 4811
rect 17132 4768 17184 4777
rect 19892 4768 19944 4820
rect 20076 4768 20128 4820
rect 26700 4811 26752 4820
rect 26700 4777 26709 4811
rect 26709 4777 26743 4811
rect 26743 4777 26752 4811
rect 26700 4768 26752 4777
rect 4712 4700 4764 4752
rect 6276 4743 6328 4752
rect 6276 4709 6310 4743
rect 6310 4709 6328 4743
rect 6276 4700 6328 4709
rect 6368 4700 6420 4752
rect 16212 4700 16264 4752
rect 17040 4743 17092 4752
rect 17040 4709 17049 4743
rect 17049 4709 17083 4743
rect 17083 4709 17092 4743
rect 17040 4700 17092 4709
rect 2780 4632 2832 4684
rect 5540 4632 5592 4684
rect 10600 4632 10652 4684
rect 16948 4632 17000 4684
rect 4620 4564 4672 4616
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 17408 4632 17460 4684
rect 26424 4632 26476 4684
rect 1676 4496 1728 4548
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 11704 4428 11756 4480
rect 13636 4471 13688 4480
rect 13636 4437 13645 4471
rect 13645 4437 13679 4471
rect 13679 4437 13688 4471
rect 13636 4428 13688 4437
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 2780 4088 2832 4140
rect 4988 4088 5040 4140
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 6276 4224 6328 4276
rect 6368 4224 6420 4276
rect 14096 4267 14148 4276
rect 14096 4233 14105 4267
rect 14105 4233 14139 4267
rect 14139 4233 14148 4267
rect 14096 4224 14148 4233
rect 17040 4267 17092 4276
rect 17040 4233 17049 4267
rect 17049 4233 17083 4267
rect 17083 4233 17092 4267
rect 17040 4224 17092 4233
rect 17408 4267 17460 4276
rect 17408 4233 17417 4267
rect 17417 4233 17451 4267
rect 17451 4233 17460 4267
rect 17408 4224 17460 4233
rect 26424 4224 26476 4276
rect 5356 4088 5408 4097
rect 14280 4156 14332 4208
rect 15476 4156 15528 4208
rect 17132 4156 17184 4208
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 5080 4063 5132 4072
rect 4528 4020 4580 4029
rect 2596 3952 2648 4004
rect 4620 3952 4672 4004
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 10232 4020 10284 4072
rect 15292 4020 15344 4072
rect 16304 4020 16356 4072
rect 26424 4063 26476 4072
rect 26424 4029 26433 4063
rect 26433 4029 26467 4063
rect 26467 4029 26476 4063
rect 26424 4020 26476 4029
rect 13728 3952 13780 4004
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 2780 3884 2832 3936
rect 3792 3927 3844 3936
rect 3792 3893 3801 3927
rect 3801 3893 3835 3927
rect 3835 3893 3844 3927
rect 3792 3884 3844 3893
rect 4712 3927 4764 3936
rect 4712 3893 4721 3927
rect 4721 3893 4755 3927
rect 4755 3893 4764 3927
rect 4712 3884 4764 3893
rect 10600 3884 10652 3936
rect 26608 3927 26660 3936
rect 26608 3893 26617 3927
rect 26617 3893 26651 3927
rect 26651 3893 26660 3927
rect 26608 3884 26660 3893
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 4712 3680 4764 3732
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 10600 3723 10652 3732
rect 10600 3689 10609 3723
rect 10609 3689 10643 3723
rect 10643 3689 10652 3723
rect 10600 3680 10652 3689
rect 15292 3680 15344 3732
rect 26700 3723 26752 3732
rect 26700 3689 26709 3723
rect 26709 3689 26743 3723
rect 26743 3689 26752 3723
rect 26700 3680 26752 3689
rect 4896 3612 4948 3664
rect 1768 3544 1820 3596
rect 2964 3544 3016 3596
rect 4068 3544 4120 3596
rect 10232 3544 10284 3596
rect 11612 3544 11664 3596
rect 11796 3587 11848 3596
rect 11796 3553 11830 3587
rect 11830 3553 11848 3587
rect 11796 3544 11848 3553
rect 15200 3544 15252 3596
rect 25320 3587 25372 3596
rect 25320 3553 25329 3587
rect 25329 3553 25363 3587
rect 25363 3553 25372 3587
rect 25320 3544 25372 3553
rect 26792 3544 26844 3596
rect 1492 3476 1544 3528
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 22100 3476 22152 3528
rect 23204 3476 23256 3528
rect 4620 3408 4672 3460
rect 10784 3408 10836 3460
rect 2872 3383 2924 3392
rect 2872 3349 2881 3383
rect 2881 3349 2915 3383
rect 2915 3349 2924 3383
rect 2872 3340 2924 3349
rect 12900 3383 12952 3392
rect 12900 3349 12909 3383
rect 12909 3349 12943 3383
rect 12943 3349 12952 3383
rect 12900 3340 12952 3349
rect 13084 3340 13136 3392
rect 16948 3340 17000 3392
rect 25872 3340 25924 3392
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2688 3136 2740 3188
rect 2964 3136 3016 3188
rect 3884 3136 3936 3188
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 5172 3136 5224 3188
rect 5356 3136 5408 3188
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 8852 3179 8904 3188
rect 8852 3145 8861 3179
rect 8861 3145 8895 3179
rect 8895 3145 8904 3179
rect 8852 3136 8904 3145
rect 25136 3179 25188 3188
rect 25136 3145 25145 3179
rect 25145 3145 25179 3179
rect 25179 3145 25188 3179
rect 25136 3136 25188 3145
rect 25320 3136 25372 3188
rect 26608 3179 26660 3188
rect 26608 3145 26617 3179
rect 26617 3145 26651 3179
rect 26651 3145 26660 3179
rect 26608 3136 26660 3145
rect 26792 3136 26844 3188
rect 4988 3068 5040 3120
rect 11612 3068 11664 3120
rect 6276 3043 6328 3052
rect 6276 3009 6285 3043
rect 6285 3009 6319 3043
rect 6319 3009 6328 3043
rect 6276 3000 6328 3009
rect 8852 2932 8904 2984
rect 10232 2932 10284 2984
rect 13084 2975 13136 2984
rect 13084 2941 13093 2975
rect 13093 2941 13127 2975
rect 13127 2941 13136 2975
rect 15200 2975 15252 2984
rect 13084 2932 13136 2941
rect 15200 2941 15209 2975
rect 15209 2941 15243 2975
rect 15243 2941 15252 2975
rect 15200 2932 15252 2941
rect 15384 2932 15436 2984
rect 17592 2932 17644 2984
rect 25136 2932 25188 2984
rect 26424 2975 26476 2984
rect 26424 2941 26433 2975
rect 26433 2941 26467 2975
rect 26467 2941 26476 2975
rect 26424 2932 26476 2941
rect 27528 2975 27580 2984
rect 27528 2941 27537 2975
rect 27537 2941 27571 2975
rect 27571 2941 27580 2975
rect 27528 2932 27580 2941
rect 480 2864 532 2916
rect 5632 2864 5684 2916
rect 8300 2907 8352 2916
rect 8300 2873 8309 2907
rect 8309 2873 8343 2907
rect 8343 2873 8352 2907
rect 8300 2864 8352 2873
rect 10600 2864 10652 2916
rect 12900 2907 12952 2916
rect 12900 2873 12909 2907
rect 12909 2873 12943 2907
rect 12943 2873 12952 2907
rect 12900 2864 12952 2873
rect 3332 2839 3384 2848
rect 3332 2805 3341 2839
rect 3341 2805 3375 2839
rect 3375 2805 3384 2839
rect 3332 2796 3384 2805
rect 10876 2796 10928 2848
rect 11796 2839 11848 2848
rect 11796 2805 11805 2839
rect 11805 2805 11839 2839
rect 11839 2805 11848 2839
rect 11796 2796 11848 2805
rect 13820 2796 13872 2848
rect 16580 2796 16632 2848
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 18420 2839 18472 2848
rect 18420 2805 18429 2839
rect 18429 2805 18463 2839
rect 18463 2805 18472 2839
rect 18420 2796 18472 2805
rect 25504 2839 25556 2848
rect 25504 2805 25513 2839
rect 25513 2805 25547 2839
rect 25547 2805 25556 2839
rect 25504 2796 25556 2805
rect 27712 2839 27764 2848
rect 27712 2805 27721 2839
rect 27721 2805 27755 2839
rect 27755 2805 27764 2839
rect 27712 2796 27764 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 1768 2592 1820 2644
rect 3516 2592 3568 2644
rect 5816 2592 5868 2644
rect 2504 2388 2556 2440
rect 5448 2524 5500 2576
rect 7748 2567 7800 2576
rect 7748 2533 7757 2567
rect 7757 2533 7791 2567
rect 7791 2533 7800 2567
rect 7748 2524 7800 2533
rect 6644 2456 6696 2508
rect 9588 2592 9640 2644
rect 10232 2635 10284 2644
rect 10232 2601 10241 2635
rect 10241 2601 10275 2635
rect 10275 2601 10284 2635
rect 10232 2592 10284 2601
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 11612 2635 11664 2644
rect 11612 2601 11621 2635
rect 11621 2601 11655 2635
rect 11655 2601 11664 2635
rect 11612 2592 11664 2601
rect 13820 2635 13872 2644
rect 13820 2601 13829 2635
rect 13829 2601 13863 2635
rect 13863 2601 13872 2635
rect 13820 2592 13872 2601
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 17040 2592 17092 2644
rect 19616 2635 19668 2644
rect 19616 2601 19625 2635
rect 19625 2601 19659 2635
rect 19659 2601 19668 2635
rect 19616 2592 19668 2601
rect 23020 2635 23072 2644
rect 23020 2601 23029 2635
rect 23029 2601 23063 2635
rect 23063 2601 23072 2635
rect 23020 2592 23072 2601
rect 12900 2456 12952 2508
rect 16488 2524 16540 2576
rect 15384 2456 15436 2508
rect 18144 2456 18196 2508
rect 19432 2499 19484 2508
rect 19432 2465 19441 2499
rect 19441 2465 19475 2499
rect 19475 2465 19484 2499
rect 19432 2456 19484 2465
rect 22836 2499 22888 2508
rect 22836 2465 22845 2499
rect 22845 2465 22879 2499
rect 22879 2465 22888 2499
rect 22836 2456 22888 2465
rect 24584 2499 24636 2508
rect 24584 2465 24593 2499
rect 24593 2465 24627 2499
rect 24627 2465 24636 2499
rect 24584 2456 24636 2465
rect 25688 2499 25740 2508
rect 25688 2465 25697 2499
rect 25697 2465 25731 2499
rect 25731 2465 25740 2499
rect 25688 2456 25740 2465
rect 26884 2499 26936 2508
rect 26884 2465 26893 2499
rect 26893 2465 26927 2499
rect 26927 2465 26936 2499
rect 26884 2456 26936 2465
rect 12808 2320 12860 2372
rect 18512 2363 18564 2372
rect 14740 2252 14792 2304
rect 18512 2329 18521 2363
rect 18521 2329 18555 2363
rect 18555 2329 18564 2363
rect 18512 2320 18564 2329
rect 15844 2252 15896 2304
rect 24768 2295 24820 2304
rect 24768 2261 24777 2295
rect 24777 2261 24811 2295
rect 24811 2261 24820 2295
rect 24768 2252 24820 2261
rect 25872 2295 25924 2304
rect 25872 2261 25881 2295
rect 25881 2261 25915 2295
rect 25915 2261 25924 2295
rect 25872 2252 25924 2261
rect 27068 2295 27120 2304
rect 27068 2261 27077 2295
rect 27077 2261 27111 2295
rect 27111 2261 27120 2295
rect 27068 2252 27120 2261
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
<< metal2 >>
rect 754 23520 810 24000
rect 2226 23520 2282 24000
rect 3698 23520 3754 24000
rect 4066 23624 4122 23633
rect 4066 23559 4122 23568
rect 768 20369 796 23520
rect 754 20360 810 20369
rect 754 20295 810 20304
rect 2240 19825 2268 23520
rect 3330 23080 3386 23089
rect 3330 23015 3386 23024
rect 3344 22574 3372 23015
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 2870 22400 2926 22409
rect 2870 22335 2926 22344
rect 2226 19816 2282 19825
rect 2226 19751 2282 19760
rect 2686 13832 2742 13841
rect 2686 13767 2742 13776
rect 2700 13394 2728 13767
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 1412 11121 1440 13126
rect 1688 12986 1716 13330
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 2608 12782 2636 13262
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2686 12744 2742 12753
rect 2136 12708 2188 12714
rect 2686 12679 2688 12688
rect 2136 12650 2188 12656
rect 2740 12679 2742 12688
rect 2688 12650 2740 12656
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1582 11656 1638 11665
rect 1582 11591 1638 11600
rect 1398 11112 1454 11121
rect 1398 11047 1454 11056
rect 1596 10810 1624 11591
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1964 11393 1992 11494
rect 1950 11384 2006 11393
rect 1950 11319 2006 11328
rect 2056 11268 2084 11834
rect 1964 11240 2084 11268
rect 1766 11112 1822 11121
rect 1766 11047 1822 11056
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1582 10432 1638 10441
rect 1582 10367 1638 10376
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 1412 9178 1440 9823
rect 1596 9654 1624 10367
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1490 9344 1546 9353
rect 1490 9279 1546 9288
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1504 8634 1532 9279
rect 1582 8664 1638 8673
rect 1492 8628 1544 8634
rect 1582 8599 1638 8608
rect 1492 8570 1544 8576
rect 1596 8090 1624 8599
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1584 7472 1636 7478
rect 1582 7440 1584 7449
rect 1636 7440 1638 7449
rect 1582 7375 1638 7384
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1596 6730 1624 6831
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5681 1624 6054
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1596 5137 1624 5510
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 480 2916 532 2922
rect 480 2858 532 2864
rect 492 480 520 2858
rect 1412 1465 1440 4966
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1584 4480 1636 4486
rect 1582 4448 1584 4457
rect 1636 4448 1638 4457
rect 1582 4383 1638 4392
rect 1584 3936 1636 3942
rect 1582 3904 1584 3913
rect 1636 3904 1638 3913
rect 1582 3839 1638 3848
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1398 1456 1454 1465
rect 1398 1391 1454 1400
rect 1504 480 1532 3470
rect 1688 921 1716 4490
rect 1780 3602 1808 11047
rect 1964 6866 1992 11240
rect 2042 10704 2098 10713
rect 2042 10639 2044 10648
rect 2096 10639 2098 10648
rect 2044 10610 2096 10616
rect 2148 9654 2176 12650
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2240 11694 2268 12582
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2424 11762 2452 12038
rect 2792 11898 2820 12378
rect 2884 12306 2912 22335
rect 3330 21856 3386 21865
rect 3330 21791 3386 21800
rect 3344 20806 3372 21791
rect 3712 21146 3740 23520
rect 4080 22166 4108 23559
rect 5170 23520 5226 24000
rect 6734 23520 6790 24000
rect 8206 23520 8262 24000
rect 9678 23520 9734 24000
rect 11242 23520 11298 24000
rect 12714 23520 12770 24000
rect 14186 23520 14242 24000
rect 15750 23520 15806 24000
rect 17222 23520 17278 24000
rect 18694 23520 18750 24000
rect 20166 23520 20222 24000
rect 21730 23520 21786 24000
rect 23202 23520 23258 24000
rect 24674 23520 24730 24000
rect 25686 23624 25742 23633
rect 25686 23559 25742 23568
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 3882 21312 3938 21321
rect 3882 21247 3938 21256
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3896 21010 3924 21247
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 5184 20874 5212 23520
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 6368 21072 6420 21078
rect 6368 21014 6420 21020
rect 5172 20868 5224 20874
rect 5172 20810 5224 20816
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 4066 20088 4122 20097
rect 4066 20023 4122 20032
rect 2962 18864 3018 18873
rect 2962 18799 3018 18808
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2594 11792 2650 11801
rect 2412 11756 2464 11762
rect 2594 11727 2596 11736
rect 2412 11698 2464 11704
rect 2648 11727 2650 11736
rect 2596 11698 2648 11704
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2608 11286 2636 11698
rect 2596 11280 2648 11286
rect 2596 11222 2648 11228
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2332 10266 2360 11154
rect 2608 10810 2636 11222
rect 2686 11112 2742 11121
rect 2742 11082 2820 11098
rect 2742 11076 2832 11082
rect 2742 11070 2780 11076
rect 2686 11047 2742 11056
rect 2780 11018 2832 11024
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2884 10810 2912 10950
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2884 10198 2912 10746
rect 2976 10198 3004 18799
rect 3422 16416 3478 16425
rect 3422 16351 3478 16360
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3068 11558 3096 12242
rect 3146 12200 3202 12209
rect 3146 12135 3202 12144
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3068 10441 3096 11494
rect 3054 10432 3110 10441
rect 3054 10367 3110 10376
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2424 9178 2452 9930
rect 2516 9382 2544 10066
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2792 9654 2820 9998
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2332 8634 2360 8978
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2332 8401 2360 8570
rect 2318 8392 2374 8401
rect 2318 8327 2374 8336
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2424 7857 2452 7890
rect 2410 7848 2466 7857
rect 2410 7783 2466 7792
rect 2424 7546 2452 7783
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2516 7449 2544 9318
rect 3068 8838 3096 9318
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2700 8129 2728 8502
rect 2686 8120 2742 8129
rect 2686 8055 2742 8064
rect 2686 7984 2742 7993
rect 2686 7919 2742 7928
rect 2502 7440 2558 7449
rect 2502 7375 2558 7384
rect 2134 7304 2190 7313
rect 2134 7239 2190 7248
rect 2044 7200 2096 7206
rect 2042 7168 2044 7177
rect 2096 7168 2098 7177
rect 2042 7103 2098 7112
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1964 6458 1992 6802
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 2148 6254 2176 7239
rect 2700 7018 2728 7919
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2976 7410 3004 7686
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2332 6990 2728 7018
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2148 5914 2176 6190
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2044 5024 2096 5030
rect 2042 4992 2044 5001
rect 2096 4992 2098 5001
rect 2042 4927 2098 4936
rect 2332 4826 2360 6990
rect 2596 6928 2648 6934
rect 2502 6896 2558 6905
rect 2596 6870 2648 6876
rect 2502 6831 2504 6840
rect 2556 6831 2558 6840
rect 2504 6802 2556 6808
rect 2410 6760 2466 6769
rect 2410 6695 2466 6704
rect 2424 5778 2452 6695
rect 2516 6458 2544 6802
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2424 5370 2452 5714
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2410 4720 2466 4729
rect 2410 4655 2466 4664
rect 2424 4146 2452 4655
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2608 4010 2636 6870
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6361 2728 6598
rect 2686 6352 2742 6361
rect 2686 6287 2742 6296
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2596 4004 2648 4010
rect 2596 3946 2648 3952
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 2650 1808 3538
rect 2700 3194 2728 6054
rect 3068 5760 3096 8774
rect 3160 8634 3188 12135
rect 3238 11520 3294 11529
rect 3238 11455 3294 11464
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3160 8430 3188 8570
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3252 6934 3280 11455
rect 3436 11257 3464 16351
rect 3698 15328 3754 15337
rect 3698 15263 3754 15272
rect 3606 14648 3662 14657
rect 3606 14583 3662 14592
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3528 12238 3556 12786
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3528 11558 3556 12174
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3422 11248 3478 11257
rect 3422 11183 3478 11192
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3344 10470 3372 10950
rect 3528 10674 3556 11494
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3528 10577 3556 10610
rect 3514 10568 3570 10577
rect 3424 10532 3476 10538
rect 3514 10503 3570 10512
rect 3424 10474 3476 10480
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 9178 3372 10406
rect 3436 9926 3464 10474
rect 3528 10062 3556 10503
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3436 9722 3464 9862
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3436 7041 3464 9318
rect 3422 7032 3478 7041
rect 3422 6967 3478 6976
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6254 3464 6802
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3528 5914 3556 6054
rect 3620 5953 3648 14583
rect 3712 9450 3740 15263
rect 4080 15065 4108 20023
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 4066 14104 4122 14113
rect 4066 14039 4122 14048
rect 3974 13424 4030 13433
rect 3974 13359 4030 13368
rect 3882 12880 3938 12889
rect 3882 12815 3938 12824
rect 3896 11937 3924 12815
rect 3882 11928 3938 11937
rect 3882 11863 3938 11872
rect 3988 10305 4016 13359
rect 3974 10296 4030 10305
rect 3974 10231 4030 10240
rect 4080 10248 4108 14039
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4172 12238 4200 12718
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4526 11928 4582 11937
rect 4724 11898 4752 12174
rect 4526 11863 4582 11872
rect 4712 11892 4764 11898
rect 4342 11384 4398 11393
rect 4342 11319 4398 11328
rect 4436 11348 4488 11354
rect 4356 11218 4384 11319
rect 4436 11290 4488 11296
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4356 10674 4384 11154
rect 4448 10742 4476 11290
rect 4436 10736 4488 10742
rect 4436 10678 4488 10684
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4080 10220 4200 10248
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3804 9110 3832 9522
rect 4172 9518 4200 10220
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4540 9178 4568 11863
rect 4712 11834 4764 11840
rect 4908 11830 4936 12310
rect 4896 11824 4948 11830
rect 4894 11792 4896 11801
rect 4948 11792 4950 11801
rect 4894 11727 4950 11736
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4632 11150 4660 11562
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4632 10810 4660 11086
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4618 10296 4674 10305
rect 4618 10231 4674 10240
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3804 8634 3832 9046
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 4448 8362 4476 8978
rect 4540 8634 4568 9114
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3988 7002 4016 7822
rect 4172 7206 4200 7890
rect 4160 7200 4212 7206
rect 4080 7160 4160 7188
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 4080 6322 4108 7160
rect 4160 7142 4212 7148
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3606 5944 3662 5953
rect 3516 5908 3568 5914
rect 3606 5879 3662 5888
rect 3516 5850 3568 5856
rect 2976 5732 3096 5760
rect 4344 5772 4396 5778
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 2792 4690 2820 5199
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2792 4146 2820 4626
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 2516 480 2544 2382
rect 2792 2145 2820 3878
rect 2976 3602 3004 5732
rect 4344 5714 4396 5720
rect 3882 5672 3938 5681
rect 3882 5607 3938 5616
rect 4068 5636 4120 5642
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2872 3392 2924 3398
rect 2870 3360 2872 3369
rect 2924 3360 2926 3369
rect 2870 3295 2926 3304
rect 2976 3194 3004 3538
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 3606 2952 3662 2961
rect 3606 2887 3662 2896
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 3344 2689 3372 2790
rect 3330 2680 3386 2689
rect 3330 2615 3386 2624
rect 3514 2680 3570 2689
rect 3514 2615 3516 2624
rect 3568 2615 3570 2624
rect 3516 2586 3568 2592
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 3620 1714 3648 2887
rect 3528 1686 3648 1714
rect 3528 480 3556 1686
rect 478 0 534 480
rect 1490 0 1546 480
rect 2502 0 2558 480
rect 3514 0 3570 480
rect 3804 377 3832 3878
rect 3896 3194 3924 5607
rect 4068 5578 4120 5584
rect 4080 5370 4108 5578
rect 4356 5370 4384 5714
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4448 5273 4476 8298
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4434 5264 4490 5273
rect 4434 5199 4490 5208
rect 4540 4826 4568 5646
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4632 4706 4660 10231
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4986 10024 5042 10033
rect 4724 9722 4752 9998
rect 4986 9959 5042 9968
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4908 9364 4936 9862
rect 5000 9518 5028 9959
rect 5092 9625 5120 20742
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5814 20632 5870 20641
rect 5956 20624 6252 20644
rect 5814 20567 5870 20576
rect 5354 18320 5410 18329
rect 5354 18255 5410 18264
rect 5630 18320 5686 18329
rect 5630 18255 5686 18264
rect 5078 9616 5134 9625
rect 5078 9551 5134 9560
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4988 9376 5040 9382
rect 4908 9336 4988 9364
rect 4988 9318 5040 9324
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8362 4936 8774
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4724 5710 4752 7346
rect 4908 6905 4936 8298
rect 4894 6896 4950 6905
rect 4894 6831 4950 6840
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4816 5234 4844 5510
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4712 5160 4764 5166
rect 4710 5128 4712 5137
rect 4764 5128 4766 5137
rect 4710 5063 4766 5072
rect 4540 4678 4660 4706
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4540 4078 4568 4678
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4632 4010 4660 4558
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4066 3904 4122 3913
rect 4066 3839 4122 3848
rect 4080 3602 4108 3839
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4632 3466 4660 3946
rect 4724 3942 4752 4694
rect 4908 4622 4936 5170
rect 5000 4729 5028 9318
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5184 7188 5212 8230
rect 5264 7200 5316 7206
rect 5184 7160 5264 7188
rect 5092 6934 5120 7142
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 5184 6866 5212 7160
rect 5264 7142 5316 7148
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5368 5137 5396 18255
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12374 5580 12582
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5460 9586 5488 10066
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5460 9382 5488 9522
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 8974 5488 9318
rect 5644 9058 5672 18255
rect 5828 10169 5856 20567
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 6274 18728 6330 18737
rect 6274 18663 6330 18672
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 6288 12442 6316 18663
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 6288 11626 6316 12038
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 6090 10568 6146 10577
rect 6090 10503 6146 10512
rect 6104 10266 6132 10503
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 5814 10160 5870 10169
rect 5814 10095 5870 10104
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 5722 9616 5778 9625
rect 5722 9551 5778 9560
rect 5552 9030 5672 9058
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5460 8090 5488 8910
rect 5552 8838 5580 9030
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5644 8090 5672 8910
rect 5736 8430 5764 9551
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 5724 8424 5776 8430
rect 6380 8401 6408 21014
rect 6748 20505 6776 23520
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 6734 20496 6790 20505
rect 6734 20431 6790 20440
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7116 12442 7144 12786
rect 7392 12782 7420 13466
rect 7668 13394 7696 22510
rect 8220 20942 8248 23520
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 9588 20596 9640 20602
rect 9692 20584 9720 23520
rect 11256 21434 11284 23520
rect 11256 21406 11376 21434
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 11348 20602 11376 21406
rect 12728 20602 12756 23520
rect 14200 23474 14228 23520
rect 13832 23446 14228 23474
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 9640 20556 9720 20584
rect 11336 20596 11388 20602
rect 9588 20538 9640 20544
rect 11336 20538 11388 20544
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12728 20398 12756 20538
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 8758 14512 8814 14521
rect 8024 14476 8076 14482
rect 8758 14447 8814 14456
rect 8024 14418 8076 14424
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 13530 7788 14214
rect 7840 13864 7892 13870
rect 7838 13832 7840 13841
rect 7892 13832 7894 13841
rect 7838 13767 7894 13776
rect 7944 13530 7972 14282
rect 8036 14074 8064 14418
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8220 14074 8248 14350
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8220 13530 8248 14010
rect 8482 13968 8538 13977
rect 8300 13932 8352 13938
rect 8482 13903 8538 13912
rect 8300 13874 8352 13880
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 7562 13152 7618 13161
rect 7562 13087 7618 13096
rect 7576 12850 7604 13087
rect 8128 12986 8156 13330
rect 8312 13258 8340 13874
rect 8496 13870 8524 13903
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8772 13530 8800 14447
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6840 11354 6868 11698
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6840 9722 6868 10202
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6734 9480 6790 9489
rect 6734 9415 6790 9424
rect 5724 8366 5776 8372
rect 6366 8392 6422 8401
rect 6366 8327 6422 8336
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 6380 8022 6408 8327
rect 6368 8016 6420 8022
rect 6368 7958 6420 7964
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5644 7002 5672 7278
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5828 6934 5856 7346
rect 6288 7342 6316 7686
rect 6380 7546 6408 7958
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 6472 6866 6500 7142
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 6288 6458 6316 6802
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6380 6390 6408 6734
rect 6368 6384 6420 6390
rect 6090 6352 6146 6361
rect 6368 6326 6420 6332
rect 6090 6287 6146 6296
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 5302 5580 6054
rect 6104 5953 6132 6287
rect 5722 5944 5778 5953
rect 5722 5879 5778 5888
rect 6090 5944 6146 5953
rect 6090 5879 6092 5888
rect 5736 5370 5764 5879
rect 6144 5879 6146 5888
rect 6092 5850 6144 5856
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 6012 5681 6040 5782
rect 6276 5704 6328 5710
rect 5998 5672 6054 5681
rect 6276 5646 6328 5652
rect 5998 5607 6054 5616
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 6288 5370 6316 5646
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5354 5128 5410 5137
rect 5354 5063 5410 5072
rect 5078 4992 5134 5001
rect 5078 4927 5134 4936
rect 4986 4720 5042 4729
rect 4986 4655 5042 4664
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4724 3738 4752 3878
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4908 3670 4936 4558
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5000 3754 5028 4082
rect 5092 4078 5120 4927
rect 6288 4758 6316 5306
rect 6380 4758 6408 6326
rect 6472 6118 6500 6802
rect 6550 6488 6606 6497
rect 6550 6423 6606 6432
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6564 5846 6592 6423
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6564 5302 6592 5782
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 6748 5001 6776 9415
rect 6932 9382 6960 10066
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 8566 6960 9318
rect 6920 8560 6972 8566
rect 6840 8520 6920 8548
rect 6840 6458 6868 8520
rect 6920 8502 6972 8508
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 7886 6960 8230
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6932 7206 6960 7822
rect 7024 7546 7052 8026
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6734 4992 6790 5001
rect 6734 4927 6790 4936
rect 6840 4808 6868 6054
rect 6920 4820 6972 4826
rect 6840 4780 6920 4808
rect 6920 4762 6972 4768
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6368 4752 6420 4758
rect 6368 4694 6420 4700
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5078 3768 5134 3777
rect 5000 3726 5078 3754
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4526 2816 4582 2825
rect 4526 2751 4582 2760
rect 4540 480 4568 2751
rect 4816 2553 4844 3130
rect 5000 3126 5028 3726
rect 5078 3703 5080 3712
rect 5132 3703 5134 3712
rect 5080 3674 5132 3680
rect 5368 3534 5396 4082
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5184 3194 5212 3470
rect 5368 3194 5396 3470
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5552 2802 5580 4626
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 6288 4282 6316 4694
rect 6380 4282 6408 4694
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5460 2774 5580 2802
rect 5460 2582 5488 2774
rect 5448 2576 5500 2582
rect 4802 2544 4858 2553
rect 5448 2518 5500 2524
rect 4802 2479 4858 2488
rect 5644 480 5672 2858
rect 5828 2650 5856 3130
rect 6274 3088 6330 3097
rect 6274 3023 6276 3032
rect 6328 3023 6330 3032
rect 6276 2994 6328 3000
rect 7208 2689 7236 12582
rect 8312 12442 8340 13194
rect 8588 12782 8616 13398
rect 8772 12986 8800 13466
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8588 12442 8616 12718
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 11218 7512 11494
rect 8312 11354 8340 12378
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7392 10742 7420 11154
rect 7484 10810 7512 11154
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7392 10266 7420 10678
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7484 8634 7512 9046
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7668 8090 7696 8366
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7852 7886 7880 10202
rect 8390 10160 8446 10169
rect 8390 10095 8446 10104
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 9586 8340 9862
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8401 8064 8774
rect 8128 8634 8156 8910
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8206 8528 8262 8537
rect 8206 8463 8208 8472
rect 8260 8463 8262 8472
rect 8208 8434 8260 8440
rect 8022 8392 8078 8401
rect 8022 8327 8078 8336
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7562 7712 7618 7721
rect 7562 7647 7618 7656
rect 7576 7313 7604 7647
rect 7852 7546 7880 7822
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7562 7304 7618 7313
rect 7562 7239 7618 7248
rect 8312 6769 8340 9522
rect 8404 9450 8432 10095
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8496 9178 8524 9318
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8496 8634 8524 9114
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8588 7546 8616 8910
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8298 6760 8354 6769
rect 8298 6695 8354 6704
rect 8588 6458 8616 7482
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8298 2952 8354 2961
rect 7668 2910 7880 2938
rect 7194 2680 7250 2689
rect 5816 2644 5868 2650
rect 7194 2615 7250 2624
rect 5816 2586 5868 2592
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 6656 480 6684 2450
rect 7668 480 7696 2910
rect 7746 2816 7802 2825
rect 7852 2802 7880 2910
rect 8298 2887 8300 2896
rect 8352 2887 8354 2896
rect 8300 2858 8352 2864
rect 7930 2816 7986 2825
rect 7852 2774 7930 2802
rect 7746 2751 7802 2760
rect 7930 2751 7986 2760
rect 7760 2582 7788 2751
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 8680 480 8708 8298
rect 8772 8072 8800 12922
rect 9140 12714 9168 13126
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 9048 12170 9076 12582
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9128 11552 9180 11558
rect 9126 11520 9128 11529
rect 9180 11520 9182 11529
rect 9126 11455 9182 11464
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8956 10810 8984 10950
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 10305 9168 10406
rect 9126 10296 9182 10305
rect 9126 10231 9182 10240
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8956 8129 8984 9318
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9232 8922 9260 20198
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 9954 19952 10010 19961
rect 9954 19887 10010 19896
rect 9310 17096 9366 17105
rect 9310 17031 9366 17040
rect 9324 9926 9352 17031
rect 9678 15872 9734 15881
rect 9678 15807 9734 15816
rect 9494 13424 9550 13433
rect 9494 13359 9496 13368
rect 9548 13359 9550 13368
rect 9496 13330 9548 13336
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9048 8498 9076 8910
rect 9232 8894 9352 8922
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8942 8120 8998 8129
rect 8772 8044 8892 8072
rect 8942 8055 8998 8064
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8772 7478 8800 7890
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8772 7342 8800 7414
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8864 7177 8892 8044
rect 9048 7857 9076 8434
rect 9232 8362 9260 8774
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9034 7848 9090 7857
rect 9034 7783 9090 7792
rect 9128 7336 9180 7342
rect 9126 7304 9128 7313
rect 9180 7304 9182 7313
rect 9036 7268 9088 7274
rect 9126 7239 9182 7248
rect 9036 7210 9088 7216
rect 8944 7200 8996 7206
rect 8850 7168 8906 7177
rect 8944 7142 8996 7148
rect 8850 7103 8906 7112
rect 8956 6934 8984 7142
rect 9048 7002 9076 7210
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 9140 6866 9168 7239
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8956 5914 8984 6190
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9324 4049 9352 8894
rect 9310 4040 9366 4049
rect 9310 3975 9366 3984
rect 9416 3777 9444 10950
rect 9600 10248 9628 12650
rect 9692 11626 9720 15807
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9692 11150 9720 11181
rect 9680 11144 9732 11150
rect 9678 11112 9680 11121
rect 9732 11112 9734 11121
rect 9678 11047 9734 11056
rect 9692 10810 9720 11047
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9784 10266 9812 11494
rect 9968 11370 9996 19887
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 10598 16688 10654 16697
rect 10598 16623 10654 16632
rect 10230 16008 10286 16017
rect 10230 15943 10286 15952
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10152 12850 10180 13330
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 9876 11342 9996 11370
rect 10060 11354 10088 12242
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10152 11898 10180 12174
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10048 11348 10100 11354
rect 9680 10260 9732 10266
rect 9600 10220 9680 10248
rect 9680 10202 9732 10208
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9876 10130 9904 11342
rect 10048 11290 10100 11296
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9770 10024 9826 10033
rect 9770 9959 9826 9968
rect 9784 7993 9812 9959
rect 9876 9382 9904 10066
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9770 7984 9826 7993
rect 9770 7919 9826 7928
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7410 9536 7686
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9402 3768 9458 3777
rect 9402 3703 9458 3712
rect 8850 3224 8906 3233
rect 8850 3159 8852 3168
rect 8904 3159 8906 3168
rect 8852 3130 8904 3136
rect 8864 2990 8892 3130
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 9588 2644 9640 2650
rect 9692 2632 9720 6598
rect 9876 6225 9904 9318
rect 9968 8974 9996 11222
rect 10060 10810 10088 11290
rect 10152 11082 10180 11834
rect 10244 11694 10272 15943
rect 10506 14920 10562 14929
rect 10506 14855 10562 14864
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10336 12306 10364 12650
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10336 11914 10364 12242
rect 10336 11886 10456 11914
rect 10428 11830 10456 11886
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10244 11121 10272 11494
rect 10336 11150 10364 11698
rect 10324 11144 10376 11150
rect 10230 11112 10286 11121
rect 10140 11076 10192 11082
rect 10324 11086 10376 11092
rect 10230 11047 10286 11056
rect 10140 11018 10192 11024
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10336 10674 10364 11086
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10428 10554 10456 11766
rect 10520 11286 10548 14855
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10336 10526 10456 10554
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10152 9489 10180 10406
rect 10336 10062 10364 10526
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 9654 10364 9998
rect 10428 9722 10456 10202
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10324 9512 10376 9518
rect 10138 9480 10194 9489
rect 10324 9454 10376 9460
rect 10138 9415 10194 9424
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 10060 8090 10088 8978
rect 10152 8945 10180 9415
rect 10336 8974 10364 9454
rect 10324 8968 10376 8974
rect 10138 8936 10194 8945
rect 10324 8910 10376 8916
rect 10138 8871 10194 8880
rect 10138 8256 10194 8265
rect 10138 8191 10194 8200
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10152 7002 10180 8191
rect 10336 7818 10364 8910
rect 10520 7857 10548 11018
rect 10506 7848 10562 7857
rect 10324 7812 10376 7818
rect 10506 7783 10562 7792
rect 10324 7754 10376 7760
rect 10612 7585 10640 16623
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10690 12880 10746 12889
rect 10690 12815 10746 12824
rect 10704 10713 10732 12815
rect 11072 12714 11100 13330
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10888 12442 10916 12582
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 11348 12442 11376 13398
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12176 13190 12204 13330
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12164 13184 12216 13190
rect 12162 13152 12164 13161
rect 12216 13152 12218 13161
rect 12162 13087 12218 13096
rect 12176 12986 12204 13087
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11348 12102 11376 12378
rect 12912 12102 12940 13262
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 10782 11656 10838 11665
rect 10782 11591 10838 11600
rect 10796 11354 10824 11591
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 11520 11076 11572 11082
rect 11520 11018 11572 11024
rect 10690 10704 10746 10713
rect 10690 10639 10746 10648
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 11348 8634 11376 10542
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10598 7576 10654 7585
rect 10598 7511 10654 7520
rect 10612 7342 10640 7511
rect 10704 7410 10732 7686
rect 10888 7410 10916 7754
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 11348 7342 11376 8230
rect 11532 8090 11560 11018
rect 12912 10130 12940 12038
rect 13096 11778 13124 20198
rect 13464 12374 13492 22102
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13452 12368 13504 12374
rect 13450 12336 13452 12345
rect 13504 12336 13506 12345
rect 13450 12271 13506 12280
rect 13176 12232 13228 12238
rect 13174 12200 13176 12209
rect 13228 12200 13230 12209
rect 13174 12135 13230 12144
rect 13188 11898 13216 12135
rect 13464 11898 13492 12271
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 11898 13584 12038
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13096 11750 13584 11778
rect 12990 11520 13046 11529
rect 12990 11455 13046 11464
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12912 9586 12940 10066
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11624 8498 11652 8978
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11624 8294 11652 8434
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11520 8084 11572 8090
rect 11440 8044 11520 8072
rect 11440 7546 11468 8044
rect 11520 8026 11572 8032
rect 11624 7886 11652 8230
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 10140 6996 10192 7002
rect 10192 6956 10272 6984
rect 10140 6938 10192 6944
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10152 6390 10180 6734
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10244 6322 10272 6956
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 6458 10364 6734
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 9862 6216 9918 6225
rect 9862 6151 9918 6160
rect 10336 5914 10364 6394
rect 11348 6361 11376 7142
rect 11440 6497 11468 7482
rect 11532 7206 11560 7822
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11624 7002 11652 7822
rect 11808 7546 11836 9454
rect 12084 9382 12112 9522
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 9110 12112 9318
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 12084 8090 12112 9046
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12254 8664 12310 8673
rect 12254 8599 12310 8608
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11426 6488 11482 6497
rect 11426 6423 11482 6432
rect 11334 6352 11390 6361
rect 11334 6287 11390 6296
rect 11808 6254 11836 7482
rect 12268 7478 12296 8599
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11900 7002 11928 7278
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10336 5370 10364 5850
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10428 5370 10456 5714
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10428 4826 10456 5306
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10244 4078 10272 4762
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10232 4072 10284 4078
rect 9770 4040 9826 4049
rect 10232 4014 10284 4020
rect 9770 3975 9826 3984
rect 9640 2604 9720 2632
rect 9588 2586 9640 2592
rect 9784 480 9812 3975
rect 10244 3602 10272 4014
rect 10612 3942 10640 4626
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3738 10640 3878
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10244 2990 10272 3538
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10244 2650 10272 2926
rect 10612 2922 10640 3674
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10796 480 10824 3402
rect 11624 3126 11652 3538
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 11610 2816 11666 2825
rect 10888 2650 10916 2790
rect 10956 2748 11252 2768
rect 11610 2751 11666 2760
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 11624 2650 11652 2751
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11716 2258 11744 4422
rect 12360 3641 12388 8298
rect 12728 8090 12756 8774
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12728 7410 12756 7686
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12820 7342 12848 8230
rect 13004 8090 13032 11455
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13096 10470 13124 11086
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13096 10130 13124 10406
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13096 9722 13124 10066
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13082 8936 13138 8945
rect 13082 8871 13084 8880
rect 13136 8871 13138 8880
rect 13084 8842 13136 8848
rect 13096 8430 13124 8842
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13004 7970 13032 8026
rect 12912 7942 13032 7970
rect 13084 7948 13136 7954
rect 12808 7336 12860 7342
rect 12438 7304 12494 7313
rect 12808 7278 12860 7284
rect 12438 7239 12494 7248
rect 12452 7206 12480 7239
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12912 7002 12940 7942
rect 13084 7890 13136 7896
rect 13096 7857 13124 7890
rect 13082 7848 13138 7857
rect 12992 7812 13044 7818
rect 13082 7783 13138 7792
rect 12992 7754 13044 7760
rect 13004 7410 13032 7754
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5778 12480 6054
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12544 5681 12572 5782
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12530 5672 12586 5681
rect 12530 5607 12586 5616
rect 12544 5574 12572 5607
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12544 5370 12572 5510
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 13096 5030 13124 5714
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 12346 3632 12402 3641
rect 11796 3596 11848 3602
rect 12346 3567 12402 3576
rect 11796 3538 11848 3544
rect 11808 2854 11836 3538
rect 13096 3398 13124 4966
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 12912 2922 12940 3334
rect 13096 2990 13124 3334
rect 13188 3233 13216 10406
rect 13464 9722 13492 10474
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13464 9178 13492 9522
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13358 8528 13414 8537
rect 13358 8463 13360 8472
rect 13412 8463 13414 8472
rect 13360 8434 13412 8440
rect 13372 7886 13400 8434
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13372 7002 13400 7822
rect 13464 7206 13492 7890
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13464 6474 13492 7142
rect 13372 6446 13492 6474
rect 13174 3224 13230 3233
rect 13174 3159 13230 3168
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 12912 2514 12940 2858
rect 13372 2553 13400 6446
rect 13556 3233 13584 11750
rect 13648 11354 13676 12582
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13740 11218 13768 12038
rect 13832 11234 13860 23446
rect 15764 19378 15792 23520
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15658 17232 15714 17241
rect 15658 17167 15714 17176
rect 15474 15056 15530 15065
rect 15474 14991 15530 15000
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15120 12986 15148 13126
rect 15108 12980 15160 12986
rect 15160 12940 15240 12968
rect 15108 12922 15160 12928
rect 14094 12880 14150 12889
rect 14094 12815 14096 12824
rect 14148 12815 14150 12824
rect 14464 12844 14516 12850
rect 14096 12786 14148 12792
rect 14464 12786 14516 12792
rect 14476 12238 14504 12786
rect 15212 12782 15240 12940
rect 15304 12850 15332 13126
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15212 12442 15240 12582
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 14096 12232 14148 12238
rect 14094 12200 14096 12209
rect 14464 12232 14516 12238
rect 14148 12200 14150 12209
rect 14464 12174 14516 12180
rect 14094 12135 14150 12144
rect 14476 11626 14504 12174
rect 15304 11898 15332 12786
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 13728 11212 13780 11218
rect 13832 11206 14044 11234
rect 14476 11218 14504 11562
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 13728 11154 13780 11160
rect 13634 11112 13690 11121
rect 13740 11098 13768 11154
rect 13740 11070 13860 11098
rect 13634 11047 13690 11056
rect 13648 7857 13676 11047
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13740 10470 13768 10950
rect 13832 10810 13860 11070
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10266 13768 10406
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13634 7848 13690 7857
rect 13634 7783 13690 7792
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13648 6322 13676 6598
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13648 5574 13676 6258
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13924 5914 13952 6122
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 5166 13676 5510
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13542 3224 13598 3233
rect 13542 3159 13598 3168
rect 13648 3097 13676 4422
rect 13740 4010 13768 4762
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13634 3088 13690 3097
rect 13634 3023 13690 3032
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13910 2816 13966 2825
rect 13832 2650 13860 2790
rect 13910 2751 13966 2760
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13358 2544 13414 2553
rect 12900 2508 12952 2514
rect 13358 2479 13414 2488
rect 12900 2450 12952 2456
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 11716 2230 11836 2258
rect 11808 480 11836 2230
rect 12820 480 12848 2314
rect 13372 1873 13400 2479
rect 13358 1864 13414 1873
rect 13358 1799 13414 1808
rect 13924 480 13952 2751
rect 14016 2009 14044 11206
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 15120 11150 15148 11494
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15120 10826 15148 11086
rect 15120 10810 15240 10826
rect 15120 10804 15252 10810
rect 15120 10798 15200 10804
rect 15200 10746 15252 10752
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14384 10266 14412 10610
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14384 9722 14412 10202
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14384 9450 14412 9658
rect 14372 9444 14424 9450
rect 14372 9386 14424 9392
rect 15304 7970 15332 11494
rect 15488 11286 15516 14991
rect 15672 11558 15700 17167
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15856 11370 15884 20946
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 16486 20360 16542 20369
rect 16486 20295 16542 20304
rect 16500 20262 16528 20295
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 17236 19378 17264 23520
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 18234 20360 18290 20369
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 17328 19446 17356 19858
rect 17498 19816 17554 19825
rect 17498 19751 17500 19760
rect 17552 19751 17554 19760
rect 17500 19722 17552 19728
rect 17316 19440 17368 19446
rect 17316 19382 17368 19388
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 16396 12776 16448 12782
rect 16396 12718 16448 12724
rect 16408 12442 16436 12718
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 15580 11342 15884 11370
rect 16304 11348 16356 11354
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15580 11098 15608 11342
rect 16304 11290 16356 11296
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15396 11070 15608 11098
rect 15396 8090 15424 11070
rect 15672 10606 15700 11222
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15764 10606 15792 10950
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15580 8537 15608 9318
rect 15566 8528 15622 8537
rect 15672 8514 15700 10542
rect 15764 10266 15792 10542
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15856 10198 15884 11086
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 16316 10198 16344 11290
rect 16408 10606 16436 11494
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 15844 10192 15896 10198
rect 15750 10160 15806 10169
rect 15844 10134 15896 10140
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 15750 10095 15806 10104
rect 15764 9761 15792 10095
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15750 9752 15806 9761
rect 15956 9744 16252 9764
rect 15750 9687 15806 9696
rect 16394 9072 16450 9081
rect 16394 9007 16450 9016
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 15750 8528 15806 8537
rect 15672 8486 15750 8514
rect 15566 8463 15622 8472
rect 15750 8463 15806 8472
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15304 7942 15424 7970
rect 15106 7712 15162 7721
rect 15106 7647 15162 7656
rect 15120 7546 15148 7647
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14292 4622 14320 4966
rect 15212 4842 15240 6598
rect 15396 5778 15424 7942
rect 15580 7478 15608 8026
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15658 7576 15714 7585
rect 15658 7511 15714 7520
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 15672 6905 15700 7511
rect 15764 6934 15792 7686
rect 15856 7546 15884 7822
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15856 7313 15884 7482
rect 16316 7342 16344 8230
rect 16408 8090 16436 9007
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16500 7562 16528 19314
rect 16578 14240 16634 14249
rect 16578 14175 16634 14184
rect 16592 11082 16620 14175
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16684 11898 16712 12582
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16684 11150 16712 11834
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16578 10160 16634 10169
rect 16578 10095 16634 10104
rect 16408 7534 16528 7562
rect 16304 7336 16356 7342
rect 15842 7304 15898 7313
rect 16304 7278 16356 7284
rect 15842 7239 15898 7248
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15948 7002 15976 7142
rect 16316 7002 16344 7278
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 15752 6928 15804 6934
rect 15658 6896 15714 6905
rect 15752 6870 15804 6876
rect 15658 6831 15714 6840
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15488 6458 15516 6734
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15120 4826 15240 4842
rect 15108 4820 15240 4826
rect 15160 4814 15240 4820
rect 15108 4762 15160 4768
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14108 4282 14136 4558
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14292 4214 14320 4558
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 15304 4078 15332 5510
rect 15396 5030 15424 5714
rect 15488 5166 15516 6394
rect 15764 5914 15792 6870
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16040 6118 16068 6258
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 16040 5846 16068 6054
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 16210 5672 16266 5681
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15396 4185 15424 4966
rect 15488 4214 15516 5102
rect 15764 4826 15792 5646
rect 15856 5370 15884 5646
rect 16210 5607 16212 5616
rect 16264 5607 16266 5616
rect 16212 5578 16264 5584
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 16224 4758 16252 5102
rect 16212 4752 16264 4758
rect 16210 4720 16212 4729
rect 16264 4720 16266 4729
rect 16210 4655 16266 4664
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 15476 4208 15528 4214
rect 15382 4176 15438 4185
rect 15476 4150 15528 4156
rect 15382 4111 15438 4120
rect 16316 4078 16344 6054
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 15304 3738 15332 4014
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 15212 2990 15240 3538
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 15200 2984 15252 2990
rect 15198 2952 15200 2961
rect 15384 2984 15436 2990
rect 15252 2952 15254 2961
rect 15384 2926 15436 2932
rect 15198 2887 15254 2896
rect 15396 2514 15424 2926
rect 16408 2553 16436 7534
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16500 5370 16528 6190
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16592 5302 16620 10095
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16684 7410 16712 7822
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16684 7206 16712 7346
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16684 6662 16712 7142
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16684 6322 16712 6598
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 16592 5098 16620 5238
rect 16776 5166 16804 12242
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 16868 11626 16896 12038
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 16960 11762 16988 11834
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 17420 11694 17448 12038
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 17408 11552 17460 11558
rect 17512 11506 17540 12174
rect 17696 11898 17724 12242
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17682 11792 17738 11801
rect 17682 11727 17684 11736
rect 17736 11727 17738 11736
rect 17684 11698 17736 11704
rect 17460 11500 17540 11506
rect 17408 11494 17540 11500
rect 17420 11478 17540 11494
rect 17420 10169 17448 11478
rect 17696 11370 17724 11698
rect 17604 11342 17724 11370
rect 17498 11248 17554 11257
rect 17498 11183 17554 11192
rect 17512 11150 17540 11183
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17512 10470 17540 11086
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17406 10160 17462 10169
rect 17406 10095 17462 10104
rect 17130 7032 17186 7041
rect 17130 6967 17186 6976
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17052 6254 17080 6598
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16868 5914 16896 6054
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 16960 5234 16988 5578
rect 17038 5400 17094 5409
rect 17038 5335 17094 5344
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16960 4690 16988 5170
rect 17052 4758 17080 5335
rect 17144 4826 17172 6967
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17236 5370 17264 5714
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17236 5273 17264 5306
rect 17222 5264 17278 5273
rect 17222 5199 17278 5208
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 17052 4282 17080 4694
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 17052 4049 17080 4218
rect 17144 4214 17172 4762
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17420 4282 17448 4626
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 17038 4040 17094 4049
rect 17038 3975 17094 3984
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16854 2952 16910 2961
rect 16854 2887 16910 2896
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16592 2666 16620 2790
rect 16500 2638 16620 2666
rect 16868 2650 16896 2887
rect 16856 2644 16908 2650
rect 16500 2582 16528 2638
rect 16856 2586 16908 2592
rect 16488 2576 16540 2582
rect 16394 2544 16450 2553
rect 15384 2508 15436 2514
rect 16488 2518 16540 2524
rect 16394 2479 16450 2488
rect 15384 2450 15436 2456
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 14002 2000 14058 2009
rect 14002 1935 14058 1944
rect 14752 1170 14780 2246
rect 15856 1170 15884 2246
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 14752 1142 14964 1170
rect 15856 1142 15976 1170
rect 14936 480 14964 1142
rect 15948 480 15976 1142
rect 16960 480 16988 3334
rect 17144 2961 17172 4150
rect 17512 3369 17540 10406
rect 17604 5914 17632 11342
rect 17880 11234 17908 19314
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17788 11206 17908 11234
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 17696 10985 17724 11154
rect 17682 10976 17738 10985
rect 17682 10911 17738 10920
rect 17696 10470 17724 10911
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17696 10033 17724 10406
rect 17682 10024 17738 10033
rect 17682 9959 17738 9968
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17604 5302 17632 5850
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17498 3360 17554 3369
rect 17498 3295 17554 3304
rect 17604 2990 17632 5238
rect 17788 4049 17816 11206
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17880 10810 17908 11086
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17972 8242 18000 11222
rect 17880 8214 18000 8242
rect 17880 5370 17908 8214
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17774 4040 17830 4049
rect 17774 3975 17830 3984
rect 17592 2984 17644 2990
rect 17130 2952 17186 2961
rect 17592 2926 17644 2932
rect 17130 2887 17186 2896
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 2650 17080 2790
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 18064 480 18092 20334
rect 18234 20295 18290 20304
rect 18248 20262 18276 20295
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18708 19378 18736 23520
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 19524 21004 19576 21010
rect 19524 20946 19576 20952
rect 19076 20262 19104 20946
rect 19430 20632 19486 20641
rect 19430 20567 19432 20576
rect 19484 20567 19486 20576
rect 19432 20538 19484 20544
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 19168 19446 19196 20334
rect 19536 20330 19564 20946
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19444 19922 19472 20198
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19156 19440 19208 19446
rect 19156 19382 19208 19388
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18418 13016 18474 13025
rect 18418 12951 18474 12960
rect 18432 11558 18460 12951
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18616 11762 18644 12174
rect 19062 11928 19118 11937
rect 19062 11863 19064 11872
rect 19116 11863 19118 11872
rect 19064 11834 19116 11840
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11286 18460 11494
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 18616 11150 18644 11698
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18142 9480 18198 9489
rect 18142 9415 18198 9424
rect 18156 7478 18184 9415
rect 19168 7562 19196 19382
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19076 7534 19196 7562
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18156 2514 18184 5034
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18144 2508 18196 2514
rect 18144 2450 18196 2456
rect 18432 921 18460 2790
rect 18510 2408 18566 2417
rect 18510 2343 18512 2352
rect 18564 2343 18566 2352
rect 18512 2314 18564 2320
rect 18418 912 18474 921
rect 18418 847 18474 856
rect 19076 480 19104 7534
rect 19260 3233 19288 19314
rect 19444 19174 19472 19858
rect 19614 19816 19670 19825
rect 19614 19751 19616 19760
rect 19668 19751 19670 19760
rect 19616 19722 19668 19728
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19340 18760 19392 18766
rect 19338 18728 19340 18737
rect 19392 18728 19394 18737
rect 19338 18663 19394 18672
rect 19338 12472 19394 12481
rect 19338 12407 19394 12416
rect 19352 4321 19380 12407
rect 19720 12322 19748 19110
rect 20180 12481 20208 23520
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21652 20602 21680 20946
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 20536 20528 20588 20534
rect 20534 20496 20536 20505
rect 20588 20496 20590 20505
rect 20534 20431 20590 20440
rect 21652 20330 21680 20538
rect 21744 20369 21772 23520
rect 23216 20641 23244 23520
rect 23202 20632 23258 20641
rect 23202 20567 23258 20576
rect 23848 20528 23900 20534
rect 23846 20496 23848 20505
rect 23900 20496 23902 20505
rect 23846 20431 23902 20440
rect 23664 20392 23716 20398
rect 21730 20360 21786 20369
rect 20720 20324 20772 20330
rect 20720 20266 20772 20272
rect 21640 20324 21692 20330
rect 21730 20295 21786 20304
rect 22006 20360 22062 20369
rect 23664 20334 23716 20340
rect 22006 20295 22062 20304
rect 22100 20324 22152 20330
rect 21640 20266 21692 20272
rect 20732 19922 20760 20266
rect 22020 20262 22048 20295
rect 22100 20266 22152 20272
rect 22008 20256 22060 20262
rect 22112 20233 22140 20266
rect 22376 20256 22428 20262
rect 22008 20198 22060 20204
rect 22098 20224 22154 20233
rect 20956 20156 21252 20176
rect 23676 20233 23704 20334
rect 22376 20198 22428 20204
rect 23662 20224 23718 20233
rect 22098 20159 22154 20168
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 21560 19961 21588 19994
rect 21546 19952 21602 19961
rect 20720 19916 20772 19922
rect 21546 19887 21602 19896
rect 20720 19858 20772 19864
rect 20732 19174 20760 19858
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20166 12472 20222 12481
rect 20166 12407 20222 12416
rect 19720 12294 19932 12322
rect 19904 4826 19932 12294
rect 19892 4820 19944 4826
rect 19892 4762 19944 4768
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 19338 4312 19394 4321
rect 19338 4247 19394 4256
rect 19614 3496 19670 3505
rect 19614 3431 19670 3440
rect 19246 3224 19302 3233
rect 19246 3159 19302 3168
rect 19628 2650 19656 3431
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 19430 2544 19486 2553
rect 19430 2479 19432 2488
rect 19484 2479 19486 2488
rect 19432 2450 19484 2456
rect 20088 480 20116 4762
rect 20732 1306 20760 19110
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 22006 14648 22062 14657
rect 22006 14583 22062 14592
rect 22020 14249 22048 14583
rect 22006 14240 22062 14249
rect 22006 14175 22062 14184
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 21914 13424 21970 13433
rect 21914 13359 21970 13368
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 21928 11218 21956 13359
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 22112 3534 22140 20159
rect 22100 3528 22152 3534
rect 22388 3482 22416 20198
rect 23662 20159 23718 20168
rect 24688 19825 24716 23520
rect 25410 23080 25466 23089
rect 25410 23015 25466 23024
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 24674 19816 24730 19825
rect 24674 19751 24730 19760
rect 25042 16144 25098 16153
rect 25042 16079 25098 16088
rect 24858 13424 24914 13433
rect 24858 13359 24914 13368
rect 24872 8945 24900 13359
rect 25056 10985 25084 16079
rect 25148 12753 25176 20402
rect 25318 20088 25374 20097
rect 25318 20023 25374 20032
rect 25226 17640 25282 17649
rect 25226 17575 25282 17584
rect 25134 12744 25190 12753
rect 25134 12679 25190 12688
rect 25042 10976 25098 10985
rect 25042 10911 25098 10920
rect 24858 8936 24914 8945
rect 24858 8871 24914 8880
rect 25240 7313 25268 17575
rect 25332 12209 25360 20023
rect 25424 13977 25452 23015
rect 25594 21584 25650 21593
rect 25594 21519 25650 21528
rect 25502 21312 25558 21321
rect 25502 21247 25558 21256
rect 25410 13968 25466 13977
rect 25410 13903 25466 13912
rect 25318 12200 25374 12209
rect 25318 12135 25374 12144
rect 25516 9489 25544 21247
rect 25608 21078 25636 21519
rect 25596 21072 25648 21078
rect 25596 21014 25648 21020
rect 25700 20312 25728 23559
rect 26238 23520 26294 24000
rect 27710 23520 27766 24000
rect 29182 23520 29238 24000
rect 26252 23474 26280 23520
rect 26252 23446 26464 23474
rect 25870 22400 25926 22409
rect 25870 22335 25926 22344
rect 25884 20466 25912 22335
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 25872 20460 25924 20466
rect 25872 20402 25924 20408
rect 25700 20284 25912 20312
rect 25778 20224 25834 20233
rect 25778 20159 25834 20168
rect 25686 19408 25742 19417
rect 25686 19343 25742 19352
rect 25594 15464 25650 15473
rect 25594 15399 25650 15408
rect 25502 9480 25558 9489
rect 25502 9415 25558 9424
rect 25226 7304 25282 7313
rect 25226 7239 25282 7248
rect 25608 5409 25636 15399
rect 25700 14521 25728 19343
rect 25792 14929 25820 20159
rect 25778 14920 25834 14929
rect 25778 14855 25834 14864
rect 25686 14512 25742 14521
rect 25686 14447 25742 14456
rect 25884 14090 25912 20284
rect 26436 19961 26464 23446
rect 27724 20369 27752 23520
rect 29196 20505 29224 23520
rect 29182 20496 29238 20505
rect 29182 20431 29238 20440
rect 27710 20360 27766 20369
rect 27710 20295 27766 20304
rect 26422 19952 26478 19961
rect 26422 19887 26478 19896
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 29366 18864 29422 18873
rect 29366 18799 29422 18808
rect 29380 18766 29408 18799
rect 29368 18760 29420 18766
rect 29368 18702 29420 18708
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 25700 14062 25912 14090
rect 25700 12889 25728 14062
rect 25778 13968 25834 13977
rect 25778 13903 25834 13912
rect 25686 12880 25742 12889
rect 25686 12815 25742 12824
rect 25792 11937 25820 13903
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 26422 12336 26478 12345
rect 26422 12271 26478 12280
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25778 11928 25834 11937
rect 25956 11920 26252 11940
rect 25778 11863 25834 11872
rect 26436 11694 26464 12271
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26606 11656 26662 11665
rect 26606 11591 26662 11600
rect 26620 11558 26648 11591
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 27344 11212 27396 11218
rect 27344 11154 27396 11160
rect 26698 11112 26754 11121
rect 26698 11047 26700 11056
rect 26752 11047 26754 11056
rect 26700 11018 26752 11024
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 27356 10810 27384 11154
rect 27344 10804 27396 10810
rect 27344 10746 27396 10752
rect 26424 10600 26476 10606
rect 26422 10568 26424 10577
rect 26476 10568 26478 10577
rect 26422 10503 26478 10512
rect 26608 10464 26660 10470
rect 26606 10432 26608 10441
rect 26660 10432 26662 10441
rect 26606 10367 26662 10376
rect 26698 9888 26754 9897
rect 25956 9820 26252 9840
rect 26698 9823 26754 9832
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 26514 9616 26570 9625
rect 26514 9551 26570 9560
rect 26422 9072 26478 9081
rect 26528 9042 26556 9551
rect 26606 9344 26662 9353
rect 26606 9279 26662 9288
rect 26422 9007 26478 9016
rect 26516 9036 26568 9042
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 26436 8430 26464 9007
rect 26516 8978 26568 8984
rect 26528 8634 26556 8978
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26620 8566 26648 9279
rect 26712 9178 26740 9823
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26698 8664 26754 8673
rect 26698 8599 26754 8608
rect 26608 8560 26660 8566
rect 26608 8502 26660 8508
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26712 8090 26740 8599
rect 27712 8560 27764 8566
rect 27526 8528 27582 8537
rect 27712 8502 27764 8508
rect 27526 8463 27582 8472
rect 27540 8430 27568 8463
rect 27528 8424 27580 8430
rect 27724 8401 27752 8502
rect 27528 8366 27580 8372
rect 27710 8392 27766 8401
rect 27710 8327 27766 8336
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 26514 7984 26570 7993
rect 26514 7919 26516 7928
rect 26568 7919 26570 7928
rect 26516 7890 26568 7896
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 26528 7546 26556 7890
rect 26790 7848 26846 7857
rect 26790 7783 26846 7792
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 26422 7440 26478 7449
rect 26422 7375 26478 7384
rect 26698 7440 26754 7449
rect 26698 7375 26754 7384
rect 26436 7342 26464 7375
rect 26424 7336 26476 7342
rect 26424 7278 26476 7284
rect 26608 7200 26660 7206
rect 26608 7142 26660 7148
rect 26620 7041 26648 7142
rect 26606 7032 26662 7041
rect 26606 6967 26662 6976
rect 26422 6896 26478 6905
rect 26422 6831 26478 6840
rect 26516 6860 26568 6866
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25594 5400 25650 5409
rect 25956 5392 26252 5412
rect 25594 5335 25650 5344
rect 26332 5024 26384 5030
rect 26332 4966 26384 4972
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 24582 4312 24638 4321
rect 25956 4304 26252 4324
rect 24582 4247 24638 4256
rect 22100 3470 22152 3476
rect 22204 3454 22416 3482
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 20732 1278 21128 1306
rect 21100 480 21128 1278
rect 22204 480 22232 3454
rect 23018 2816 23074 2825
rect 23018 2751 23074 2760
rect 23032 2650 23060 2751
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22848 2009 22876 2450
rect 22834 2000 22890 2009
rect 22834 1935 22890 1944
rect 23216 480 23244 3470
rect 24214 3088 24270 3097
rect 24214 3023 24270 3032
rect 24228 480 24256 3023
rect 24596 2514 24624 4247
rect 26344 4185 26372 4966
rect 26436 4690 26464 6831
rect 26516 6802 26568 6808
rect 26528 6254 26556 6802
rect 26712 6730 26740 7375
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26698 6352 26754 6361
rect 26698 6287 26754 6296
rect 26516 6248 26568 6254
rect 26514 6216 26516 6225
rect 26568 6216 26570 6225
rect 26514 6151 26570 6160
rect 26712 5914 26740 6287
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 26516 5772 26568 5778
rect 26516 5714 26568 5720
rect 26528 5166 26556 5714
rect 26606 5672 26662 5681
rect 26606 5607 26662 5616
rect 26620 5370 26648 5607
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26516 5160 26568 5166
rect 26514 5128 26516 5137
rect 26568 5128 26570 5137
rect 26514 5063 26570 5072
rect 26698 5128 26754 5137
rect 26698 5063 26754 5072
rect 26712 4826 26740 5063
rect 26700 4820 26752 4826
rect 26700 4762 26752 4768
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 26436 4282 26464 4626
rect 26606 4448 26662 4457
rect 26606 4383 26662 4392
rect 26424 4276 26476 4282
rect 26424 4218 26476 4224
rect 26330 4176 26386 4185
rect 26330 4111 26386 4120
rect 26424 4072 26476 4078
rect 25318 4040 25374 4049
rect 25318 3975 25374 3984
rect 25502 4040 25558 4049
rect 25502 3975 25558 3984
rect 26422 4040 26424 4049
rect 26476 4040 26478 4049
rect 26422 3975 26478 3984
rect 25332 3602 25360 3975
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25134 3224 25190 3233
rect 25332 3194 25360 3538
rect 25516 3369 25544 3975
rect 26620 3942 26648 4383
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26698 3904 26754 3913
rect 26698 3839 26754 3848
rect 26712 3738 26740 3839
rect 26700 3732 26752 3738
rect 26700 3674 26752 3680
rect 26804 3602 26832 7783
rect 27526 6488 27582 6497
rect 27526 6423 27582 6432
rect 26882 3632 26938 3641
rect 26792 3596 26844 3602
rect 26882 3567 26938 3576
rect 26792 3538 26844 3544
rect 26330 3496 26386 3505
rect 26330 3431 26386 3440
rect 25872 3392 25924 3398
rect 25502 3360 25558 3369
rect 25872 3334 25924 3340
rect 25502 3295 25558 3304
rect 25134 3159 25136 3168
rect 25188 3159 25190 3168
rect 25320 3188 25372 3194
rect 25136 3130 25188 3136
rect 25320 3130 25372 3136
rect 25148 2990 25176 3130
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 25502 2952 25558 2961
rect 25502 2887 25558 2896
rect 25516 2854 25544 2887
rect 25504 2848 25556 2854
rect 25226 2816 25282 2825
rect 25884 2825 25912 3334
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 25504 2790 25556 2796
rect 25870 2816 25926 2825
rect 25226 2751 25282 2760
rect 25870 2751 25926 2760
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24780 1601 24808 2246
rect 24766 1592 24822 1601
rect 24766 1527 24822 1536
rect 25240 480 25268 2751
rect 25688 2508 25740 2514
rect 25688 2450 25740 2456
rect 25700 1873 25728 2450
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25686 1864 25742 1873
rect 25686 1799 25742 1808
rect 3790 368 3846 377
rect 3790 303 3846 312
rect 4526 0 4582 480
rect 5630 0 5686 480
rect 6642 0 6698 480
rect 7654 0 7710 480
rect 8666 0 8722 480
rect 9770 0 9826 480
rect 10782 0 10838 480
rect 11794 0 11850 480
rect 12806 0 12862 480
rect 13910 0 13966 480
rect 14922 0 14978 480
rect 15934 0 15990 480
rect 16946 0 17002 480
rect 18050 0 18106 480
rect 19062 0 19118 480
rect 20074 0 20130 480
rect 21086 0 21142 480
rect 22190 0 22246 480
rect 23202 0 23258 480
rect 24214 0 24270 480
rect 25226 0 25282 480
rect 25884 377 25912 2246
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 26344 480 26372 3431
rect 26606 3360 26662 3369
rect 26606 3295 26662 3304
rect 26620 3194 26648 3295
rect 26804 3194 26832 3538
rect 26608 3188 26660 3194
rect 26608 3130 26660 3136
rect 26792 3188 26844 3194
rect 26792 3130 26844 3136
rect 26422 3088 26478 3097
rect 26422 3023 26478 3032
rect 26436 2990 26464 3023
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26896 2514 26924 3567
rect 27540 2990 27568 6423
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 28354 2952 28410 2961
rect 28354 2887 28410 2896
rect 27712 2848 27764 2854
rect 27342 2816 27398 2825
rect 27342 2751 27398 2760
rect 27710 2816 27712 2825
rect 27764 2816 27766 2825
rect 27710 2751 27766 2760
rect 26884 2508 26936 2514
rect 26884 2450 26936 2456
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 27080 1465 27108 2246
rect 27066 1456 27122 1465
rect 27066 1391 27122 1400
rect 27356 480 27384 2751
rect 28368 480 28396 2887
rect 29366 1592 29422 1601
rect 29366 1527 29422 1536
rect 29380 480 29408 1527
rect 25870 368 25926 377
rect 25870 303 25926 312
rect 26330 0 26386 480
rect 27342 0 27398 480
rect 28354 0 28410 480
rect 29366 0 29422 480
<< via2 >>
rect 4066 23568 4122 23624
rect 754 20304 810 20360
rect 3330 23024 3386 23080
rect 2870 22344 2926 22400
rect 2226 19760 2282 19816
rect 2686 13776 2742 13832
rect 2686 12708 2742 12744
rect 2686 12688 2688 12708
rect 2688 12688 2740 12708
rect 2740 12688 2742 12708
rect 1582 11600 1638 11656
rect 1398 11056 1454 11112
rect 1950 11328 2006 11384
rect 1766 11056 1822 11112
rect 1582 10376 1638 10432
rect 1398 9832 1454 9888
rect 1490 9288 1546 9344
rect 1582 8608 1638 8664
rect 1582 7420 1584 7440
rect 1584 7420 1636 7440
rect 1636 7420 1638 7440
rect 1582 7384 1638 7420
rect 1582 6840 1638 6896
rect 1582 5616 1638 5672
rect 1582 5072 1638 5128
rect 1582 4428 1584 4448
rect 1584 4428 1636 4448
rect 1636 4428 1638 4448
rect 1582 4392 1638 4428
rect 1582 3884 1584 3904
rect 1584 3884 1636 3904
rect 1636 3884 1638 3904
rect 1582 3848 1638 3884
rect 1398 1400 1454 1456
rect 2042 10668 2098 10704
rect 2042 10648 2044 10668
rect 2044 10648 2096 10668
rect 2096 10648 2098 10668
rect 3330 21800 3386 21856
rect 25686 23568 25742 23624
rect 3882 21256 3938 21312
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 4066 20032 4122 20088
rect 2962 18808 3018 18864
rect 2594 11756 2650 11792
rect 2594 11736 2596 11756
rect 2596 11736 2648 11756
rect 2648 11736 2650 11756
rect 2686 11056 2742 11112
rect 3422 16360 3478 16416
rect 3146 12144 3202 12200
rect 3054 10376 3110 10432
rect 2318 8336 2374 8392
rect 2410 7792 2466 7848
rect 2686 8064 2742 8120
rect 2686 7928 2742 7984
rect 2502 7384 2558 7440
rect 2134 7248 2190 7304
rect 2042 7148 2044 7168
rect 2044 7148 2096 7168
rect 2096 7148 2098 7168
rect 2042 7112 2098 7148
rect 2042 4972 2044 4992
rect 2044 4972 2096 4992
rect 2096 4972 2098 4992
rect 2042 4936 2098 4972
rect 2502 6860 2558 6896
rect 2502 6840 2504 6860
rect 2504 6840 2556 6860
rect 2556 6840 2558 6860
rect 2410 6704 2466 6760
rect 2410 4664 2466 4720
rect 2686 6296 2742 6352
rect 3238 11464 3294 11520
rect 3698 15272 3754 15328
rect 3606 14592 3662 14648
rect 3422 11192 3478 11248
rect 3514 10512 3570 10568
rect 3422 6976 3478 7032
rect 4066 15000 4122 15056
rect 4066 14048 4122 14104
rect 3974 13368 4030 13424
rect 3882 12824 3938 12880
rect 3882 11872 3938 11928
rect 3974 10240 4030 10296
rect 4526 11872 4582 11928
rect 4342 11328 4398 11384
rect 4894 11772 4896 11792
rect 4896 11772 4948 11792
rect 4948 11772 4950 11792
rect 4894 11736 4950 11772
rect 4618 10240 4674 10296
rect 3606 5888 3662 5944
rect 2778 5208 2834 5264
rect 1674 856 1730 912
rect 3882 5616 3938 5672
rect 2870 3340 2872 3360
rect 2872 3340 2924 3360
rect 2924 3340 2926 3360
rect 2870 3304 2926 3340
rect 3606 2896 3662 2952
rect 3330 2624 3386 2680
rect 3514 2644 3570 2680
rect 3514 2624 3516 2644
rect 3516 2624 3568 2644
rect 3568 2624 3570 2644
rect 2778 2080 2834 2136
rect 4434 5208 4490 5264
rect 4986 9968 5042 10024
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 5814 20576 5870 20632
rect 5354 18264 5410 18320
rect 5630 18264 5686 18320
rect 5078 9560 5134 9616
rect 4894 6840 4950 6896
rect 4710 5108 4712 5128
rect 4712 5108 4764 5128
rect 4764 5108 4766 5128
rect 4710 5072 4766 5108
rect 4066 3848 4122 3904
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 6274 18672 6330 18728
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 6090 10512 6146 10568
rect 5814 10104 5870 10160
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 5722 9560 5778 9616
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 6734 20440 6790 20496
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 8758 14456 8814 14512
rect 7838 13812 7840 13832
rect 7840 13812 7892 13832
rect 7892 13812 7894 13832
rect 7838 13776 7894 13812
rect 8482 13912 8538 13968
rect 7562 13096 7618 13152
rect 6734 9424 6790 9480
rect 6366 8336 6422 8392
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 6090 6296 6146 6352
rect 5722 5888 5778 5944
rect 6090 5908 6146 5944
rect 6090 5888 6092 5908
rect 6092 5888 6144 5908
rect 6144 5888 6146 5908
rect 5998 5616 6054 5672
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5354 5072 5410 5128
rect 5078 4936 5134 4992
rect 4986 4664 5042 4720
rect 6550 6432 6606 6488
rect 6734 4936 6790 4992
rect 5078 3732 5134 3768
rect 4526 2760 4582 2816
rect 5078 3712 5080 3732
rect 5080 3712 5132 3732
rect 5132 3712 5134 3732
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 4802 2488 4858 2544
rect 6274 3052 6330 3088
rect 6274 3032 6276 3052
rect 6276 3032 6328 3052
rect 6328 3032 6330 3052
rect 8390 10104 8446 10160
rect 8206 8492 8262 8528
rect 8206 8472 8208 8492
rect 8208 8472 8260 8492
rect 8260 8472 8262 8492
rect 8022 8336 8078 8392
rect 7562 7656 7618 7712
rect 7562 7248 7618 7304
rect 8298 6704 8354 6760
rect 7194 2624 7250 2680
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 7746 2760 7802 2816
rect 8298 2916 8354 2952
rect 8298 2896 8300 2916
rect 8300 2896 8352 2916
rect 8352 2896 8354 2916
rect 7930 2760 7986 2816
rect 9126 11500 9128 11520
rect 9128 11500 9180 11520
rect 9180 11500 9182 11520
rect 9126 11464 9182 11500
rect 9126 10240 9182 10296
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 9954 19896 10010 19952
rect 9310 17040 9366 17096
rect 9678 15816 9734 15872
rect 9494 13388 9550 13424
rect 9494 13368 9496 13388
rect 9496 13368 9548 13388
rect 9548 13368 9550 13388
rect 8942 8064 8998 8120
rect 9034 7792 9090 7848
rect 9126 7284 9128 7304
rect 9128 7284 9180 7304
rect 9180 7284 9182 7304
rect 9126 7248 9182 7284
rect 8850 7112 8906 7168
rect 9310 3984 9366 4040
rect 9678 11092 9680 11112
rect 9680 11092 9732 11112
rect 9732 11092 9734 11112
rect 9678 11056 9734 11092
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 10598 16632 10654 16688
rect 10230 15952 10286 16008
rect 9770 9968 9826 10024
rect 9770 7928 9826 7984
rect 9402 3712 9458 3768
rect 8850 3188 8906 3224
rect 8850 3168 8852 3188
rect 8852 3168 8904 3188
rect 8904 3168 8906 3188
rect 10506 14864 10562 14920
rect 10230 11056 10286 11112
rect 10138 9424 10194 9480
rect 10138 8880 10194 8936
rect 10138 8200 10194 8256
rect 10506 7792 10562 7848
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 10690 12824 10746 12880
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 12162 13132 12164 13152
rect 12164 13132 12216 13152
rect 12216 13132 12218 13152
rect 12162 13096 12218 13132
rect 10782 11600 10838 11656
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 10690 10648 10746 10704
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 10598 7520 10654 7576
rect 13450 12316 13452 12336
rect 13452 12316 13504 12336
rect 13504 12316 13506 12336
rect 13450 12280 13506 12316
rect 13174 12180 13176 12200
rect 13176 12180 13228 12200
rect 13228 12180 13230 12200
rect 13174 12144 13230 12180
rect 12990 11464 13046 11520
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 9862 6160 9918 6216
rect 12254 8608 12310 8664
rect 11426 6432 11482 6488
rect 11334 6296 11390 6352
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 9770 3984 9826 4040
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 11610 2760 11666 2816
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 13082 8900 13138 8936
rect 13082 8880 13084 8900
rect 13084 8880 13136 8900
rect 13136 8880 13138 8900
rect 12438 7248 12494 7304
rect 13082 7792 13138 7848
rect 12530 5616 12586 5672
rect 12346 3576 12402 3632
rect 13358 8492 13414 8528
rect 13358 8472 13360 8492
rect 13360 8472 13412 8492
rect 13412 8472 13414 8492
rect 13174 3168 13230 3224
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 15658 17176 15714 17232
rect 15474 15000 15530 15056
rect 14094 12844 14150 12880
rect 14094 12824 14096 12844
rect 14096 12824 14148 12844
rect 14148 12824 14150 12844
rect 14094 12180 14096 12200
rect 14096 12180 14148 12200
rect 14148 12180 14150 12200
rect 14094 12144 14150 12180
rect 13634 11056 13690 11112
rect 13634 7792 13690 7848
rect 13542 3168 13598 3224
rect 13634 3032 13690 3088
rect 13910 2760 13966 2816
rect 13358 2488 13414 2544
rect 13358 1808 13414 1864
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 16486 20304 16542 20360
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 17498 19780 17554 19816
rect 17498 19760 17500 19780
rect 17500 19760 17552 19780
rect 17552 19760 17554 19780
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 15566 8472 15622 8528
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 15750 10104 15806 10160
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 15750 9696 15806 9752
rect 16394 9016 16450 9072
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 15750 8472 15806 8528
rect 15106 7656 15162 7712
rect 15658 7520 15714 7576
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 16578 14184 16634 14240
rect 16578 10104 16634 10160
rect 15842 7248 15898 7304
rect 15658 6840 15714 6896
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 16210 5636 16266 5672
rect 16210 5616 16212 5636
rect 16212 5616 16264 5636
rect 16264 5616 16266 5636
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 16210 4700 16212 4720
rect 16212 4700 16264 4720
rect 16264 4700 16266 4720
rect 16210 4664 16266 4700
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 15382 4120 15438 4176
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 15198 2932 15200 2952
rect 15200 2932 15252 2952
rect 15252 2932 15254 2952
rect 15198 2896 15254 2932
rect 17682 11756 17738 11792
rect 17682 11736 17684 11756
rect 17684 11736 17736 11756
rect 17736 11736 17738 11756
rect 17498 11192 17554 11248
rect 17406 10104 17462 10160
rect 17130 6976 17186 7032
rect 17038 5344 17094 5400
rect 17222 5208 17278 5264
rect 17038 3984 17094 4040
rect 16854 2896 16910 2952
rect 16394 2488 16450 2544
rect 14002 1944 14058 2000
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 17682 10920 17738 10976
rect 17682 9968 17738 10024
rect 17498 3304 17554 3360
rect 17774 3984 17830 4040
rect 17130 2896 17186 2952
rect 18234 20304 18290 20360
rect 19430 20596 19486 20632
rect 19430 20576 19432 20596
rect 19432 20576 19484 20596
rect 19484 20576 19486 20596
rect 18418 12960 18474 13016
rect 19062 11892 19118 11928
rect 19062 11872 19064 11892
rect 19064 11872 19116 11892
rect 19116 11872 19118 11892
rect 18142 9424 18198 9480
rect 18510 2372 18566 2408
rect 18510 2352 18512 2372
rect 18512 2352 18564 2372
rect 18564 2352 18566 2372
rect 18418 856 18474 912
rect 19614 19780 19670 19816
rect 19614 19760 19616 19780
rect 19616 19760 19668 19780
rect 19668 19760 19670 19780
rect 19338 18708 19340 18728
rect 19340 18708 19392 18728
rect 19392 18708 19394 18728
rect 19338 18672 19394 18708
rect 19338 12416 19394 12472
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 20534 20476 20536 20496
rect 20536 20476 20588 20496
rect 20588 20476 20590 20496
rect 20534 20440 20590 20476
rect 23202 20576 23258 20632
rect 23846 20476 23848 20496
rect 23848 20476 23900 20496
rect 23900 20476 23902 20496
rect 23846 20440 23902 20476
rect 21730 20304 21786 20360
rect 22006 20304 22062 20360
rect 22098 20168 22154 20224
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 21546 19896 21602 19952
rect 20166 12416 20222 12472
rect 19338 4256 19394 4312
rect 19614 3440 19670 3496
rect 19246 3168 19302 3224
rect 19430 2508 19486 2544
rect 19430 2488 19432 2508
rect 19432 2488 19484 2508
rect 19484 2488 19486 2508
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 22006 14592 22062 14648
rect 22006 14184 22062 14240
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 21914 13368 21970 13424
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 23662 20168 23718 20224
rect 25410 23024 25466 23080
rect 24674 19760 24730 19816
rect 25042 16088 25098 16144
rect 24858 13368 24914 13424
rect 25318 20032 25374 20088
rect 25226 17584 25282 17640
rect 25134 12688 25190 12744
rect 25042 10920 25098 10976
rect 24858 8880 24914 8936
rect 25594 21528 25650 21584
rect 25502 21256 25558 21312
rect 25410 13912 25466 13968
rect 25318 12144 25374 12200
rect 25870 22344 25926 22400
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 25778 20168 25834 20224
rect 25686 19352 25742 19408
rect 25594 15408 25650 15464
rect 25502 9424 25558 9480
rect 25226 7248 25282 7304
rect 25778 14864 25834 14920
rect 25686 14456 25742 14512
rect 29182 20440 29238 20496
rect 27710 20304 27766 20360
rect 26422 19896 26478 19952
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 29366 18808 29422 18864
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 25778 13912 25834 13968
rect 25686 12824 25742 12880
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 26422 12280 26478 12336
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 25778 11872 25834 11928
rect 26606 11600 26662 11656
rect 26698 11076 26754 11112
rect 26698 11056 26700 11076
rect 26700 11056 26752 11076
rect 26752 11056 26754 11076
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 26422 10548 26424 10568
rect 26424 10548 26476 10568
rect 26476 10548 26478 10568
rect 26422 10512 26478 10548
rect 26606 10412 26608 10432
rect 26608 10412 26660 10432
rect 26660 10412 26662 10432
rect 26606 10376 26662 10412
rect 26698 9832 26754 9888
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 26514 9560 26570 9616
rect 26422 9016 26478 9072
rect 26606 9288 26662 9344
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 26698 8608 26754 8664
rect 27526 8472 27582 8528
rect 27710 8336 27766 8392
rect 26514 7948 26570 7984
rect 26514 7928 26516 7948
rect 26516 7928 26568 7948
rect 26568 7928 26570 7948
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 26790 7792 26846 7848
rect 26422 7384 26478 7440
rect 26698 7384 26754 7440
rect 26606 6976 26662 7032
rect 26422 6840 26478 6896
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 25594 5344 25650 5400
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 24582 4256 24638 4312
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 23018 2760 23074 2816
rect 22834 1944 22890 2000
rect 24214 3032 24270 3088
rect 26698 6296 26754 6352
rect 26514 6196 26516 6216
rect 26516 6196 26568 6216
rect 26568 6196 26570 6216
rect 26514 6160 26570 6196
rect 26606 5616 26662 5672
rect 26514 5108 26516 5128
rect 26516 5108 26568 5128
rect 26568 5108 26570 5128
rect 26514 5072 26570 5108
rect 26698 5072 26754 5128
rect 26606 4392 26662 4448
rect 26330 4120 26386 4176
rect 25318 3984 25374 4040
rect 25502 3984 25558 4040
rect 26422 4020 26424 4040
rect 26424 4020 26476 4040
rect 26476 4020 26478 4040
rect 26422 3984 26478 4020
rect 25134 3188 25190 3224
rect 26698 3848 26754 3904
rect 27526 6432 27582 6488
rect 26882 3576 26938 3632
rect 26330 3440 26386 3496
rect 25502 3304 25558 3360
rect 25134 3168 25136 3188
rect 25136 3168 25188 3188
rect 25188 3168 25190 3188
rect 25502 2896 25558 2952
rect 25226 2760 25282 2816
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 25870 2760 25926 2816
rect 24766 1536 24822 1592
rect 25686 1808 25742 1864
rect 3790 312 3846 368
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 26606 3304 26662 3360
rect 26422 3032 26478 3088
rect 28354 2896 28410 2952
rect 27342 2760 27398 2816
rect 27710 2796 27712 2816
rect 27712 2796 27764 2816
rect 27764 2796 27766 2816
rect 27710 2760 27766 2796
rect 27066 1400 27122 1456
rect 29366 1536 29422 1592
rect 25870 312 25926 368
<< metal3 >>
rect 0 23626 480 23656
rect 4061 23626 4127 23629
rect 0 23624 4127 23626
rect 0 23568 4066 23624
rect 4122 23568 4127 23624
rect 0 23566 4127 23568
rect 0 23536 480 23566
rect 4061 23563 4127 23566
rect 25681 23626 25747 23629
rect 29520 23626 30000 23656
rect 25681 23624 30000 23626
rect 25681 23568 25686 23624
rect 25742 23568 30000 23624
rect 25681 23566 30000 23568
rect 25681 23563 25747 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 3325 23082 3391 23085
rect 0 23080 3391 23082
rect 0 23024 3330 23080
rect 3386 23024 3391 23080
rect 0 23022 3391 23024
rect 0 22992 480 23022
rect 3325 23019 3391 23022
rect 25405 23082 25471 23085
rect 29520 23082 30000 23112
rect 25405 23080 30000 23082
rect 25405 23024 25410 23080
rect 25466 23024 30000 23080
rect 25405 23022 30000 23024
rect 25405 23019 25471 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 2865 22402 2931 22405
rect 0 22400 2931 22402
rect 0 22344 2870 22400
rect 2926 22344 2931 22400
rect 0 22342 2931 22344
rect 0 22312 480 22342
rect 2865 22339 2931 22342
rect 25865 22402 25931 22405
rect 29520 22402 30000 22432
rect 25865 22400 30000 22402
rect 25865 22344 25870 22400
rect 25926 22344 30000 22400
rect 25865 22342 30000 22344
rect 25865 22339 25931 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 3325 21858 3391 21861
rect 29520 21858 30000 21888
rect 0 21856 3391 21858
rect 0 21800 3330 21856
rect 3386 21800 3391 21856
rect 0 21798 3391 21800
rect 0 21768 480 21798
rect 3325 21795 3391 21798
rect 26374 21798 30000 21858
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 25589 21586 25655 21589
rect 26374 21586 26434 21798
rect 29520 21768 30000 21798
rect 25589 21584 26434 21586
rect 25589 21528 25594 21584
rect 25650 21528 26434 21584
rect 25589 21526 26434 21528
rect 25589 21523 25655 21526
rect 0 21314 480 21344
rect 3877 21314 3943 21317
rect 0 21312 3943 21314
rect 0 21256 3882 21312
rect 3938 21256 3943 21312
rect 0 21254 3943 21256
rect 0 21224 480 21254
rect 3877 21251 3943 21254
rect 25497 21314 25563 21317
rect 29520 21314 30000 21344
rect 25497 21312 30000 21314
rect 25497 21256 25502 21312
rect 25558 21256 30000 21312
rect 25497 21254 30000 21256
rect 25497 21251 25563 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 5809 20634 5875 20637
rect 0 20632 5875 20634
rect 0 20576 5814 20632
rect 5870 20576 5875 20632
rect 0 20574 5875 20576
rect 0 20544 480 20574
rect 5809 20571 5875 20574
rect 19425 20634 19491 20637
rect 23197 20634 23263 20637
rect 29520 20634 30000 20664
rect 19425 20632 23263 20634
rect 19425 20576 19430 20632
rect 19486 20576 23202 20632
rect 23258 20576 23263 20632
rect 19425 20574 23263 20576
rect 19425 20571 19491 20574
rect 23197 20571 23263 20574
rect 29318 20574 30000 20634
rect 6729 20498 6795 20501
rect 20529 20498 20595 20501
rect 6729 20496 20595 20498
rect 6729 20440 6734 20496
rect 6790 20440 20534 20496
rect 20590 20440 20595 20496
rect 6729 20438 20595 20440
rect 6729 20435 6795 20438
rect 20529 20435 20595 20438
rect 23841 20498 23907 20501
rect 29177 20498 29243 20501
rect 23841 20496 29243 20498
rect 23841 20440 23846 20496
rect 23902 20440 29182 20496
rect 29238 20440 29243 20496
rect 23841 20438 29243 20440
rect 23841 20435 23907 20438
rect 29177 20435 29243 20438
rect 749 20362 815 20365
rect 16481 20362 16547 20365
rect 749 20360 16547 20362
rect 749 20304 754 20360
rect 810 20304 16486 20360
rect 16542 20304 16547 20360
rect 749 20302 16547 20304
rect 749 20299 815 20302
rect 16481 20299 16547 20302
rect 18229 20362 18295 20365
rect 21725 20362 21791 20365
rect 18229 20360 21791 20362
rect 18229 20304 18234 20360
rect 18290 20304 21730 20360
rect 21786 20304 21791 20360
rect 18229 20302 21791 20304
rect 18229 20299 18295 20302
rect 21725 20299 21791 20302
rect 22001 20362 22067 20365
rect 27705 20362 27771 20365
rect 22001 20360 27771 20362
rect 22001 20304 22006 20360
rect 22062 20304 27710 20360
rect 27766 20304 27771 20360
rect 22001 20302 27771 20304
rect 22001 20299 22067 20302
rect 27705 20299 27771 20302
rect 22093 20226 22159 20229
rect 23657 20226 23723 20229
rect 22093 20224 23723 20226
rect 22093 20168 22098 20224
rect 22154 20168 23662 20224
rect 23718 20168 23723 20224
rect 22093 20166 23723 20168
rect 22093 20163 22159 20166
rect 23657 20163 23723 20166
rect 25773 20226 25839 20229
rect 29318 20226 29378 20574
rect 29520 20544 30000 20574
rect 25773 20224 29378 20226
rect 25773 20168 25778 20224
rect 25834 20168 29378 20224
rect 25773 20166 29378 20168
rect 25773 20163 25839 20166
rect 10944 20160 11264 20161
rect 0 20090 480 20120
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 4061 20090 4127 20093
rect 0 20088 4127 20090
rect 0 20032 4066 20088
rect 4122 20032 4127 20088
rect 0 20030 4127 20032
rect 0 20000 480 20030
rect 4061 20027 4127 20030
rect 25313 20090 25379 20093
rect 29520 20090 30000 20120
rect 25313 20088 30000 20090
rect 25313 20032 25318 20088
rect 25374 20032 30000 20088
rect 25313 20030 30000 20032
rect 25313 20027 25379 20030
rect 29520 20000 30000 20030
rect 9949 19954 10015 19957
rect 1350 19952 10015 19954
rect 1350 19896 9954 19952
rect 10010 19896 10015 19952
rect 1350 19894 10015 19896
rect 0 19410 480 19440
rect 1350 19410 1410 19894
rect 9949 19891 10015 19894
rect 21541 19954 21607 19957
rect 26417 19954 26483 19957
rect 21541 19952 26483 19954
rect 21541 19896 21546 19952
rect 21602 19896 26422 19952
rect 26478 19896 26483 19952
rect 21541 19894 26483 19896
rect 21541 19891 21607 19894
rect 26417 19891 26483 19894
rect 2221 19818 2287 19821
rect 17493 19818 17559 19821
rect 2221 19816 17559 19818
rect 2221 19760 2226 19816
rect 2282 19760 17498 19816
rect 17554 19760 17559 19816
rect 2221 19758 17559 19760
rect 2221 19755 2287 19758
rect 17493 19755 17559 19758
rect 19609 19818 19675 19821
rect 24669 19818 24735 19821
rect 19609 19816 24735 19818
rect 19609 19760 19614 19816
rect 19670 19760 24674 19816
rect 24730 19760 24735 19816
rect 19609 19758 24735 19760
rect 19609 19755 19675 19758
rect 24669 19755 24735 19758
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 0 19350 1410 19410
rect 25681 19410 25747 19413
rect 29520 19410 30000 19440
rect 25681 19408 30000 19410
rect 25681 19352 25686 19408
rect 25742 19352 30000 19408
rect 25681 19350 30000 19352
rect 0 19320 480 19350
rect 25681 19347 25747 19350
rect 29520 19320 30000 19350
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 0 18866 480 18896
rect 2957 18866 3023 18869
rect 0 18864 3023 18866
rect 0 18808 2962 18864
rect 3018 18808 3023 18864
rect 0 18806 3023 18808
rect 0 18776 480 18806
rect 2957 18803 3023 18806
rect 29361 18866 29427 18869
rect 29520 18866 30000 18896
rect 29361 18864 30000 18866
rect 29361 18808 29366 18864
rect 29422 18808 30000 18864
rect 29361 18806 30000 18808
rect 29361 18803 29427 18806
rect 29520 18776 30000 18806
rect 6269 18730 6335 18733
rect 19333 18730 19399 18733
rect 6269 18728 19399 18730
rect 6269 18672 6274 18728
rect 6330 18672 19338 18728
rect 19394 18672 19399 18728
rect 6269 18670 19399 18672
rect 6269 18667 6335 18670
rect 19333 18667 19399 18670
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 0 18322 480 18352
rect 5349 18322 5415 18325
rect 0 18320 5415 18322
rect 0 18264 5354 18320
rect 5410 18264 5415 18320
rect 0 18262 5415 18264
rect 0 18232 480 18262
rect 5349 18259 5415 18262
rect 5625 18322 5691 18325
rect 29520 18322 30000 18352
rect 5625 18320 11530 18322
rect 5625 18264 5630 18320
rect 5686 18264 11530 18320
rect 5625 18262 11530 18264
rect 5625 18259 5691 18262
rect 11470 18050 11530 18262
rect 29318 18262 30000 18322
rect 29318 18186 29378 18262
rect 29520 18232 30000 18262
rect 17174 18126 29378 18186
rect 17174 18050 17234 18126
rect 11470 17990 17234 18050
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 0 17642 480 17672
rect 25221 17642 25287 17645
rect 29520 17642 30000 17672
rect 0 17582 674 17642
rect 0 17552 480 17582
rect 614 17234 674 17582
rect 25221 17640 30000 17642
rect 25221 17584 25226 17640
rect 25282 17584 30000 17640
rect 25221 17582 30000 17584
rect 25221 17579 25287 17582
rect 29520 17552 30000 17582
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 15653 17234 15719 17237
rect 614 17232 15719 17234
rect 614 17176 15658 17232
rect 15714 17176 15719 17232
rect 614 17174 15719 17176
rect 15653 17171 15719 17174
rect 0 17098 480 17128
rect 9305 17098 9371 17101
rect 29520 17098 30000 17128
rect 0 17038 674 17098
rect 0 17008 480 17038
rect 614 16690 674 17038
rect 9305 17096 30000 17098
rect 9305 17040 9310 17096
rect 9366 17040 30000 17096
rect 9305 17038 30000 17040
rect 9305 17035 9371 17038
rect 29520 17008 30000 17038
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 10593 16690 10659 16693
rect 614 16688 10659 16690
rect 614 16632 10598 16688
rect 10654 16632 10659 16688
rect 614 16630 10659 16632
rect 10593 16627 10659 16630
rect 0 16418 480 16448
rect 3417 16418 3483 16421
rect 29520 16418 30000 16448
rect 0 16416 3483 16418
rect 0 16360 3422 16416
rect 3478 16360 3483 16416
rect 0 16358 3483 16360
rect 0 16328 480 16358
rect 3417 16355 3483 16358
rect 26558 16358 30000 16418
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 25037 16146 25103 16149
rect 26558 16146 26618 16358
rect 29520 16328 30000 16358
rect 25037 16144 26618 16146
rect 25037 16088 25042 16144
rect 25098 16088 26618 16144
rect 25037 16086 26618 16088
rect 25037 16083 25103 16086
rect 10225 16010 10291 16013
rect 10225 16008 29378 16010
rect 10225 15952 10230 16008
rect 10286 15952 29378 16008
rect 10225 15950 29378 15952
rect 10225 15947 10291 15950
rect 0 15874 480 15904
rect 9673 15874 9739 15877
rect 0 15872 9739 15874
rect 0 15816 9678 15872
rect 9734 15816 9739 15872
rect 0 15814 9739 15816
rect 29318 15874 29378 15950
rect 29520 15874 30000 15904
rect 29318 15814 30000 15874
rect 0 15784 480 15814
rect 9673 15811 9739 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 29520 15784 30000 15814
rect 20944 15743 21264 15744
rect 25589 15466 25655 15469
rect 25589 15464 26480 15466
rect 25589 15408 25594 15464
rect 25650 15408 26480 15464
rect 25589 15406 26480 15408
rect 25589 15403 25655 15406
rect 0 15330 480 15360
rect 3693 15330 3759 15333
rect 0 15328 3759 15330
rect 0 15272 3698 15328
rect 3754 15272 3759 15328
rect 0 15270 3759 15272
rect 26420 15330 26480 15406
rect 29520 15330 30000 15360
rect 26420 15270 30000 15330
rect 0 15240 480 15270
rect 3693 15267 3759 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 4061 15058 4127 15061
rect 15469 15058 15535 15061
rect 4061 15056 15535 15058
rect 4061 15000 4066 15056
rect 4122 15000 15474 15056
rect 15530 15000 15535 15056
rect 4061 14998 15535 15000
rect 4061 14995 4127 14998
rect 15469 14995 15535 14998
rect 10501 14922 10567 14925
rect 25773 14922 25839 14925
rect 10501 14920 25839 14922
rect 10501 14864 10506 14920
rect 10562 14864 25778 14920
rect 25834 14864 25839 14920
rect 10501 14862 25839 14864
rect 10501 14859 10567 14862
rect 25773 14859 25839 14862
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 3601 14650 3667 14653
rect 0 14648 3667 14650
rect 0 14592 3606 14648
rect 3662 14592 3667 14648
rect 0 14590 3667 14592
rect 0 14560 480 14590
rect 3601 14587 3667 14590
rect 22001 14650 22067 14653
rect 29520 14650 30000 14680
rect 22001 14648 30000 14650
rect 22001 14592 22006 14648
rect 22062 14592 30000 14648
rect 22001 14590 30000 14592
rect 22001 14587 22067 14590
rect 29520 14560 30000 14590
rect 8753 14514 8819 14517
rect 25681 14514 25747 14517
rect 8753 14512 25747 14514
rect 8753 14456 8758 14512
rect 8814 14456 25686 14512
rect 25742 14456 25747 14512
rect 8753 14454 25747 14456
rect 8753 14451 8819 14454
rect 25681 14451 25747 14454
rect 16573 14242 16639 14245
rect 22001 14242 22067 14245
rect 16573 14240 22067 14242
rect 16573 14184 16578 14240
rect 16634 14184 22006 14240
rect 22062 14184 22067 14240
rect 16573 14182 22067 14184
rect 16573 14179 16639 14182
rect 22001 14179 22067 14182
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 4061 14106 4127 14109
rect 29520 14106 30000 14136
rect 0 14104 4127 14106
rect 0 14048 4066 14104
rect 4122 14048 4127 14104
rect 0 14046 4127 14048
rect 0 14016 480 14046
rect 4061 14043 4127 14046
rect 26420 14046 30000 14106
rect 8477 13970 8543 13973
rect 25405 13970 25471 13973
rect 8477 13968 25471 13970
rect 8477 13912 8482 13968
rect 8538 13912 25410 13968
rect 25466 13912 25471 13968
rect 8477 13910 25471 13912
rect 8477 13907 8543 13910
rect 25405 13907 25471 13910
rect 25773 13970 25839 13973
rect 26420 13970 26480 14046
rect 29520 14016 30000 14046
rect 25773 13968 26480 13970
rect 25773 13912 25778 13968
rect 25834 13912 26480 13968
rect 25773 13910 26480 13912
rect 25773 13907 25839 13910
rect 2681 13834 2747 13837
rect 7833 13834 7899 13837
rect 2681 13832 7899 13834
rect 2681 13776 2686 13832
rect 2742 13776 7838 13832
rect 7894 13776 7899 13832
rect 2681 13774 7899 13776
rect 2681 13771 2747 13774
rect 7833 13771 7899 13774
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 0 13426 480 13456
rect 3969 13426 4035 13429
rect 0 13424 4035 13426
rect 0 13368 3974 13424
rect 4030 13368 4035 13424
rect 0 13366 4035 13368
rect 0 13336 480 13366
rect 3969 13363 4035 13366
rect 9489 13426 9555 13429
rect 21909 13426 21975 13429
rect 9489 13424 21975 13426
rect 9489 13368 9494 13424
rect 9550 13368 21914 13424
rect 21970 13368 21975 13424
rect 9489 13366 21975 13368
rect 9489 13363 9555 13366
rect 21909 13363 21975 13366
rect 24853 13426 24919 13429
rect 29520 13426 30000 13456
rect 24853 13424 30000 13426
rect 24853 13368 24858 13424
rect 24914 13368 30000 13424
rect 24853 13366 30000 13368
rect 24853 13363 24919 13366
rect 29520 13336 30000 13366
rect 7557 13154 7623 13157
rect 12157 13154 12223 13157
rect 7557 13152 12223 13154
rect 7557 13096 7562 13152
rect 7618 13096 12162 13152
rect 12218 13096 12223 13152
rect 7557 13094 12223 13096
rect 7557 13091 7623 13094
rect 12157 13091 12223 13094
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 18413 13018 18479 13021
rect 18413 13016 25882 13018
rect 18413 12960 18418 13016
rect 18474 12960 25882 13016
rect 18413 12958 25882 12960
rect 18413 12955 18479 12958
rect 0 12882 480 12912
rect 3877 12882 3943 12885
rect 0 12880 3943 12882
rect 0 12824 3882 12880
rect 3938 12824 3943 12880
rect 0 12822 3943 12824
rect 0 12792 480 12822
rect 3877 12819 3943 12822
rect 10685 12882 10751 12885
rect 14089 12882 14155 12885
rect 25681 12882 25747 12885
rect 10685 12880 25747 12882
rect 10685 12824 10690 12880
rect 10746 12824 14094 12880
rect 14150 12824 25686 12880
rect 25742 12824 25747 12880
rect 10685 12822 25747 12824
rect 25822 12882 25882 12958
rect 29520 12882 30000 12912
rect 25822 12822 30000 12882
rect 10685 12819 10751 12822
rect 14089 12819 14155 12822
rect 25681 12819 25747 12822
rect 29520 12792 30000 12822
rect 2681 12746 2747 12749
rect 25129 12746 25195 12749
rect 2681 12744 25195 12746
rect 2681 12688 2686 12744
rect 2742 12688 25134 12744
rect 25190 12688 25195 12744
rect 2681 12686 25195 12688
rect 2681 12683 2747 12686
rect 25129 12683 25195 12686
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 19333 12474 19399 12477
rect 20161 12474 20227 12477
rect 19333 12472 20227 12474
rect 19333 12416 19338 12472
rect 19394 12416 20166 12472
rect 20222 12416 20227 12472
rect 19333 12414 20227 12416
rect 19333 12411 19399 12414
rect 20161 12411 20227 12414
rect 0 12338 480 12368
rect 13445 12338 13511 12341
rect 26417 12338 26483 12341
rect 29520 12338 30000 12368
rect 0 12278 1778 12338
rect 0 12248 480 12278
rect 0 11658 480 11688
rect 1577 11658 1643 11661
rect 0 11656 1643 11658
rect 0 11600 1582 11656
rect 1638 11600 1643 11656
rect 0 11598 1643 11600
rect 0 11568 480 11598
rect 1577 11595 1643 11598
rect 1718 11250 1778 12278
rect 13445 12336 26483 12338
rect 13445 12280 13450 12336
rect 13506 12280 26422 12336
rect 26478 12280 26483 12336
rect 13445 12278 26483 12280
rect 13445 12275 13511 12278
rect 26417 12275 26483 12278
rect 27846 12278 30000 12338
rect 3141 12202 3207 12205
rect 13169 12202 13235 12205
rect 3141 12200 13235 12202
rect 3141 12144 3146 12200
rect 3202 12144 13174 12200
rect 13230 12144 13235 12200
rect 3141 12142 13235 12144
rect 3141 12139 3207 12142
rect 13169 12139 13235 12142
rect 14089 12202 14155 12205
rect 25313 12202 25379 12205
rect 14089 12200 25379 12202
rect 14089 12144 14094 12200
rect 14150 12144 25318 12200
rect 25374 12144 25379 12200
rect 14089 12142 25379 12144
rect 14089 12139 14155 12142
rect 25313 12139 25379 12142
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 3877 11930 3943 11933
rect 4521 11930 4587 11933
rect 19057 11930 19123 11933
rect 25773 11930 25839 11933
rect 3877 11928 5090 11930
rect 3877 11872 3882 11928
rect 3938 11872 4526 11928
rect 4582 11872 5090 11928
rect 3877 11870 5090 11872
rect 3877 11867 3943 11870
rect 4521 11867 4587 11870
rect 2589 11794 2655 11797
rect 4889 11794 4955 11797
rect 2589 11792 4955 11794
rect 2589 11736 2594 11792
rect 2650 11736 4894 11792
rect 4950 11736 4955 11792
rect 2589 11734 4955 11736
rect 5030 11794 5090 11870
rect 19057 11928 25839 11930
rect 19057 11872 19062 11928
rect 19118 11872 25778 11928
rect 25834 11872 25839 11928
rect 19057 11870 25839 11872
rect 19057 11867 19123 11870
rect 25773 11867 25839 11870
rect 17677 11794 17743 11797
rect 27846 11794 27906 12278
rect 29520 12248 30000 12278
rect 5030 11792 17743 11794
rect 5030 11736 17682 11792
rect 17738 11736 17743 11792
rect 5030 11734 17743 11736
rect 2589 11731 2655 11734
rect 4889 11731 4955 11734
rect 17677 11731 17743 11734
rect 17910 11734 27906 11794
rect 10777 11658 10843 11661
rect 10777 11656 11530 11658
rect 10777 11600 10782 11656
rect 10838 11600 11530 11656
rect 10777 11598 11530 11600
rect 10777 11595 10843 11598
rect 3233 11522 3299 11525
rect 9121 11522 9187 11525
rect 3233 11520 9187 11522
rect 3233 11464 3238 11520
rect 3294 11464 9126 11520
rect 9182 11464 9187 11520
rect 3233 11462 9187 11464
rect 11470 11522 11530 11598
rect 12985 11522 13051 11525
rect 17910 11522 17970 11734
rect 26601 11658 26667 11661
rect 29520 11658 30000 11688
rect 26601 11656 30000 11658
rect 26601 11600 26606 11656
rect 26662 11600 30000 11656
rect 26601 11598 30000 11600
rect 26601 11595 26667 11598
rect 29520 11568 30000 11598
rect 11470 11520 17970 11522
rect 11470 11464 12990 11520
rect 13046 11464 17970 11520
rect 11470 11462 17970 11464
rect 3233 11459 3299 11462
rect 9121 11459 9187 11462
rect 12985 11459 13051 11462
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 1945 11386 2011 11389
rect 4337 11386 4403 11389
rect 1945 11384 4403 11386
rect 1945 11328 1950 11384
rect 2006 11328 4342 11384
rect 4398 11328 4403 11384
rect 1945 11326 4403 11328
rect 1945 11323 2011 11326
rect 4337 11323 4403 11326
rect 3417 11250 3483 11253
rect 17493 11250 17559 11253
rect 1718 11190 3250 11250
rect 0 11114 480 11144
rect 1393 11114 1459 11117
rect 0 11112 1459 11114
rect 0 11056 1398 11112
rect 1454 11056 1459 11112
rect 0 11054 1459 11056
rect 0 11024 480 11054
rect 1393 11051 1459 11054
rect 1761 11114 1827 11117
rect 2681 11114 2747 11117
rect 1761 11112 2747 11114
rect 1761 11056 1766 11112
rect 1822 11056 2686 11112
rect 2742 11056 2747 11112
rect 1761 11054 2747 11056
rect 3190 11114 3250 11190
rect 3417 11248 17559 11250
rect 3417 11192 3422 11248
rect 3478 11192 17498 11248
rect 17554 11192 17559 11248
rect 3417 11190 17559 11192
rect 3417 11187 3483 11190
rect 17493 11187 17559 11190
rect 9673 11114 9739 11117
rect 3190 11112 9739 11114
rect 3190 11056 9678 11112
rect 9734 11056 9739 11112
rect 3190 11054 9739 11056
rect 1761 11051 1827 11054
rect 2681 11051 2747 11054
rect 9673 11051 9739 11054
rect 10225 11114 10291 11117
rect 13629 11114 13695 11117
rect 10225 11112 13695 11114
rect 10225 11056 10230 11112
rect 10286 11056 13634 11112
rect 13690 11056 13695 11112
rect 10225 11054 13695 11056
rect 10225 11051 10291 11054
rect 13629 11051 13695 11054
rect 26693 11114 26759 11117
rect 29520 11114 30000 11144
rect 26693 11112 30000 11114
rect 26693 11056 26698 11112
rect 26754 11056 30000 11112
rect 26693 11054 30000 11056
rect 26693 11051 26759 11054
rect 29520 11024 30000 11054
rect 17677 10978 17743 10981
rect 25037 10978 25103 10981
rect 17677 10976 25103 10978
rect 17677 10920 17682 10976
rect 17738 10920 25042 10976
rect 25098 10920 25103 10976
rect 17677 10918 25103 10920
rect 17677 10915 17743 10918
rect 25037 10915 25103 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 2037 10706 2103 10709
rect 10685 10706 10751 10709
rect 2037 10704 10751 10706
rect 2037 10648 2042 10704
rect 2098 10648 10690 10704
rect 10746 10648 10751 10704
rect 2037 10646 10751 10648
rect 2037 10643 2103 10646
rect 10685 10643 10751 10646
rect 3509 10570 3575 10573
rect 6085 10570 6151 10573
rect 26417 10570 26483 10573
rect 3509 10568 6151 10570
rect 3509 10512 3514 10568
rect 3570 10512 6090 10568
rect 6146 10512 6151 10568
rect 3509 10510 6151 10512
rect 3509 10507 3575 10510
rect 6085 10507 6151 10510
rect 6318 10568 26483 10570
rect 6318 10512 26422 10568
rect 26478 10512 26483 10568
rect 6318 10510 26483 10512
rect 0 10434 480 10464
rect 1577 10434 1643 10437
rect 0 10432 1643 10434
rect 0 10376 1582 10432
rect 1638 10376 1643 10432
rect 0 10374 1643 10376
rect 0 10344 480 10374
rect 1577 10371 1643 10374
rect 3049 10434 3115 10437
rect 6318 10434 6378 10510
rect 26417 10507 26483 10510
rect 3049 10432 6378 10434
rect 3049 10376 3054 10432
rect 3110 10376 6378 10432
rect 3049 10374 6378 10376
rect 26601 10434 26667 10437
rect 29520 10434 30000 10464
rect 26601 10432 30000 10434
rect 26601 10376 26606 10432
rect 26662 10376 30000 10432
rect 26601 10374 30000 10376
rect 3049 10371 3115 10374
rect 26601 10371 26667 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 3969 10298 4035 10301
rect 4613 10298 4679 10301
rect 9121 10298 9187 10301
rect 3969 10296 9187 10298
rect 3969 10240 3974 10296
rect 4030 10240 4618 10296
rect 4674 10240 9126 10296
rect 9182 10240 9187 10296
rect 3969 10238 9187 10240
rect 3969 10235 4035 10238
rect 4613 10235 4679 10238
rect 9121 10235 9187 10238
rect 5809 10162 5875 10165
rect 8385 10162 8451 10165
rect 5809 10160 8451 10162
rect 5809 10104 5814 10160
rect 5870 10104 8390 10160
rect 8446 10104 8451 10160
rect 5809 10102 8451 10104
rect 5809 10099 5875 10102
rect 8385 10099 8451 10102
rect 15745 10162 15811 10165
rect 16573 10162 16639 10165
rect 17401 10162 17467 10165
rect 15745 10160 17467 10162
rect 15745 10104 15750 10160
rect 15806 10104 16578 10160
rect 16634 10104 17406 10160
rect 17462 10104 17467 10160
rect 15745 10102 17467 10104
rect 15745 10099 15811 10102
rect 16573 10099 16639 10102
rect 17401 10099 17467 10102
rect 4981 10026 5047 10029
rect 9765 10026 9831 10029
rect 17677 10026 17743 10029
rect 4981 10024 6562 10026
rect 4981 9968 4986 10024
rect 5042 9968 6562 10024
rect 4981 9966 6562 9968
rect 4981 9963 5047 9966
rect 0 9890 480 9920
rect 1393 9890 1459 9893
rect 0 9888 1459 9890
rect 0 9832 1398 9888
rect 1454 9832 1459 9888
rect 0 9830 1459 9832
rect 0 9800 480 9830
rect 1393 9827 1459 9830
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 6502 9754 6562 9966
rect 9765 10024 17743 10026
rect 9765 9968 9770 10024
rect 9826 9968 17682 10024
rect 17738 9968 17743 10024
rect 9765 9966 17743 9968
rect 9765 9963 9831 9966
rect 17677 9963 17743 9966
rect 26693 9890 26759 9893
rect 29520 9890 30000 9920
rect 26693 9888 30000 9890
rect 26693 9832 26698 9888
rect 26754 9832 30000 9888
rect 26693 9830 30000 9832
rect 26693 9827 26759 9830
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 29520 9800 30000 9830
rect 25944 9759 26264 9760
rect 15745 9754 15811 9757
rect 6502 9752 15811 9754
rect 6502 9696 15750 9752
rect 15806 9696 15811 9752
rect 6502 9694 15811 9696
rect 15745 9691 15811 9694
rect 5073 9618 5139 9621
rect 5717 9618 5783 9621
rect 26509 9618 26575 9621
rect 5073 9616 26575 9618
rect 5073 9560 5078 9616
rect 5134 9560 5722 9616
rect 5778 9560 26514 9616
rect 26570 9560 26575 9616
rect 5073 9558 26575 9560
rect 5073 9555 5139 9558
rect 5717 9555 5783 9558
rect 26509 9555 26575 9558
rect 6729 9482 6795 9485
rect 10133 9482 10199 9485
rect 6729 9480 10199 9482
rect 6729 9424 6734 9480
rect 6790 9424 10138 9480
rect 10194 9424 10199 9480
rect 6729 9422 10199 9424
rect 6729 9419 6795 9422
rect 10133 9419 10199 9422
rect 18137 9482 18203 9485
rect 25497 9482 25563 9485
rect 18137 9480 25563 9482
rect 18137 9424 18142 9480
rect 18198 9424 25502 9480
rect 25558 9424 25563 9480
rect 18137 9422 25563 9424
rect 18137 9419 18203 9422
rect 25497 9419 25563 9422
rect 0 9346 480 9376
rect 1485 9346 1551 9349
rect 0 9344 1551 9346
rect 0 9288 1490 9344
rect 1546 9288 1551 9344
rect 0 9286 1551 9288
rect 0 9256 480 9286
rect 1485 9283 1551 9286
rect 26601 9346 26667 9349
rect 29520 9346 30000 9376
rect 26601 9344 30000 9346
rect 26601 9288 26606 9344
rect 26662 9288 30000 9344
rect 26601 9286 30000 9288
rect 26601 9283 26667 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 16389 9074 16455 9077
rect 26417 9074 26483 9077
rect 16389 9072 26483 9074
rect 16389 9016 16394 9072
rect 16450 9016 26422 9072
rect 26478 9016 26483 9072
rect 16389 9014 26483 9016
rect 16389 9011 16455 9014
rect 26417 9011 26483 9014
rect 10133 8938 10199 8941
rect 13077 8938 13143 8941
rect 24853 8938 24919 8941
rect 10133 8936 24919 8938
rect 10133 8880 10138 8936
rect 10194 8880 13082 8936
rect 13138 8880 24858 8936
rect 24914 8880 24919 8936
rect 10133 8878 24919 8880
rect 10133 8875 10199 8878
rect 13077 8875 13143 8878
rect 24853 8875 24919 8878
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 1577 8666 1643 8669
rect 12249 8666 12315 8669
rect 0 8664 1643 8666
rect 0 8608 1582 8664
rect 1638 8608 1643 8664
rect 9768 8664 12315 8666
rect 9768 8632 12254 8664
rect 0 8606 1643 8608
rect 0 8576 480 8606
rect 1577 8603 1643 8606
rect 9630 8608 12254 8632
rect 12310 8608 12315 8664
rect 9630 8606 12315 8608
rect 9630 8572 9828 8606
rect 12249 8603 12315 8606
rect 26693 8666 26759 8669
rect 29520 8666 30000 8696
rect 26693 8664 30000 8666
rect 26693 8608 26698 8664
rect 26754 8608 30000 8664
rect 26693 8606 30000 8608
rect 26693 8603 26759 8606
rect 29520 8576 30000 8606
rect 8201 8530 8267 8533
rect 9630 8530 9690 8572
rect 8201 8528 9690 8530
rect 8201 8472 8206 8528
rect 8262 8472 9690 8528
rect 8201 8470 9690 8472
rect 13353 8530 13419 8533
rect 15561 8530 15627 8533
rect 13353 8528 15627 8530
rect 13353 8472 13358 8528
rect 13414 8472 15566 8528
rect 15622 8472 15627 8528
rect 13353 8470 15627 8472
rect 8201 8467 8267 8470
rect 13353 8467 13419 8470
rect 15561 8467 15627 8470
rect 15745 8530 15811 8533
rect 27521 8530 27587 8533
rect 15745 8528 27587 8530
rect 15745 8472 15750 8528
rect 15806 8472 27526 8528
rect 27582 8472 27587 8528
rect 15745 8470 27587 8472
rect 15745 8467 15811 8470
rect 27521 8467 27587 8470
rect 2313 8394 2379 8397
rect 6361 8394 6427 8397
rect 2313 8392 6427 8394
rect 2313 8336 2318 8392
rect 2374 8336 6366 8392
rect 6422 8336 6427 8392
rect 2313 8334 6427 8336
rect 2313 8331 2379 8334
rect 6361 8331 6427 8334
rect 8017 8394 8083 8397
rect 27705 8394 27771 8397
rect 8017 8392 9690 8394
rect 8017 8336 8022 8392
rect 8078 8336 9690 8392
rect 8017 8334 9690 8336
rect 8017 8331 8083 8334
rect 9630 8292 9690 8334
rect 27705 8392 28642 8394
rect 27705 8336 27710 8392
rect 27766 8336 28642 8392
rect 27705 8334 28642 8336
rect 27705 8331 27771 8334
rect 9630 8258 10058 8292
rect 10133 8258 10199 8261
rect 9630 8256 10199 8258
rect 9630 8232 10138 8256
rect 9998 8200 10138 8232
rect 10194 8200 10199 8256
rect 9998 8198 10199 8200
rect 10133 8195 10199 8198
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 2681 8122 2747 8125
rect 0 8120 2747 8122
rect 0 8064 2686 8120
rect 2742 8064 2747 8120
rect 0 8062 2747 8064
rect 0 8032 480 8062
rect 2681 8059 2747 8062
rect 8937 8122 9003 8125
rect 28582 8122 28642 8334
rect 29520 8122 30000 8152
rect 8937 8120 10058 8122
rect 8937 8064 8942 8120
rect 8998 8064 10058 8120
rect 8937 8062 10058 8064
rect 28582 8062 30000 8122
rect 8937 8059 9003 8062
rect 2681 7986 2747 7989
rect 9765 7986 9831 7989
rect 2681 7984 9831 7986
rect 2681 7928 2686 7984
rect 2742 7928 9770 7984
rect 9826 7928 9831 7984
rect 2681 7926 9831 7928
rect 9998 7986 10058 8062
rect 29520 8032 30000 8062
rect 26509 7986 26575 7989
rect 9998 7984 26575 7986
rect 9998 7928 26514 7984
rect 26570 7928 26575 7984
rect 9998 7926 26575 7928
rect 2681 7923 2747 7926
rect 9765 7923 9831 7926
rect 26509 7923 26575 7926
rect 2405 7850 2471 7853
rect 9029 7850 9095 7853
rect 2405 7848 9095 7850
rect 2405 7792 2410 7848
rect 2466 7792 9034 7848
rect 9090 7792 9095 7848
rect 2405 7790 9095 7792
rect 2405 7787 2471 7790
rect 9029 7787 9095 7790
rect 10501 7850 10567 7853
rect 13077 7850 13143 7853
rect 10501 7848 13143 7850
rect 10501 7792 10506 7848
rect 10562 7792 13082 7848
rect 13138 7792 13143 7848
rect 10501 7790 13143 7792
rect 10501 7787 10567 7790
rect 13077 7787 13143 7790
rect 13629 7850 13695 7853
rect 26785 7850 26851 7853
rect 13629 7848 26851 7850
rect 13629 7792 13634 7848
rect 13690 7792 26790 7848
rect 26846 7792 26851 7848
rect 13629 7790 26851 7792
rect 13629 7787 13695 7790
rect 26785 7787 26851 7790
rect 7557 7714 7623 7717
rect 15101 7714 15167 7717
rect 7557 7712 15167 7714
rect 7557 7656 7562 7712
rect 7618 7656 15106 7712
rect 15162 7656 15167 7712
rect 7557 7654 15167 7656
rect 7557 7651 7623 7654
rect 15101 7651 15167 7654
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 10593 7578 10659 7581
rect 15653 7578 15719 7581
rect 10593 7576 15719 7578
rect 10593 7520 10598 7576
rect 10654 7520 15658 7576
rect 15714 7520 15719 7576
rect 10593 7518 15719 7520
rect 10593 7515 10659 7518
rect 15653 7515 15719 7518
rect 0 7442 480 7472
rect 1577 7442 1643 7445
rect 0 7440 1643 7442
rect 0 7384 1582 7440
rect 1638 7384 1643 7440
rect 0 7382 1643 7384
rect 0 7352 480 7382
rect 1577 7379 1643 7382
rect 2497 7442 2563 7445
rect 26417 7442 26483 7445
rect 2497 7440 26483 7442
rect 2497 7384 2502 7440
rect 2558 7384 26422 7440
rect 26478 7384 26483 7440
rect 2497 7382 26483 7384
rect 2497 7379 2563 7382
rect 26417 7379 26483 7382
rect 26693 7442 26759 7445
rect 29520 7442 30000 7472
rect 26693 7440 30000 7442
rect 26693 7384 26698 7440
rect 26754 7384 30000 7440
rect 26693 7382 30000 7384
rect 26693 7379 26759 7382
rect 29520 7352 30000 7382
rect 2129 7306 2195 7309
rect 7557 7306 7623 7309
rect 2129 7304 7623 7306
rect 2129 7248 2134 7304
rect 2190 7248 7562 7304
rect 7618 7248 7623 7304
rect 2129 7246 7623 7248
rect 2129 7243 2195 7246
rect 7557 7243 7623 7246
rect 9121 7306 9187 7309
rect 12433 7306 12499 7309
rect 9121 7304 12499 7306
rect 9121 7248 9126 7304
rect 9182 7248 12438 7304
rect 12494 7248 12499 7304
rect 9121 7246 12499 7248
rect 9121 7243 9187 7246
rect 12433 7243 12499 7246
rect 15837 7306 15903 7309
rect 25221 7306 25287 7309
rect 15837 7304 25287 7306
rect 15837 7248 15842 7304
rect 15898 7248 25226 7304
rect 25282 7248 25287 7304
rect 15837 7246 25287 7248
rect 15837 7243 15903 7246
rect 25221 7243 25287 7246
rect 2037 7170 2103 7173
rect 8845 7170 8911 7173
rect 2037 7168 8911 7170
rect 2037 7112 2042 7168
rect 2098 7112 8850 7168
rect 8906 7112 8911 7168
rect 2037 7110 8911 7112
rect 2037 7107 2103 7110
rect 8845 7107 8911 7110
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 3417 7034 3483 7037
rect 17125 7034 17191 7037
rect 3417 7032 10794 7034
rect 3417 6976 3422 7032
rect 3478 6976 10794 7032
rect 3417 6974 10794 6976
rect 3417 6971 3483 6974
rect 0 6898 480 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 480 6838
rect 1577 6835 1643 6838
rect 2497 6898 2563 6901
rect 4889 6898 4955 6901
rect 2497 6896 4955 6898
rect 2497 6840 2502 6896
rect 2558 6840 4894 6896
rect 4950 6840 4955 6896
rect 2497 6838 4955 6840
rect 10734 6898 10794 6974
rect 11470 7032 17191 7034
rect 11470 6976 17130 7032
rect 17186 6976 17191 7032
rect 11470 6974 17191 6976
rect 11470 6898 11530 6974
rect 17125 6971 17191 6974
rect 26601 7034 26667 7037
rect 26601 7032 26802 7034
rect 26601 6976 26606 7032
rect 26662 6976 26802 7032
rect 26601 6974 26802 6976
rect 26601 6971 26667 6974
rect 10734 6838 11530 6898
rect 15653 6898 15719 6901
rect 26417 6898 26483 6901
rect 15653 6896 26483 6898
rect 15653 6840 15658 6896
rect 15714 6840 26422 6896
rect 26478 6840 26483 6896
rect 15653 6838 26483 6840
rect 26742 6898 26802 6974
rect 29520 6898 30000 6928
rect 26742 6838 30000 6898
rect 2497 6835 2563 6838
rect 4889 6835 4955 6838
rect 15653 6835 15719 6838
rect 26417 6835 26483 6838
rect 29520 6808 30000 6838
rect 2405 6762 2471 6765
rect 8293 6762 8359 6765
rect 2405 6760 8359 6762
rect 2405 6704 2410 6760
rect 2466 6704 8298 6760
rect 8354 6704 8359 6760
rect 2405 6702 8359 6704
rect 2405 6699 2471 6702
rect 8293 6699 8359 6702
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 6545 6490 6611 6493
rect 11421 6490 11487 6493
rect 27521 6490 27587 6493
rect 6545 6488 11487 6490
rect 6545 6432 6550 6488
rect 6606 6432 11426 6488
rect 11482 6432 11487 6488
rect 6545 6430 11487 6432
rect 6545 6427 6611 6430
rect 11421 6427 11487 6430
rect 26558 6488 27587 6490
rect 26558 6432 27526 6488
rect 27582 6432 27587 6488
rect 26558 6430 27587 6432
rect 0 6354 480 6384
rect 2681 6354 2747 6357
rect 0 6352 2747 6354
rect 0 6296 2686 6352
rect 2742 6296 2747 6352
rect 0 6294 2747 6296
rect 0 6264 480 6294
rect 2681 6291 2747 6294
rect 6085 6354 6151 6357
rect 11329 6354 11395 6357
rect 26558 6354 26618 6430
rect 27521 6427 27587 6430
rect 6085 6352 26618 6354
rect 6085 6296 6090 6352
rect 6146 6296 11334 6352
rect 11390 6296 26618 6352
rect 6085 6294 26618 6296
rect 26693 6354 26759 6357
rect 29520 6354 30000 6384
rect 26693 6352 30000 6354
rect 26693 6296 26698 6352
rect 26754 6296 30000 6352
rect 26693 6294 30000 6296
rect 6085 6291 6151 6294
rect 11329 6291 11395 6294
rect 26693 6291 26759 6294
rect 29520 6264 30000 6294
rect 9857 6218 9923 6221
rect 26509 6218 26575 6221
rect 9857 6216 26575 6218
rect 9857 6160 9862 6216
rect 9918 6160 26514 6216
rect 26570 6160 26575 6216
rect 9857 6158 26575 6160
rect 9857 6155 9923 6158
rect 26509 6155 26575 6158
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 3601 5946 3667 5949
rect 5717 5946 5783 5949
rect 6085 5946 6151 5949
rect 3601 5944 6151 5946
rect 3601 5888 3606 5944
rect 3662 5888 5722 5944
rect 5778 5888 6090 5944
rect 6146 5888 6151 5944
rect 3601 5886 6151 5888
rect 3601 5883 3667 5886
rect 5717 5883 5783 5886
rect 6085 5883 6151 5886
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 3877 5674 3943 5677
rect 5993 5674 6059 5677
rect 3877 5672 6059 5674
rect 3877 5616 3882 5672
rect 3938 5616 5998 5672
rect 6054 5616 6059 5672
rect 3877 5614 6059 5616
rect 3877 5611 3943 5614
rect 5993 5611 6059 5614
rect 12525 5674 12591 5677
rect 16205 5674 16271 5677
rect 12525 5672 16271 5674
rect 12525 5616 12530 5672
rect 12586 5616 16210 5672
rect 16266 5616 16271 5672
rect 12525 5614 16271 5616
rect 12525 5611 12591 5614
rect 16205 5611 16271 5614
rect 26601 5674 26667 5677
rect 29520 5674 30000 5704
rect 26601 5672 30000 5674
rect 26601 5616 26606 5672
rect 26662 5616 30000 5672
rect 26601 5614 30000 5616
rect 26601 5611 26667 5614
rect 29520 5584 30000 5614
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 17033 5402 17099 5405
rect 25589 5402 25655 5405
rect 17033 5400 25655 5402
rect 17033 5344 17038 5400
rect 17094 5344 25594 5400
rect 25650 5344 25655 5400
rect 17033 5342 25655 5344
rect 17033 5339 17099 5342
rect 25589 5339 25655 5342
rect 2773 5266 2839 5269
rect 4429 5266 4495 5269
rect 17217 5266 17283 5269
rect 2773 5264 17283 5266
rect 2773 5208 2778 5264
rect 2834 5208 4434 5264
rect 4490 5208 17222 5264
rect 17278 5208 17283 5264
rect 2773 5206 17283 5208
rect 2773 5203 2839 5206
rect 4429 5203 4495 5206
rect 17217 5203 17283 5206
rect 0 5130 480 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 480 5070
rect 1577 5067 1643 5070
rect 4705 5130 4771 5133
rect 5349 5130 5415 5133
rect 26509 5130 26575 5133
rect 4705 5128 26575 5130
rect 4705 5072 4710 5128
rect 4766 5072 5354 5128
rect 5410 5072 26514 5128
rect 26570 5072 26575 5128
rect 4705 5070 26575 5072
rect 4705 5067 4771 5070
rect 5349 5067 5415 5070
rect 26509 5067 26575 5070
rect 26693 5130 26759 5133
rect 29520 5130 30000 5160
rect 26693 5128 30000 5130
rect 26693 5072 26698 5128
rect 26754 5072 30000 5128
rect 26693 5070 30000 5072
rect 26693 5067 26759 5070
rect 29520 5040 30000 5070
rect 2037 4994 2103 4997
rect 5073 4994 5139 4997
rect 6729 4994 6795 4997
rect 2037 4992 6795 4994
rect 2037 4936 2042 4992
rect 2098 4936 5078 4992
rect 5134 4936 6734 4992
rect 6790 4936 6795 4992
rect 2037 4934 6795 4936
rect 2037 4931 2103 4934
rect 5073 4931 5139 4934
rect 6729 4931 6795 4934
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 2405 4722 2471 4725
rect 4981 4722 5047 4725
rect 16205 4722 16271 4725
rect 2405 4720 16271 4722
rect 2405 4664 2410 4720
rect 2466 4664 4986 4720
rect 5042 4664 16210 4720
rect 16266 4664 16271 4720
rect 2405 4662 16271 4664
rect 2405 4659 2471 4662
rect 4981 4659 5047 4662
rect 16205 4659 16271 4662
rect 0 4450 480 4480
rect 1577 4450 1643 4453
rect 0 4448 1643 4450
rect 0 4392 1582 4448
rect 1638 4392 1643 4448
rect 0 4390 1643 4392
rect 0 4360 480 4390
rect 1577 4387 1643 4390
rect 26601 4450 26667 4453
rect 29520 4450 30000 4480
rect 26601 4448 30000 4450
rect 26601 4392 26606 4448
rect 26662 4392 30000 4448
rect 26601 4390 30000 4392
rect 26601 4387 26667 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 19333 4314 19399 4317
rect 24577 4314 24643 4317
rect 19333 4312 24643 4314
rect 19333 4256 19338 4312
rect 19394 4256 24582 4312
rect 24638 4256 24643 4312
rect 19333 4254 24643 4256
rect 19333 4251 19399 4254
rect 24577 4251 24643 4254
rect 15377 4178 15443 4181
rect 26325 4178 26391 4181
rect 15377 4176 26391 4178
rect 15377 4120 15382 4176
rect 15438 4120 26330 4176
rect 26386 4120 26391 4176
rect 15377 4118 26391 4120
rect 15377 4115 15443 4118
rect 26325 4115 26391 4118
rect 9305 4042 9371 4045
rect 9765 4042 9831 4045
rect 17033 4042 17099 4045
rect 9305 4040 9831 4042
rect 9305 3984 9310 4040
rect 9366 3984 9770 4040
rect 9826 3984 9831 4040
rect 9305 3982 9831 3984
rect 9305 3979 9371 3982
rect 9765 3979 9831 3982
rect 9998 4040 17099 4042
rect 9998 3984 17038 4040
rect 17094 3984 17099 4040
rect 9998 3982 17099 3984
rect 0 3906 480 3936
rect 1577 3906 1643 3909
rect 0 3904 1643 3906
rect 0 3848 1582 3904
rect 1638 3848 1643 3904
rect 0 3846 1643 3848
rect 0 3816 480 3846
rect 1577 3843 1643 3846
rect 4061 3906 4127 3909
rect 9998 3906 10058 3982
rect 17033 3979 17099 3982
rect 17769 4042 17835 4045
rect 25313 4042 25379 4045
rect 17769 4040 25379 4042
rect 17769 3984 17774 4040
rect 17830 3984 25318 4040
rect 25374 3984 25379 4040
rect 17769 3982 25379 3984
rect 17769 3979 17835 3982
rect 25313 3979 25379 3982
rect 25497 4042 25563 4045
rect 26417 4042 26483 4045
rect 25497 4040 26483 4042
rect 25497 3984 25502 4040
rect 25558 3984 26422 4040
rect 26478 3984 26483 4040
rect 25497 3982 26483 3984
rect 25497 3979 25563 3982
rect 26417 3979 26483 3982
rect 4061 3904 10058 3906
rect 4061 3848 4066 3904
rect 4122 3848 10058 3904
rect 4061 3846 10058 3848
rect 26693 3906 26759 3909
rect 29520 3906 30000 3936
rect 26693 3904 30000 3906
rect 26693 3848 26698 3904
rect 26754 3848 30000 3904
rect 26693 3846 30000 3848
rect 4061 3843 4127 3846
rect 26693 3843 26759 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 5073 3770 5139 3773
rect 9397 3770 9463 3773
rect 5073 3768 9463 3770
rect 5073 3712 5078 3768
rect 5134 3712 9402 3768
rect 9458 3712 9463 3768
rect 5073 3710 9463 3712
rect 5073 3707 5139 3710
rect 9397 3707 9463 3710
rect 12341 3634 12407 3637
rect 26877 3634 26943 3637
rect 12341 3632 26943 3634
rect 12341 3576 12346 3632
rect 12402 3576 26882 3632
rect 26938 3576 26943 3632
rect 12341 3574 26943 3576
rect 12341 3571 12407 3574
rect 26877 3571 26943 3574
rect 19609 3498 19675 3501
rect 26325 3498 26391 3501
rect 19609 3496 26391 3498
rect 19609 3440 19614 3496
rect 19670 3440 26330 3496
rect 26386 3440 26391 3496
rect 19609 3438 26391 3440
rect 19609 3435 19675 3438
rect 26325 3435 26391 3438
rect 0 3362 480 3392
rect 2865 3362 2931 3365
rect 0 3360 2931 3362
rect 0 3304 2870 3360
rect 2926 3304 2931 3360
rect 0 3302 2931 3304
rect 0 3272 480 3302
rect 2865 3299 2931 3302
rect 17493 3362 17559 3365
rect 25497 3362 25563 3365
rect 17493 3360 25563 3362
rect 17493 3304 17498 3360
rect 17554 3304 25502 3360
rect 25558 3304 25563 3360
rect 17493 3302 25563 3304
rect 17493 3299 17559 3302
rect 25497 3299 25563 3302
rect 26601 3362 26667 3365
rect 29520 3362 30000 3392
rect 26601 3360 30000 3362
rect 26601 3304 26606 3360
rect 26662 3304 30000 3360
rect 26601 3302 30000 3304
rect 26601 3299 26667 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 8845 3226 8911 3229
rect 13169 3226 13235 3229
rect 8845 3224 13235 3226
rect 8845 3168 8850 3224
rect 8906 3168 13174 3224
rect 13230 3168 13235 3224
rect 8845 3166 13235 3168
rect 8845 3163 8911 3166
rect 13169 3163 13235 3166
rect 13537 3226 13603 3229
rect 19241 3226 19307 3229
rect 25129 3226 25195 3229
rect 13537 3224 13922 3226
rect 13537 3168 13542 3224
rect 13598 3168 13922 3224
rect 13537 3166 13922 3168
rect 13537 3163 13603 3166
rect 6269 3090 6335 3093
rect 13629 3090 13695 3093
rect 6269 3088 13695 3090
rect 6269 3032 6274 3088
rect 6330 3032 13634 3088
rect 13690 3032 13695 3088
rect 6269 3030 13695 3032
rect 13862 3090 13922 3166
rect 19241 3224 25195 3226
rect 19241 3168 19246 3224
rect 19302 3168 25134 3224
rect 25190 3168 25195 3224
rect 19241 3166 25195 3168
rect 19241 3163 19307 3166
rect 25129 3163 25195 3166
rect 24209 3090 24275 3093
rect 26417 3090 26483 3093
rect 13862 3088 24275 3090
rect 13862 3032 24214 3088
rect 24270 3032 24275 3088
rect 13862 3030 24275 3032
rect 6269 3027 6335 3030
rect 13629 3027 13695 3030
rect 24209 3027 24275 3030
rect 24350 3088 26483 3090
rect 24350 3032 26422 3088
rect 26478 3032 26483 3088
rect 24350 3030 26483 3032
rect 3601 2954 3667 2957
rect 8293 2954 8359 2957
rect 15193 2954 15259 2957
rect 16849 2954 16915 2957
rect 3601 2952 8359 2954
rect 3601 2896 3606 2952
rect 3662 2896 8298 2952
rect 8354 2896 8359 2952
rect 3601 2894 8359 2896
rect 3601 2891 3667 2894
rect 8293 2891 8359 2894
rect 8526 2952 16915 2954
rect 8526 2896 15198 2952
rect 15254 2896 16854 2952
rect 16910 2896 16915 2952
rect 8526 2894 16915 2896
rect 4521 2818 4587 2821
rect 7741 2818 7807 2821
rect 4521 2816 7807 2818
rect 4521 2760 4526 2816
rect 4582 2760 7746 2816
rect 7802 2760 7807 2816
rect 4521 2758 7807 2760
rect 4521 2755 4587 2758
rect 7741 2755 7807 2758
rect 7925 2818 7991 2821
rect 8526 2818 8586 2894
rect 15193 2891 15259 2894
rect 16849 2891 16915 2894
rect 17125 2954 17191 2957
rect 24350 2954 24410 3030
rect 26417 3027 26483 3030
rect 17125 2952 24410 2954
rect 17125 2896 17130 2952
rect 17186 2896 24410 2952
rect 17125 2894 24410 2896
rect 25497 2954 25563 2957
rect 28349 2954 28415 2957
rect 25497 2952 28415 2954
rect 25497 2896 25502 2952
rect 25558 2896 28354 2952
rect 28410 2896 28415 2952
rect 25497 2894 28415 2896
rect 17125 2891 17191 2894
rect 25497 2891 25563 2894
rect 28349 2891 28415 2894
rect 7925 2816 8586 2818
rect 7925 2760 7930 2816
rect 7986 2760 8586 2816
rect 7925 2758 8586 2760
rect 11605 2818 11671 2821
rect 13905 2818 13971 2821
rect 11605 2816 13971 2818
rect 11605 2760 11610 2816
rect 11666 2760 13910 2816
rect 13966 2760 13971 2816
rect 11605 2758 13971 2760
rect 7925 2755 7991 2758
rect 11605 2755 11671 2758
rect 13905 2755 13971 2758
rect 23013 2818 23079 2821
rect 25221 2818 25287 2821
rect 23013 2816 25287 2818
rect 23013 2760 23018 2816
rect 23074 2760 25226 2816
rect 25282 2760 25287 2816
rect 23013 2758 25287 2760
rect 23013 2755 23079 2758
rect 25221 2755 25287 2758
rect 25865 2818 25931 2821
rect 27337 2818 27403 2821
rect 25865 2816 27403 2818
rect 25865 2760 25870 2816
rect 25926 2760 27342 2816
rect 27398 2760 27403 2816
rect 25865 2758 27403 2760
rect 25865 2755 25931 2758
rect 27337 2755 27403 2758
rect 27705 2818 27771 2821
rect 27705 2816 27906 2818
rect 27705 2760 27710 2816
rect 27766 2760 27906 2816
rect 27705 2758 27906 2760
rect 27705 2755 27771 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 3325 2682 3391 2685
rect 0 2680 3391 2682
rect 0 2624 3330 2680
rect 3386 2624 3391 2680
rect 0 2622 3391 2624
rect 0 2592 480 2622
rect 3325 2619 3391 2622
rect 3509 2682 3575 2685
rect 7189 2682 7255 2685
rect 3509 2680 7255 2682
rect 3509 2624 3514 2680
rect 3570 2624 7194 2680
rect 7250 2624 7255 2680
rect 3509 2622 7255 2624
rect 27846 2682 27906 2758
rect 29520 2682 30000 2712
rect 27846 2622 30000 2682
rect 3509 2619 3575 2622
rect 7189 2619 7255 2622
rect 29520 2592 30000 2622
rect 4797 2546 4863 2549
rect 13353 2546 13419 2549
rect 4797 2544 13419 2546
rect 4797 2488 4802 2544
rect 4858 2488 13358 2544
rect 13414 2488 13419 2544
rect 4797 2486 13419 2488
rect 4797 2483 4863 2486
rect 13353 2483 13419 2486
rect 16389 2546 16455 2549
rect 19425 2546 19491 2549
rect 16389 2544 19491 2546
rect 16389 2488 16394 2544
rect 16450 2488 19430 2544
rect 19486 2488 19491 2544
rect 16389 2486 19491 2488
rect 16389 2483 16455 2486
rect 19425 2483 19491 2486
rect 18505 2410 18571 2413
rect 18505 2408 27906 2410
rect 18505 2352 18510 2408
rect 18566 2352 27906 2408
rect 18505 2350 27906 2352
rect 18505 2347 18571 2350
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 27846 2138 27906 2350
rect 29520 2138 30000 2168
rect 27846 2078 30000 2138
rect 0 2048 480 2078
rect 2773 2075 2839 2078
rect 29520 2048 30000 2078
rect 13997 2002 14063 2005
rect 22829 2002 22895 2005
rect 13997 2000 22895 2002
rect 13997 1944 14002 2000
rect 14058 1944 22834 2000
rect 22890 1944 22895 2000
rect 13997 1942 22895 1944
rect 13997 1939 14063 1942
rect 22829 1939 22895 1942
rect 13353 1866 13419 1869
rect 25681 1866 25747 1869
rect 13353 1864 25747 1866
rect 13353 1808 13358 1864
rect 13414 1808 25686 1864
rect 25742 1808 25747 1864
rect 13353 1806 25747 1808
rect 13353 1803 13419 1806
rect 25681 1803 25747 1806
rect 24761 1594 24827 1597
rect 29361 1594 29427 1597
rect 24761 1592 29427 1594
rect 24761 1536 24766 1592
rect 24822 1536 29366 1592
rect 29422 1536 29427 1592
rect 24761 1534 29427 1536
rect 24761 1531 24827 1534
rect 29361 1531 29427 1534
rect 0 1458 480 1488
rect 1393 1458 1459 1461
rect 0 1456 1459 1458
rect 0 1400 1398 1456
rect 1454 1400 1459 1456
rect 0 1398 1459 1400
rect 0 1368 480 1398
rect 1393 1395 1459 1398
rect 27061 1458 27127 1461
rect 29520 1458 30000 1488
rect 27061 1456 30000 1458
rect 27061 1400 27066 1456
rect 27122 1400 30000 1456
rect 27061 1398 30000 1400
rect 27061 1395 27127 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 480 854
rect 1669 851 1735 854
rect 18413 914 18479 917
rect 29520 914 30000 944
rect 18413 912 30000 914
rect 18413 856 18418 912
rect 18474 856 30000 912
rect 18413 854 30000 856
rect 18413 851 18479 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 3785 370 3851 373
rect 0 368 3851 370
rect 0 312 3790 368
rect 3846 312 3851 368
rect 0 310 3851 312
rect 0 280 480 310
rect 3785 307 3851 310
rect 25865 370 25931 373
rect 29520 370 30000 400
rect 25865 368 30000 370
rect 25865 312 25870 368
rect 25926 312 30000 368
rect 25865 310 30000 312
rect 25865 307 25931 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
use sky130_fd_sc_hd__decap_3  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1840 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_14
timestamp 1604681595
transform 1 0 2392 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1604681595
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1932 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_19
timestamp 1604681595
transform 1 0 2852 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1604681595
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__15__A
timestamp 1604681595
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _15_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_41
timestamp 1604681595
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1604681595
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_34 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4232 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4600 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_49
timestamp 1604681595
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5060 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8004 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7452 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_79
timestamp 1604681595
transform 1 0 8372 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1604681595
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_93
timestamp 1604681595
transform 1 0 9660 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_85
timestamp 1604681595
transform 1 0 8924 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_104
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__1.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__1.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__1.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1604681595
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__2.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__2.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__3.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13064 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__3.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1604681595
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_139
timestamp 1604681595
transform 1 0 13892 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_127
timestamp 1604681595
transform 1 0 12788 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_150
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1604681595
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__5.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__4.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__5.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__4.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_1_174
timestamp 1604681595
transform 1 0 17112 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_170
timestamp 1604681595
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1604681595
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__5.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__4.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1604681595
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_176
timestamp 1604681595
transform 1 0 17296 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 18216 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_190
timestamp 1604681595
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_195
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 1604681595
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_207
timestamp 1604681595
transform 1 0 20148 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1604681595
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 19964 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_206
timestamp 1604681595
transform 1 0 20056 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_194
timestamp 1604681595
transform 1 0 18952 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_218
timestamp 1604681595
transform 1 0 21160 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_242
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_230
timestamp 1604681595
transform 1 0 22264 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_259
timestamp 1604681595
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_263
timestamp 1604681595
transform 1 0 25300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_267
timestamp 1604681595
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_279
timestamp 1604681595
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1604681595
transform 1 0 26036 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1604681595
transform 1 0 26404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_283
timestamp 1604681595
transform 1 0 27140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_288
timestamp 1604681595
transform 1 0 27600 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_284
timestamp 1604681595
transform 1 0 27232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1604681595
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 27416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 27508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_291
timestamp 1604681595
transform 1 0 27876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604681595
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp 1604681595
transform 1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1604681595
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1604681595
transform 1 0 2668 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_9
timestamp 1604681595
transform 1 0 1932 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4692 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_21
timestamp 1604681595
transform 1 0 3036 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_36
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_48
timestamp 1604681595
transform 1 0 5520 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_60
timestamp 1604681595
transform 1 0 6624 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_72
timestamp 1604681595
transform 1 0 7728 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1604681595
transform 1 0 10028 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1604681595
transform 1 0 10396 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_104
timestamp 1604681595
transform 1 0 10672 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__2.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11500 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_112
timestamp 1604681595
transform 1 0 11408 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__3.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_133
timestamp 1604681595
transform 1 0 13340 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 15824 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_158
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_164
timestamp 1604681595
transform 1 0 16192 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_176
timestamp 1604681595
transform 1 0 17296 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_188
timestamp 1604681595
transform 1 0 18400 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_200
timestamp 1604681595
transform 1 0 19504 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_267
timestamp 1604681595
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_280
timestamp 1604681595
transform 1 0 26864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_292
timestamp 1604681595
transform 1 0 27968 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1604681595
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__16__A
timestamp 1604681595
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_19
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1604681595
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1604681595
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_31
timestamp 1604681595
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1604681595
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_48
timestamp 1604681595
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_52
timestamp 1604681595
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_56
timestamp 1604681595
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1604681595
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_94
timestamp 1604681595
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_131
timestamp 1604681595
transform 1 0 13156 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_134
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_138
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1604681595
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15180 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_146
timestamp 1604681595
transform 1 0 14536 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1604681595
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1604681595
transform 1 0 16008 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_168
timestamp 1604681595
transform 1 0 16560 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604681595
transform 1 0 26404 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604681595
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1604681595
transform 1 0 27324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_279
timestamp 1604681595
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_283
timestamp 1604681595
transform 1 0 27140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_287
timestamp 1604681595
transform 1 0 27508 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1604681595
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1604681595
transform 1 0 2852 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4232 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5980 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_43
timestamp 1604681595
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_47
timestamp 1604681595
transform 1 0 5428 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_69
timestamp 1604681595
transform 1 0 7452 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_81
timestamp 1604681595
transform 1 0 8556 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1604681595
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_97
timestamp 1604681595
transform 1 0 10028 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_100
timestamp 1604681595
transform 1 0 10304 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_106
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_118
timestamp 1604681595
transform 1 0 11960 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_130
timestamp 1604681595
transform 1 0 13064 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_158
timestamp 1604681595
transform 1 0 15640 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16652 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_168
timestamp 1604681595
transform 1 0 16560 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_182
timestamp 1604681595
transform 1 0 17848 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_194
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604681595
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604681595
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1604681595
transform 1 0 26864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_292
timestamp 1604681595
transform 1 0 27968 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp 1604681595
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__17__A
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4324 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1604681595
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_31
timestamp 1604681595
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_48
timestamp 1604681595
transform 1 0 5520 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_55
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_102
timestamp 1604681595
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_106
timestamp 1604681595
transform 1 0 10856 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 13616 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_131
timestamp 1604681595
transform 1 0 13156 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_160
timestamp 1604681595
transform 1 0 15824 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1604681595
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1604681595
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1604681595
transform 1 0 26220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_279
timestamp 1604681595
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_283
timestamp 1604681595
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_295
timestamp 1604681595
transform 1 0 28244 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_7
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_17
timestamp 1604681595
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_11
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_19
timestamp 1604681595
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 3036 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1604681595
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_30
timestamp 1604681595
transform 1 0 3864 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_50
timestamp 1604681595
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_42
timestamp 1604681595
transform 1 0 4968 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_45
timestamp 1604681595
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_55
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_58
timestamp 1604681595
transform 1 0 6440 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_70
timestamp 1604681595
transform 1 0 7544 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_82
timestamp 1604681595
transform 1 0 8648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_66
timestamp 1604681595
transform 1 0 7176 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1604681595
transform 1 0 8280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_82
timestamp 1604681595
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604681595
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1604681595
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1604681595
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_97
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10304 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 8924 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_7_109
timestamp 1604681595
transform 1 0 11132 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_105
timestamp 1604681595
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_117
timestamp 1604681595
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_116
timestamp 1604681595
transform 1 0 11776 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12512 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 13708 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_140
timestamp 1604681595
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_144
timestamp 1604681595
transform 1 0 14352 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_127
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_153
timestamp 1604681595
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_150
timestamp 1604681595
transform 1 0 14904 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_161
timestamp 1604681595
transform 1 0 15916 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_157
timestamp 1604681595
transform 1 0 15548 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_163
timestamp 1604681595
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_168
timestamp 1604681595
transform 1 0 16560 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_180
timestamp 1604681595
transform 1 0 17664 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_173
timestamp 1604681595
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_177
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_192
timestamp 1604681595
transform 1 0 18768 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_204
timestamp 1604681595
transform 1 0 19872 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1604681595
transform 1 0 26496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_280
timestamp 1604681595
transform 1 0 26864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_275
timestamp 1604681595
transform 1 0 26404 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_278
timestamp 1604681595
transform 1 0 26680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_290
timestamp 1604681595
transform 1 0 27784 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_292
timestamp 1604681595
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1604681595
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_298
timestamp 1604681595
transform 1 0 28520 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1604681595
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6348 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 5980 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1604681595
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_50
timestamp 1604681595
transform 1 0 5704 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_73
timestamp 1604681595
transform 1 0 7820 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_81
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_110
timestamp 1604681595
transform 1 0 11224 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_118
timestamp 1604681595
transform 1 0 11960 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_132
timestamp 1604681595
transform 1 0 13248 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_136
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_139
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17020 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_167
timestamp 1604681595
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_171
timestamp 1604681595
transform 1 0 16836 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_175
timestamp 1604681595
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_187
timestamp 1604681595
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_199
timestamp 1604681595
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1604681595
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1604681595
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_292
timestamp 1604681595
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1604681595
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2944 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1604681595
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1604681595
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp 1604681595
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1604681595
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 7728 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8648 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1604681595
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_95
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_108
timestamp 1604681595
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1604681595
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1604681595
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1604681595
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_140
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_144
timestamp 1604681595
transform 1 0 14352 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15916 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_150
timestamp 1604681595
transform 1 0 14904 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_153
timestamp 1604681595
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_157
timestamp 1604681595
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 1604681595
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_174
timestamp 1604681595
transform 1 0 17112 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1604681595
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604681595
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1604681595
transform 1 0 26404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1604681595
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1604681595
transform 1 0 27324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_279
timestamp 1604681595
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1604681595
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_287
timestamp 1604681595
transform 1 0 27508 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_19
timestamp 1604681595
transform 1 0 2852 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_22
timestamp 1604681595
transform 1 0 3128 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1604681595
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_48
timestamp 1604681595
transform 1 0 5520 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _10_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7820 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 8096 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1604681595
transform 1 0 7084 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1604681595
transform 1 0 7452 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_72
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_101
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11040 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_121
timestamp 1604681595
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_125
timestamp 1604681595
transform 1 0 12604 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12696 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_135
timestamp 1604681595
transform 1 0 13524 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15824 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_147
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_169
timestamp 1604681595
transform 1 0 16652 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_181
timestamp 1604681595
transform 1 0 17756 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_193
timestamp 1604681595
transform 1 0 18860 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_205
timestamp 1604681595
transform 1 0 19964 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1604681595
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_292
timestamp 1604681595
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1604681595
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_19
timestamp 1604681595
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_23
timestamp 1604681595
transform 1 0 3220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1604681595
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp 1604681595
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_38
timestamp 1604681595
transform 1 0 4600 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 7544 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_73
timestamp 1604681595
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_81
timestamp 1604681595
transform 1 0 8556 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9200 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp 1604681595
transform 1 0 8924 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_108
timestamp 1604681595
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1604681595
transform 1 0 11500 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12696 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1604681595
transform 1 0 16100 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_166
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1604681595
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604681595
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1604681595
transform 1 0 26404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1604681595
transform 1 0 27508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1604681595
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1604681595
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_279
timestamp 1604681595
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_283
timestamp 1604681595
transform 1 0 27140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_291
timestamp 1604681595
transform 1 0 27876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1604681595
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1604681595
transform 1 0 28244 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_19
timestamp 1604681595
transform 1 0 2852 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp 1604681595
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_26
timestamp 1604681595
transform 1 0 3496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1604681595
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _06_
timestamp 1604681595
transform 1 0 5612 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_46
timestamp 1604681595
transform 1 0 5336 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_52
timestamp 1604681595
transform 1 0 5888 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_64
timestamp 1604681595
transform 1 0 6992 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_72
timestamp 1604681595
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_102
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11316 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_110
timestamp 1604681595
transform 1 0 11224 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1604681595
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_131
timestamp 1604681595
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_135
timestamp 1604681595
transform 1 0 13524 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_144
timestamp 1604681595
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1604681595
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_280
timestamp 1604681595
transform 1 0 26864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_292
timestamp 1604681595
transform 1 0 27968 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1604681595
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_9
timestamp 1604681595
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2300 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1604681595
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1604681595
transform 1 0 3496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1604681595
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1604681595
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_36
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_33
timestamp 1604681595
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4692 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp 1604681595
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1604681595
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_54
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1604681595
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_55
timestamp 1604681595
transform 1 0 6164 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_66
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_83
timestamp 1604681595
transform 1 0 8740 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_78
timestamp 1604681595
transform 1 0 8280 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1604681595
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1604681595
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1604681595
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_90
timestamp 1604681595
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1604681595
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_95
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_102
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_103
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1604681595
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_114
timestamp 1604681595
transform 1 0 11592 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_126
timestamp 1604681595
transform 1 0 12696 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_131
timestamp 1604681595
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_127
timestamp 1604681595
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_139
timestamp 1604681595
transform 1 0 13892 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14168 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_158
timestamp 1604681595
transform 1 0 15640 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_158
timestamp 1604681595
transform 1 0 15640 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_161
timestamp 1604681595
transform 1 0 15916 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_165
timestamp 1604681595
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_170
timestamp 1604681595
transform 1 0 16744 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1604681595
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_169
timestamp 1604681595
transform 1 0 16652 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_181
timestamp 1604681595
transform 1 0 17756 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_193
timestamp 1604681595
transform 1 0 18860 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1604681595
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1604681595
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_288
timestamp 1604681595
transform 1 0 27600 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1604681595
transform 1 0 28060 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_296
timestamp 1604681595
transform 1 0 28336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_28
timestamp 1604681595
transform 1 0 3680 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 1604681595
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_38
timestamp 1604681595
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_42
timestamp 1604681595
transform 1 0 4968 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_54
timestamp 1604681595
transform 1 0 6072 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1604681595
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1604681595
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_82
timestamp 1604681595
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9752 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1604681595
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_103
timestamp 1604681595
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1604681595
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_111
timestamp 1604681595
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_115
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1604681595
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13340 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_142
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_146
timestamp 1604681595
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_150
timestamp 1604681595
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_154
timestamp 1604681595
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_174
timestamp 1604681595
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_171
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_167
timestamp 1604681595
transform 1 0 16468 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1604681595
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_178
timestamp 1604681595
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17664 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_232
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1604681595
transform 1 0 26404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1604681595
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1604681595
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_279
timestamp 1604681595
transform 1 0 26772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_283
timestamp 1604681595
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_287
timestamp 1604681595
transform 1 0 27508 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_20
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_24
timestamp 1604681595
transform 1 0 3312 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1604681595
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1604681595
transform 1 0 5980 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_61
timestamp 1604681595
transform 1 0 6716 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_103
timestamp 1604681595
transform 1 0 10580 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_115
timestamp 1604681595
transform 1 0 11684 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13340 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_127
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1604681595
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15732 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_146
timestamp 1604681595
transform 1 0 14536 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1604681595
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_158
timestamp 1604681595
transform 1 0 15640 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17296 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_168
timestamp 1604681595
transform 1 0 16560 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_185
timestamp 1604681595
transform 1 0 18124 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_189
timestamp 1604681595
transform 1 0 18492 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1604681595
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_280
timestamp 1604681595
transform 1 0 26864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_292
timestamp 1604681595
transform 1 0 27968 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_298
timestamp 1604681595
transform 1 0 28520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_18
timestamp 1604681595
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_22
timestamp 1604681595
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_26
timestamp 1604681595
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_38
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_43
timestamp 1604681595
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_47
timestamp 1604681595
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_78
timestamp 1604681595
transform 1 0 8280 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9752 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_90
timestamp 1604681595
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_103
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_107
timestamp 1604681595
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_111
timestamp 1604681595
transform 1 0 11316 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_119
timestamp 1604681595
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_128
timestamp 1604681595
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_152
timestamp 1604681595
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_156
timestamp 1604681595
transform 1 0 15456 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1604681595
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1604681595
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_197
timestamp 1604681595
transform 1 0 19228 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_209
timestamp 1604681595
transform 1 0 20332 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_221
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_233
timestamp 1604681595
transform 1 0 22540 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_241
timestamp 1604681595
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1604681595
transform 1 0 26404 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1604681595
transform 1 0 26956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_279
timestamp 1604681595
transform 1 0 26772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_283
timestamp 1604681595
transform 1 0 27140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1604681595
transform 1 0 28244 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2300 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_11
timestamp 1604681595
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_22
timestamp 1604681595
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1604681595
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_40
timestamp 1604681595
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_57
timestamp 1604681595
transform 1 0 6348 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_63
timestamp 1604681595
transform 1 0 6900 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_66
timestamp 1604681595
transform 1 0 7176 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_74
timestamp 1604681595
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_77
timestamp 1604681595
transform 1 0 8188 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_83
timestamp 1604681595
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1604681595
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1604681595
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_107
timestamp 1604681595
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1604681595
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_123
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_131
timestamp 1604681595
transform 1 0 13156 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_135
timestamp 1604681595
transform 1 0 13524 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _09_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_157
timestamp 1604681595
transform 1 0 15548 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_165
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17388 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17204 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_168
timestamp 1604681595
transform 1 0 16560 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_174
timestamp 1604681595
transform 1 0 17112 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_186
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1604681595
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_288
timestamp 1604681595
transform 1 0 27600 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_296
timestamp 1604681595
transform 1 0 28336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_7
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_14
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 1604681595
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2208 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _07_
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_18
timestamp 1604681595
transform 1 0 2760 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1604681595
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_29
timestamp 1604681595
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_25
timestamp 1604681595
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1604681595
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4140 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_49
timestamp 1604681595
transform 1 0 5612 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_66
timestamp 1604681595
transform 1 0 7176 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_74
timestamp 1604681595
transform 1 0 7912 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1604681595
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_73
timestamp 1604681595
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8556 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_90
timestamp 1604681595
transform 1 0 9384 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_104
timestamp 1604681595
transform 1 0 10672 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_100
timestamp 1604681595
transform 1 0 10304 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_97
timestamp 1604681595
transform 1 0 10028 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_121
timestamp 1604681595
transform 1 0 12236 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13616 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1604681595
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1604681595
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_149
timestamp 1604681595
transform 1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_158
timestamp 1604681595
transform 1 0 15640 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_170
timestamp 1604681595
transform 1 0 16744 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1604681595
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_170
timestamp 1604681595
transform 1 0 16744 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_182
timestamp 1604681595
transform 1 0 17848 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_194
timestamp 1604681595
transform 1 0 18952 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_206
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_232
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1604681595
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1604681595
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_288
timestamp 1604681595
transform 1 0 27600 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1604681595
transform 1 0 28060 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_296
timestamp 1604681595
transform 1 0 28336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _08_
timestamp 1604681595
transform 1 0 6992 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_67
timestamp 1604681595
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_84
timestamp 1604681595
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1604681595
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_92
timestamp 1604681595
transform 1 0 9568 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_104
timestamp 1604681595
transform 1 0 10672 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_116
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1604681595
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1604681595
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1604681595
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1604681595
transform 1 0 26956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1604681595
transform 1 0 28060 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7728 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_81
timestamp 1604681595
transform 1 0 8556 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1604681595
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604681595
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1604681595
transform 1 0 27600 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_296
timestamp 1604681595
transform 1 0 28336 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1604681595
transform 1 0 26956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1604681595
transform 1 0 28060 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604681595
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_288
timestamp 1604681595
transform 1 0 27600 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_296
timestamp 1604681595
transform 1 0 28336 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1604681595
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1604681595
transform 1 0 26956 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1604681595
transform 1 0 28060 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_288
timestamp 1604681595
transform 1 0 27600 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1604681595
transform 1 0 26956 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_296
timestamp 1604681595
transform 1 0 28336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1604681595
transform 1 0 28060 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_288
timestamp 1604681595
transform 1 0 27600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1604681595
transform 1 0 28336 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1604681595
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1604681595
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1604681595
transform 1 0 26956 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1604681595
transform 1 0 28060 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_288
timestamp 1604681595
transform 1 0 27600 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1604681595
transform 1 0 28336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 17296 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1604681595
transform 1 0 17480 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1604681595
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_201
timestamp 1604681595
transform 1 0 19596 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_213
timestamp 1604681595
transform 1 0 20700 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_217
timestamp 1604681595
transform 1 0 21068 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1604681595
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_241
timestamp 1604681595
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1604681595
transform 1 0 26956 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1604681595
transform 1 0 28060 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 17296 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_174
timestamp 1604681595
transform 1 0 17112 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_180
timestamp 1604681595
transform 1 0 17664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_192
timestamp 1604681595
transform 1 0 18768 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_198
timestamp 1604681595
transform 1 0 19320 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_203
timestamp 1604681595
transform 1 0 19780 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_211
timestamp 1604681595
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_219
timestamp 1604681595
transform 1 0 21252 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_231
timestamp 1604681595
transform 1 0 22356 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_243
timestamp 1604681595
transform 1 0 23460 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_255
timestamp 1604681595
transform 1 0 24564 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_267
timestamp 1604681595
transform 1 0 25668 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_288
timestamp 1604681595
transform 1 0 27600 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_296
timestamp 1604681595
transform 1 0 28336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_80
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 10028 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_85
timestamp 1604681595
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_89
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_101
timestamp 1604681595
transform 1 0 10396 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1604681595
transform 1 0 11500 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1604681595
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_127
timestamp 1604681595
transform 1 0 12788 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_131
timestamp 1604681595
transform 1 0 13156 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_143
timestamp 1604681595
transform 1 0 14260 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 16284 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_155
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_163
timestamp 1604681595
transform 1 0 16100 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 18216 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_173
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_192
timestamp 1604681595
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_188
timestamp 1604681595
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1604681595
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_200
timestamp 1604681595
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 20056 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 19688 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 19320 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_213
timestamp 1604681595
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 20332 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_229
timestamp 1604681595
transform 1 0 22172 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 21620 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 21804 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 21620 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_233
timestamp 1604681595
transform 1 0 22540 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_241
timestamp 1604681595
transform 1 0 23276 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_249
timestamp 1604681595
transform 1 0 24012 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 24196 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_253
timestamp 1604681595
transform 1 0 24380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_265
timestamp 1604681595
transform 1 0 25484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_277
timestamp 1604681595
transform 1 0 26588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_289
timestamp 1604681595
transform 1 0 27692 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604681595
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 1604681595
transform 1 0 28428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604681595
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604681595
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604681595
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604681595
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604681595
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604681595
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604681595
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604681595
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604681595
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604681595
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604681595
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 9770 0 9826 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 9678 23520 9734 24000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 10782 0 10838 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 11242 23520 11298 24000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 478 0 534 480 6 bottom_grid_pin_0_
port 4 nsew default tristate
rlabel metal2 s 5630 0 5686 480 6 bottom_grid_pin_10_
port 5 nsew default tristate
rlabel metal2 s 1490 0 1546 480 6 bottom_grid_pin_2_
port 6 nsew default tristate
rlabel metal2 s 2502 0 2558 480 6 bottom_grid_pin_4_
port 7 nsew default tristate
rlabel metal2 s 3514 0 3570 480 6 bottom_grid_pin_6_
port 8 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 bottom_grid_pin_8_
port 9 nsew default tristate
rlabel metal2 s 6642 0 6698 480 6 ccff_head
port 10 nsew default input
rlabel metal2 s 7654 0 7710 480 6 ccff_tail
port 11 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 12 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 13 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 14 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 15 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 16 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 17 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 18 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 19 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 20 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 21 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 22 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 23 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 24 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 25 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 26 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 27 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 28 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 29 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 30 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 31 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 32 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 33 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 34 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 35 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 36 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 37 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 38 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 39 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 40 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 41 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 42 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 43 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 44 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 46 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 48 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 49 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 50 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 51 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 52 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 53 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 54 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 55 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 56 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 57 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 58 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 59 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 60 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 61 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 62 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 63 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 64 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 65 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 66 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 67 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 68 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 69 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 70 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 71 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 72 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 73 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 74 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 75 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 76 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 77 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 78 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 79 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 80 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 81 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 82 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 83 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 84 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 85 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 86 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 87 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 88 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 89 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 90 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 91 nsew default tristate
rlabel metal2 s 11794 0 11850 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
port 92 nsew default tristate
rlabel metal2 s 12806 0 12862 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
port 93 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
port 94 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
port 95 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
port 96 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
port 97 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[0]
port 98 nsew default input
rlabel metal2 s 19062 0 19118 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[1]
port 99 nsew default input
rlabel metal2 s 20074 0 20130 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[2]
port 100 nsew default input
rlabel metal2 s 21086 0 21142 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[3]
port 101 nsew default input
rlabel metal2 s 22190 0 22246 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[4]
port 102 nsew default input
rlabel metal2 s 23202 0 23258 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[5]
port 103 nsew default input
rlabel metal2 s 24214 0 24270 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
port 104 nsew default tristate
rlabel metal2 s 25226 0 25282 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
port 105 nsew default tristate
rlabel metal2 s 26330 0 26386 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
port 106 nsew default tristate
rlabel metal2 s 27342 0 27398 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
port 107 nsew default tristate
rlabel metal2 s 28354 0 28410 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
port 108 nsew default tristate
rlabel metal2 s 29366 0 29422 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
port 109 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 prog_clk
port 110 nsew default input
rlabel metal2 s 12714 23520 12770 24000 6 top_width_0_height_0__pin_0_
port 111 nsew default input
rlabel metal2 s 20166 23520 20222 24000 6 top_width_0_height_0__pin_10_
port 112 nsew default input
rlabel metal2 s 29182 23520 29238 24000 6 top_width_0_height_0__pin_11_lower
port 113 nsew default tristate
rlabel metal2 s 8206 23520 8262 24000 6 top_width_0_height_0__pin_11_upper
port 114 nsew default tristate
rlabel metal2 s 21730 23520 21786 24000 6 top_width_0_height_0__pin_1_lower
port 115 nsew default tristate
rlabel metal2 s 754 23520 810 24000 6 top_width_0_height_0__pin_1_upper
port 116 nsew default tristate
rlabel metal2 s 14186 23520 14242 24000 6 top_width_0_height_0__pin_2_
port 117 nsew default input
rlabel metal2 s 23202 23520 23258 24000 6 top_width_0_height_0__pin_3_lower
port 118 nsew default tristate
rlabel metal2 s 2226 23520 2282 24000 6 top_width_0_height_0__pin_3_upper
port 119 nsew default tristate
rlabel metal2 s 15750 23520 15806 24000 6 top_width_0_height_0__pin_4_
port 120 nsew default input
rlabel metal2 s 24674 23520 24730 24000 6 top_width_0_height_0__pin_5_lower
port 121 nsew default tristate
rlabel metal2 s 3698 23520 3754 24000 6 top_width_0_height_0__pin_5_upper
port 122 nsew default tristate
rlabel metal2 s 17222 23520 17278 24000 6 top_width_0_height_0__pin_6_
port 123 nsew default input
rlabel metal2 s 26238 23520 26294 24000 6 top_width_0_height_0__pin_7_lower
port 124 nsew default tristate
rlabel metal2 s 5170 23520 5226 24000 6 top_width_0_height_0__pin_7_upper
port 125 nsew default tristate
rlabel metal2 s 18694 23520 18750 24000 6 top_width_0_height_0__pin_8_
port 126 nsew default input
rlabel metal2 s 27710 23520 27766 24000 6 top_width_0_height_0__pin_9_lower
port 127 nsew default tristate
rlabel metal2 s 6734 23520 6790 24000 6 top_width_0_height_0__pin_9_upper
port 128 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 129 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 130 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
