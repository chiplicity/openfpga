VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__1_
  CLASS BLOCK ;
  FOREIGN sb_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.400 101.280 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 2.400 116.920 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 2.400 ;
    END
  END bottom_left_grid_pin_11_
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 2.400 ;
    END
  END bottom_left_grid_pin_15_
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN bottom_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END bottom_left_grid_pin_3_
  PIN bottom_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.400 ;
    END
  END bottom_left_grid_pin_5_
  PIN bottom_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 2.400 ;
    END
  END bottom_left_grid_pin_7_
  PIN bottom_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 2.400 ;
    END
  END bottom_left_grid_pin_9_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 2.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 73.480 140.000 74.080 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 80.280 140.000 80.880 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 87.080 140.000 87.680 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 93.880 140.000 94.480 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.360 140.000 101.960 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 108.160 140.000 108.760 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 114.960 140.000 115.560 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 122.440 140.000 123.040 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.240 140.000 129.840 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 10.240 140.000 10.840 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 17.040 140.000 17.640 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 23.840 140.000 24.440 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 31.320 140.000 31.920 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.120 140.000 38.720 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.920 140.000 45.520 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 52.400 140.000 53.000 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 59.200 140.000 59.800 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 66.000 140.000 66.600 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 137.600 44.070 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 137.600 49.130 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 137.600 54.190 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 137.600 59.250 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 137.600 64.770 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 137.600 74.890 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 137.600 79.950 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.190 137.600 85.470 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 137.600 90.530 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 137.600 95.590 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 137.600 100.650 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 137.600 106.170 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 137.600 111.230 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 137.600 116.290 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 137.600 121.350 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 137.600 126.870 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.650 137.600 131.930 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 2.400 132.560 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 2.400 8.120 ;
    END
  END enable
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 3.440 140.000 4.040 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.040 140.000 136.640 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 137.600 28.430 140.000 ;
    END
  END top_left_grid_pin_11_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 137.600 33.490 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 137.600 38.550 140.000 ;
    END
  END top_left_grid_pin_15_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 137.600 2.670 140.000 ;
    END
  END top_left_grid_pin_1_
  PIN top_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 137.600 7.730 140.000 ;
    END
  END top_left_grid_pin_3_
  PIN top_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 137.600 12.790 140.000 ;
    END
  END top_left_grid_pin_5_
  PIN top_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 137.600 17.850 140.000 ;
    END
  END top_left_grid_pin_7_
  PIN top_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 137.600 23.370 140.000 ;
    END
  END top_left_grid_pin_9_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.710 137.600 136.990 140.000 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 2.370 10.640 134.320 131.540 ;
      LAYER met2 ;
        RECT 2.950 137.320 7.170 137.600 ;
        RECT 8.010 137.320 12.230 137.600 ;
        RECT 13.070 137.320 17.290 137.600 ;
        RECT 18.130 137.320 22.810 137.600 ;
        RECT 23.650 137.320 27.870 137.600 ;
        RECT 28.710 137.320 32.930 137.600 ;
        RECT 33.770 137.320 37.990 137.600 ;
        RECT 38.830 137.320 43.510 137.600 ;
        RECT 44.350 137.320 48.570 137.600 ;
        RECT 49.410 137.320 53.630 137.600 ;
        RECT 54.470 137.320 58.690 137.600 ;
        RECT 59.530 137.320 64.210 137.600 ;
        RECT 65.050 137.320 69.270 137.600 ;
        RECT 70.110 137.320 74.330 137.600 ;
        RECT 75.170 137.320 79.390 137.600 ;
        RECT 80.230 137.320 84.910 137.600 ;
        RECT 85.750 137.320 89.970 137.600 ;
        RECT 90.810 137.320 95.030 137.600 ;
        RECT 95.870 137.320 100.090 137.600 ;
        RECT 100.930 137.320 105.610 137.600 ;
        RECT 106.450 137.320 110.670 137.600 ;
        RECT 111.510 137.320 115.730 137.600 ;
        RECT 116.570 137.320 120.790 137.600 ;
        RECT 121.630 137.320 126.310 137.600 ;
        RECT 127.150 137.320 131.370 137.600 ;
        RECT 132.210 137.320 136.430 137.600 ;
        RECT 2.390 2.680 136.990 137.320 ;
        RECT 2.950 2.400 7.170 2.680 ;
        RECT 8.010 2.400 12.230 2.680 ;
        RECT 13.070 2.400 17.290 2.680 ;
        RECT 18.130 2.400 22.810 2.680 ;
        RECT 23.650 2.400 27.870 2.680 ;
        RECT 28.710 2.400 32.930 2.680 ;
        RECT 33.770 2.400 37.990 2.680 ;
        RECT 38.830 2.400 43.510 2.680 ;
        RECT 44.350 2.400 48.570 2.680 ;
        RECT 49.410 2.400 53.630 2.680 ;
        RECT 54.470 2.400 58.690 2.680 ;
        RECT 59.530 2.400 64.210 2.680 ;
        RECT 65.050 2.400 69.270 2.680 ;
        RECT 70.110 2.400 74.330 2.680 ;
        RECT 75.170 2.400 79.390 2.680 ;
        RECT 80.230 2.400 84.910 2.680 ;
        RECT 85.750 2.400 89.970 2.680 ;
        RECT 90.810 2.400 95.030 2.680 ;
        RECT 95.870 2.400 100.090 2.680 ;
        RECT 100.930 2.400 105.610 2.680 ;
        RECT 106.450 2.400 110.670 2.680 ;
        RECT 111.510 2.400 115.730 2.680 ;
        RECT 116.570 2.400 120.790 2.680 ;
        RECT 121.630 2.400 126.310 2.680 ;
        RECT 127.150 2.400 131.370 2.680 ;
        RECT 132.210 2.400 136.430 2.680 ;
      LAYER met3 ;
        RECT 2.365 135.640 137.200 136.505 ;
        RECT 2.365 132.960 137.690 135.640 ;
        RECT 2.800 131.560 137.690 132.960 ;
        RECT 2.365 130.240 137.690 131.560 ;
        RECT 2.365 128.840 137.200 130.240 ;
        RECT 2.365 123.440 137.690 128.840 ;
        RECT 2.365 122.040 137.200 123.440 ;
        RECT 2.365 117.320 137.690 122.040 ;
        RECT 2.800 115.960 137.690 117.320 ;
        RECT 2.800 115.920 137.200 115.960 ;
        RECT 2.365 114.560 137.200 115.920 ;
        RECT 2.365 109.160 137.690 114.560 ;
        RECT 2.365 107.760 137.200 109.160 ;
        RECT 2.365 102.360 137.690 107.760 ;
        RECT 2.365 101.680 137.200 102.360 ;
        RECT 2.800 100.960 137.200 101.680 ;
        RECT 2.800 100.280 137.690 100.960 ;
        RECT 2.365 94.880 137.690 100.280 ;
        RECT 2.365 93.480 137.200 94.880 ;
        RECT 2.365 88.080 137.690 93.480 ;
        RECT 2.365 86.680 137.200 88.080 ;
        RECT 2.365 86.040 137.690 86.680 ;
        RECT 2.800 84.640 137.690 86.040 ;
        RECT 2.365 81.280 137.690 84.640 ;
        RECT 2.365 79.880 137.200 81.280 ;
        RECT 2.365 74.480 137.690 79.880 ;
        RECT 2.365 73.080 137.200 74.480 ;
        RECT 2.365 70.400 137.690 73.080 ;
        RECT 2.800 69.000 137.690 70.400 ;
        RECT 2.365 67.000 137.690 69.000 ;
        RECT 2.365 65.600 137.200 67.000 ;
        RECT 2.365 60.200 137.690 65.600 ;
        RECT 2.365 58.800 137.200 60.200 ;
        RECT 2.365 54.760 137.690 58.800 ;
        RECT 2.800 53.400 137.690 54.760 ;
        RECT 2.800 53.360 137.200 53.400 ;
        RECT 2.365 52.000 137.200 53.360 ;
        RECT 2.365 45.920 137.690 52.000 ;
        RECT 2.365 44.520 137.200 45.920 ;
        RECT 2.365 39.120 137.690 44.520 ;
        RECT 2.800 37.720 137.200 39.120 ;
        RECT 2.365 32.320 137.690 37.720 ;
        RECT 2.365 30.920 137.200 32.320 ;
        RECT 2.365 24.840 137.690 30.920 ;
        RECT 2.365 23.480 137.200 24.840 ;
        RECT 2.800 23.440 137.200 23.480 ;
        RECT 2.800 22.080 137.690 23.440 ;
        RECT 2.365 18.040 137.690 22.080 ;
        RECT 2.365 16.640 137.200 18.040 ;
        RECT 2.365 11.240 137.690 16.640 ;
        RECT 2.365 9.840 137.200 11.240 ;
        RECT 2.365 8.520 137.690 9.840 ;
        RECT 2.800 7.120 137.690 8.520 ;
        RECT 2.365 4.440 137.690 7.120 ;
        RECT 2.365 3.575 137.200 4.440 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_0__1_
END LIBRARY

