magic
tech EFS8A
magscale 1 2
timestamp 1602873556
<< locali >>
rect 15243 23137 15370 23171
rect 7975 19873 8010 19907
rect 6653 19261 6906 19295
rect 2881 19159 2915 19261
rect 6653 19227 6687 19261
rect 9631 18785 9758 18819
rect 19843 18785 19878 18819
rect 23155 18785 23190 18819
rect 6463 17833 6469 17867
rect 17687 17833 17693 17867
rect 19435 17833 19441 17867
rect 6463 17765 6497 17833
rect 17687 17765 17721 17833
rect 19435 17765 19469 17833
rect 14105 17085 14266 17119
rect 4546 17017 4616 17051
rect 19843 16609 19878 16643
rect 23983 16609 24110 16643
rect 16123 15657 16129 15691
rect 18239 15657 18245 15691
rect 9505 15351 9539 15657
rect 16123 15589 16157 15657
rect 18239 15589 18273 15657
rect 12449 14875 12483 15113
rect 4531 14807 4565 14875
rect 22103 14807 22137 14875
rect 4531 14773 4537 14807
rect 22103 14773 22109 14807
rect 4531 14569 4537 14603
rect 6463 14569 6469 14603
rect 4531 14501 4565 14569
rect 6463 14501 6497 14569
rect 9597 13719 9631 13821
rect 20085 13719 20119 14025
rect 22603 13821 22638 13855
rect 11983 12393 11989 12427
rect 21551 12393 21557 12427
rect 11983 12325 12017 12393
rect 21551 12325 21585 12393
rect 14841 10455 14875 10557
rect 21223 10149 21268 10183
rect 15243 10081 15323 10115
rect 25271 10081 25306 10115
rect 14933 9911 14967 10081
rect 24823 9673 24869 9707
rect 19901 9435 19935 9537
rect 24593 9469 24754 9503
rect 22695 8993 22730 9027
rect 9965 8279 9999 8449
rect 2455 7905 2490 7939
rect 21775 4641 21902 4675
<< viali >>
rect 24777 24837 24811 24871
rect 24593 24701 24627 24735
rect 25145 24701 25179 24735
rect 1593 24361 1627 24395
rect 17785 24361 17819 24395
rect 24777 24361 24811 24395
rect 1409 24225 1443 24259
rect 17601 24225 17635 24259
rect 23489 24225 23523 24259
rect 24593 24225 24627 24259
rect 23673 24089 23707 24123
rect 1961 23817 1995 23851
rect 13001 23817 13035 23851
rect 14565 23817 14599 23851
rect 16589 23817 16623 23851
rect 17601 23817 17635 23851
rect 19993 23817 20027 23851
rect 22017 23817 22051 23851
rect 23857 23817 23891 23851
rect 24777 23817 24811 23851
rect 1593 23749 1627 23783
rect 18889 23749 18923 23783
rect 25145 23681 25179 23715
rect 1409 23613 1443 23647
rect 12516 23613 12550 23647
rect 14080 23613 14114 23647
rect 16405 23613 16439 23647
rect 16957 23613 16991 23647
rect 18705 23613 18739 23647
rect 19257 23613 19291 23647
rect 19809 23613 19843 23647
rect 20361 23613 20395 23647
rect 21833 23613 21867 23647
rect 24593 23613 24627 23647
rect 22385 23545 22419 23579
rect 2421 23477 2455 23511
rect 12587 23477 12621 23511
rect 14151 23477 14185 23511
rect 24409 23477 24443 23511
rect 1593 23273 1627 23307
rect 11667 23273 11701 23307
rect 15439 23273 15473 23307
rect 23489 23273 23523 23307
rect 24777 23273 24811 23307
rect 1409 23137 1443 23171
rect 11564 23137 11598 23171
rect 15209 23137 15243 23171
rect 23305 23137 23339 23171
rect 24593 23137 24627 23171
rect 23305 22729 23339 22763
rect 24777 22729 24811 22763
rect 24409 22525 24443 22559
rect 24593 22525 24627 22559
rect 25145 22457 25179 22491
rect 1685 22389 1719 22423
rect 11529 22389 11563 22423
rect 15301 22389 15335 22423
rect 1476 22049 1510 22083
rect 2488 22049 2522 22083
rect 1547 21913 1581 21947
rect 2559 21845 2593 21879
rect 1593 21641 1627 21675
rect 24777 21641 24811 21675
rect 3065 21505 3099 21539
rect 1409 21437 1443 21471
rect 24593 21437 24627 21471
rect 25145 21437 25179 21471
rect 2421 21369 2455 21403
rect 1961 21301 1995 21335
rect 2513 21301 2547 21335
rect 1593 21097 1627 21131
rect 1409 20961 1443 20995
rect 2559 20961 2593 20995
rect 2651 20757 2685 20791
rect 1593 20553 1627 20587
rect 3341 20553 3375 20587
rect 24777 20553 24811 20587
rect 3065 20417 3099 20451
rect 1409 20349 1443 20383
rect 2580 20349 2614 20383
rect 3576 20349 3610 20383
rect 3985 20349 4019 20383
rect 9597 20349 9631 20383
rect 15060 20349 15094 20383
rect 15485 20349 15519 20383
rect 24593 20349 24627 20383
rect 25145 20349 25179 20383
rect 3663 20281 3697 20315
rect 2053 20213 2087 20247
rect 2421 20213 2455 20247
rect 2651 20213 2685 20247
rect 9781 20213 9815 20247
rect 10057 20213 10091 20247
rect 15163 20213 15197 20247
rect 1593 20009 1627 20043
rect 4215 20009 4249 20043
rect 5227 20009 5261 20043
rect 1409 19873 1443 19907
rect 2513 19873 2547 19907
rect 4144 19873 4178 19907
rect 5156 19873 5190 19907
rect 6964 19873 6998 19907
rect 7941 19873 7975 19907
rect 9724 19873 9758 19907
rect 10768 19873 10802 19907
rect 14232 19873 14266 19907
rect 15368 19873 15402 19907
rect 18061 19873 18095 19907
rect 18613 19873 18647 19907
rect 19660 19873 19694 19907
rect 18797 19805 18831 19839
rect 2697 19737 2731 19771
rect 14657 19737 14691 19771
rect 15439 19737 15473 19771
rect 20085 19737 20119 19771
rect 4629 19669 4663 19703
rect 7067 19669 7101 19703
rect 8079 19669 8113 19703
rect 9827 19669 9861 19703
rect 10839 19669 10873 19703
rect 14335 19669 14369 19703
rect 16221 19669 16255 19703
rect 19763 19669 19797 19703
rect 7665 19465 7699 19499
rect 8585 19465 8619 19499
rect 8953 19465 8987 19499
rect 10241 19465 10275 19499
rect 13645 19465 13679 19499
rect 17877 19465 17911 19499
rect 24777 19465 24811 19499
rect 7389 19329 7423 19363
rect 19441 19329 19475 19363
rect 1409 19261 1443 19295
rect 2580 19261 2614 19295
rect 2881 19261 2915 19295
rect 4261 19261 4295 19295
rect 4629 19261 4663 19295
rect 4905 19261 4939 19295
rect 8192 19261 8226 19295
rect 9781 19261 9815 19295
rect 10793 19261 10827 19295
rect 11412 19261 11446 19295
rect 11805 19261 11839 19295
rect 13461 19261 13495 19295
rect 14565 19261 14599 19295
rect 15025 19261 15059 19295
rect 18061 19261 18095 19295
rect 18613 19261 18647 19295
rect 19625 19261 19659 19295
rect 20085 19261 20119 19295
rect 24593 19261 24627 19295
rect 25145 19261 25179 19295
rect 1961 19193 1995 19227
rect 2973 19193 3007 19227
rect 6653 19193 6687 19227
rect 15301 19193 15335 19227
rect 16221 19193 16255 19227
rect 16313 19193 16347 19227
rect 16865 19193 16899 19227
rect 1593 19125 1627 19159
rect 2651 19125 2685 19159
rect 2881 19125 2915 19159
rect 3433 19125 3467 19159
rect 3893 19125 3927 19159
rect 4445 19125 4479 19159
rect 5365 19125 5399 19159
rect 6975 19125 7009 19159
rect 8263 19125 8297 19159
rect 9597 19125 9631 19159
rect 9965 19125 9999 19159
rect 11483 19125 11517 19159
rect 13369 19125 13403 19159
rect 14197 19125 14231 19159
rect 15577 19125 15611 19159
rect 16037 19125 16071 19159
rect 17509 19125 17543 19159
rect 18153 19125 18187 19159
rect 19073 19125 19107 19159
rect 19717 19125 19751 19159
rect 12449 18921 12483 18955
rect 18889 18921 18923 18955
rect 19717 18921 19751 18955
rect 23259 18921 23293 18955
rect 2513 18853 2547 18887
rect 4261 18853 4295 18887
rect 6929 18853 6963 18887
rect 16313 18853 16347 18887
rect 16405 18853 16439 18887
rect 16957 18853 16991 18887
rect 17877 18853 17911 18887
rect 17969 18853 18003 18887
rect 18521 18853 18555 18887
rect 21097 18853 21131 18887
rect 5784 18785 5818 18819
rect 8344 18785 8378 18819
rect 9597 18785 9631 18819
rect 11596 18785 11630 18819
rect 12633 18785 12667 18819
rect 13829 18785 13863 18819
rect 14197 18785 14231 18819
rect 19809 18785 19843 18819
rect 23121 18785 23155 18819
rect 2421 18717 2455 18751
rect 2697 18717 2731 18751
rect 4169 18717 4203 18751
rect 4629 18717 4663 18751
rect 5871 18717 5905 18751
rect 6285 18717 6319 18751
rect 6837 18717 6871 18751
rect 7481 18717 7515 18751
rect 14381 18717 14415 18751
rect 21005 18717 21039 18751
rect 21281 18717 21315 18751
rect 8769 18649 8803 18683
rect 1685 18581 1719 18615
rect 6561 18581 6595 18615
rect 8447 18581 8481 18615
rect 9827 18581 9861 18615
rect 10241 18581 10275 18615
rect 11667 18581 11701 18615
rect 12817 18581 12851 18615
rect 14657 18581 14691 18615
rect 15761 18581 15795 18615
rect 19947 18581 19981 18615
rect 2237 18377 2271 18411
rect 5273 18377 5307 18411
rect 6561 18377 6595 18411
rect 8309 18377 8343 18411
rect 9689 18377 9723 18411
rect 16681 18377 16715 18411
rect 16957 18377 16991 18411
rect 17509 18377 17543 18411
rect 21005 18377 21039 18411
rect 24777 18377 24811 18411
rect 3433 18309 3467 18343
rect 4905 18309 4939 18343
rect 22109 18309 22143 18343
rect 2421 18241 2455 18275
rect 3065 18241 3099 18275
rect 10333 18241 10367 18275
rect 10701 18241 10735 18275
rect 12541 18241 12575 18275
rect 18429 18241 18463 18275
rect 19349 18241 19383 18275
rect 21465 18241 21499 18275
rect 23121 18241 23155 18275
rect 5784 18173 5818 18207
rect 6285 18173 6319 18207
rect 8493 18173 8527 18207
rect 9413 18173 9447 18207
rect 10057 18173 10091 18207
rect 12173 18173 12207 18207
rect 14105 18173 14139 18207
rect 14381 18173 14415 18207
rect 14749 18173 14783 18207
rect 15761 18173 15795 18207
rect 19073 18173 19107 18207
rect 24593 18173 24627 18207
rect 25145 18173 25179 18207
rect 1869 18105 1903 18139
rect 2513 18105 2547 18139
rect 3985 18105 4019 18139
rect 4077 18105 4111 18139
rect 4629 18105 4663 18139
rect 5871 18105 5905 18139
rect 6929 18105 6963 18139
rect 7021 18105 7055 18139
rect 7573 18105 7607 18139
rect 8814 18105 8848 18139
rect 10425 18105 10459 18139
rect 12633 18105 12667 18139
rect 13185 18105 13219 18139
rect 13737 18105 13771 18139
rect 14933 18105 14967 18139
rect 16082 18105 16116 18139
rect 18521 18105 18555 18139
rect 19901 18105 19935 18139
rect 21189 18105 21223 18139
rect 21281 18105 21315 18139
rect 3801 18037 3835 18071
rect 7941 18037 7975 18071
rect 11621 18037 11655 18071
rect 15577 18037 15611 18071
rect 17785 18037 17819 18071
rect 20085 18037 20119 18071
rect 20545 18037 20579 18071
rect 2973 17833 3007 17867
rect 5181 17833 5215 17867
rect 6469 17833 6503 17867
rect 7665 17833 7699 17867
rect 9781 17833 9815 17867
rect 10885 17833 10919 17867
rect 14473 17833 14507 17867
rect 16589 17833 16623 17867
rect 17693 17833 17727 17867
rect 18245 17833 18279 17867
rect 18521 17833 18555 17867
rect 18981 17833 19015 17867
rect 19441 17833 19475 17867
rect 21925 17833 21959 17867
rect 24777 17833 24811 17867
rect 2145 17765 2179 17799
rect 4582 17765 4616 17799
rect 7297 17765 7331 17799
rect 8217 17765 8251 17799
rect 11615 17765 11649 17799
rect 13185 17765 13219 17799
rect 15755 17765 15789 17799
rect 21097 17765 21131 17799
rect 22661 17765 22695 17799
rect 23213 17765 23247 17799
rect 7021 17697 7055 17731
rect 9781 17697 9815 17731
rect 10149 17697 10183 17731
rect 16313 17697 16347 17731
rect 17325 17697 17359 17731
rect 19073 17697 19107 17731
rect 19993 17697 20027 17731
rect 24593 17697 24627 17731
rect 1869 17629 1903 17663
rect 2053 17629 2087 17663
rect 4261 17629 4295 17663
rect 6101 17629 6135 17663
rect 8125 17629 8159 17663
rect 11253 17629 11287 17663
rect 13093 17629 13127 17663
rect 13737 17629 13771 17663
rect 15393 17629 15427 17663
rect 21005 17629 21039 17663
rect 21465 17629 21499 17663
rect 22569 17629 22603 17663
rect 2605 17561 2639 17595
rect 3801 17561 3835 17595
rect 8677 17561 8711 17595
rect 12173 17493 12207 17527
rect 12449 17493 12483 17527
rect 12817 17493 12851 17527
rect 14105 17493 14139 17527
rect 1685 17289 1719 17323
rect 2053 17289 2087 17323
rect 3433 17289 3467 17323
rect 5181 17289 5215 17323
rect 7757 17289 7791 17323
rect 10149 17289 10183 17323
rect 13369 17289 13403 17323
rect 13645 17289 13679 17323
rect 16405 17289 16439 17323
rect 17785 17289 17819 17323
rect 20821 17289 20855 17323
rect 22017 17289 22051 17323
rect 23121 17289 23155 17323
rect 8125 17221 8159 17255
rect 9505 17221 9539 17255
rect 14335 17221 14369 17255
rect 20177 17221 20211 17255
rect 23397 17221 23431 17255
rect 2421 17153 2455 17187
rect 3065 17153 3099 17187
rect 6101 17153 6135 17187
rect 6561 17153 6595 17187
rect 10885 17153 10919 17187
rect 16681 17153 16715 17187
rect 19257 17153 19291 17187
rect 20453 17153 20487 17187
rect 21097 17153 21131 17187
rect 21373 17153 21407 17187
rect 24041 17153 24075 17187
rect 3801 17085 3835 17119
rect 4261 17085 4295 17119
rect 6837 17085 6871 17119
rect 8585 17085 8619 17119
rect 12449 17085 12483 17119
rect 15485 17085 15519 17119
rect 18096 17085 18130 17119
rect 18521 17085 18555 17119
rect 22636 17085 22670 17119
rect 2513 17017 2547 17051
rect 4512 17017 4546 17051
rect 5825 17017 5859 17051
rect 7158 17017 7192 17051
rect 8401 17017 8435 17051
rect 8906 17017 8940 17051
rect 10701 17017 10735 17051
rect 10977 17017 11011 17051
rect 11529 17017 11563 17051
rect 11897 17017 11931 17051
rect 12265 17017 12299 17051
rect 12811 17017 12845 17051
rect 15025 17017 15059 17051
rect 15393 17017 15427 17051
rect 15847 17017 15881 17051
rect 17417 17017 17451 17051
rect 19578 17017 19612 17051
rect 21189 17017 21223 17051
rect 22385 17017 22419 17051
rect 23765 17017 23799 17051
rect 23857 17017 23891 17051
rect 4169 16949 4203 16983
rect 9873 16949 9907 16983
rect 14013 16949 14047 16983
rect 18199 16949 18233 16983
rect 19073 16949 19107 16983
rect 22707 16949 22741 16983
rect 24685 16949 24719 16983
rect 3157 16745 3191 16779
rect 3525 16745 3559 16779
rect 4537 16745 4571 16779
rect 7849 16745 7883 16779
rect 8309 16745 8343 16779
rect 9137 16745 9171 16779
rect 11253 16745 11287 16779
rect 13001 16745 13035 16779
rect 15393 16745 15427 16779
rect 16313 16745 16347 16779
rect 16773 16745 16807 16779
rect 19947 16745 19981 16779
rect 22385 16745 22419 16779
rect 24179 16745 24213 16779
rect 2237 16677 2271 16711
rect 2789 16677 2823 16711
rect 6745 16677 6779 16711
rect 7021 16677 7055 16711
rect 10977 16677 11011 16711
rect 12167 16677 12201 16711
rect 14381 16677 14415 16711
rect 19717 16677 19751 16711
rect 21005 16677 21039 16711
rect 21097 16677 21131 16711
rect 22661 16677 22695 16711
rect 23213 16677 23247 16711
rect 4629 16609 4663 16643
rect 4997 16609 5031 16643
rect 6193 16609 6227 16643
rect 6561 16609 6595 16643
rect 8033 16609 8067 16643
rect 8585 16609 8619 16643
rect 10241 16609 10275 16643
rect 10793 16609 10827 16643
rect 13921 16609 13955 16643
rect 14197 16609 14231 16643
rect 15485 16609 15519 16643
rect 15853 16609 15887 16643
rect 18153 16609 18187 16643
rect 18613 16609 18647 16643
rect 19809 16609 19843 16643
rect 23949 16609 23983 16643
rect 25104 16609 25138 16643
rect 2145 16541 2179 16575
rect 11805 16541 11839 16575
rect 16865 16541 16899 16575
rect 18889 16541 18923 16575
rect 21281 16541 21315 16575
rect 22569 16541 22603 16575
rect 23765 16541 23799 16575
rect 25191 16541 25225 16575
rect 20729 16473 20763 16507
rect 1869 16405 1903 16439
rect 4353 16405 4387 16439
rect 12725 16405 12759 16439
rect 13369 16405 13403 16439
rect 17969 16405 18003 16439
rect 19257 16405 19291 16439
rect 1869 16201 1903 16235
rect 2973 16201 3007 16235
rect 6101 16201 6135 16235
rect 8033 16201 8067 16235
rect 11897 16201 11931 16235
rect 14105 16201 14139 16235
rect 20177 16201 20211 16235
rect 21741 16201 21775 16235
rect 23121 16201 23155 16235
rect 24501 16201 24535 16235
rect 2605 16133 2639 16167
rect 18245 16133 18279 16167
rect 21373 16133 21407 16167
rect 22753 16133 22787 16167
rect 2053 16065 2087 16099
rect 3893 16065 3927 16099
rect 4997 16065 5031 16099
rect 10241 16065 10275 16099
rect 11345 16065 11379 16099
rect 12725 16065 12759 16099
rect 16497 16065 16531 16099
rect 19809 16065 19843 16099
rect 20821 16065 20855 16099
rect 22109 16065 22143 16099
rect 24225 16065 24259 16099
rect 25237 16065 25271 16099
rect 5273 15997 5307 16031
rect 5641 15997 5675 16031
rect 6837 15997 6871 16031
rect 7389 15997 7423 16031
rect 9045 15997 9079 16031
rect 9321 15997 9355 16031
rect 10701 15997 10735 16031
rect 11069 15997 11103 16031
rect 11253 15997 11287 16031
rect 15117 15997 15151 16031
rect 15301 15997 15335 16031
rect 23740 15997 23774 16031
rect 24752 15997 24786 16031
rect 2145 15929 2179 15963
rect 3617 15929 3651 15963
rect 3709 15929 3743 15963
rect 12817 15929 12851 15963
rect 13369 15929 13403 15963
rect 15577 15929 15611 15963
rect 16313 15929 16347 15963
rect 16589 15929 16623 15963
rect 17141 15929 17175 15963
rect 18613 15929 18647 15963
rect 18705 15929 18739 15963
rect 19257 15929 19291 15963
rect 20913 15929 20947 15963
rect 3433 15861 3467 15895
rect 4629 15861 4663 15895
rect 5181 15861 5215 15895
rect 6561 15861 6595 15895
rect 6929 15861 6963 15895
rect 8585 15861 8619 15895
rect 8861 15861 8895 15895
rect 9965 15861 9999 15895
rect 12265 15861 12299 15895
rect 13737 15861 13771 15895
rect 14657 15861 14691 15895
rect 15945 15861 15979 15895
rect 17785 15861 17819 15895
rect 20545 15861 20579 15895
rect 22293 15861 22327 15895
rect 23811 15861 23845 15895
rect 24823 15861 24857 15895
rect 25605 15861 25639 15895
rect 1869 15657 1903 15691
rect 3065 15657 3099 15691
rect 8309 15657 8343 15691
rect 9505 15657 9539 15691
rect 14933 15657 14967 15691
rect 15577 15657 15611 15691
rect 16129 15657 16163 15691
rect 18245 15657 18279 15691
rect 18797 15657 18831 15691
rect 19073 15657 19107 15691
rect 19441 15657 19475 15691
rect 19947 15657 19981 15691
rect 23949 15657 23983 15691
rect 24731 15657 24765 15691
rect 2145 15589 2179 15623
rect 2697 15589 2731 15623
rect 4261 15589 4295 15623
rect 5089 15589 5123 15623
rect 5825 15589 5859 15623
rect 6745 15589 6779 15623
rect 7113 15589 7147 15623
rect 7297 15589 7331 15623
rect 7389 15589 7423 15623
rect 2053 15453 2087 15487
rect 4169 15453 4203 15487
rect 5457 15453 5491 15487
rect 5733 15453 5767 15487
rect 6009 15453 6043 15487
rect 7941 15453 7975 15487
rect 4721 15385 4755 15419
rect 9873 15589 9907 15623
rect 13093 15589 13127 15623
rect 13645 15589 13679 15623
rect 21097 15589 21131 15623
rect 23121 15589 23155 15623
rect 23673 15589 23707 15623
rect 11253 15521 11287 15555
rect 11713 15521 11747 15555
rect 19876 15521 19910 15555
rect 24660 15521 24694 15555
rect 9781 15453 9815 15487
rect 11805 15453 11839 15487
rect 12265 15453 12299 15487
rect 13001 15453 13035 15487
rect 15761 15453 15795 15487
rect 17877 15453 17911 15487
rect 20729 15453 20763 15487
rect 21005 15453 21039 15487
rect 22845 15453 22879 15487
rect 23029 15453 23063 15487
rect 10333 15385 10367 15419
rect 21557 15385 21591 15419
rect 3893 15317 3927 15351
rect 8769 15317 8803 15351
rect 9505 15317 9539 15351
rect 10885 15317 10919 15351
rect 12725 15317 12759 15351
rect 16681 15317 16715 15351
rect 4077 15113 4111 15147
rect 7757 15113 7791 15147
rect 8033 15113 8067 15147
rect 9873 15113 9907 15147
rect 10149 15113 10183 15147
rect 12173 15113 12207 15147
rect 12449 15113 12483 15147
rect 13461 15113 13495 15147
rect 13829 15113 13863 15147
rect 17233 15113 17267 15147
rect 20269 15113 20303 15147
rect 22661 15113 22695 15147
rect 23029 15113 23063 15147
rect 5641 15045 5675 15079
rect 11345 15045 11379 15079
rect 2697 14977 2731 15011
rect 3341 14977 3375 15011
rect 8953 14977 8987 15011
rect 10793 14977 10827 15011
rect 11805 14977 11839 15011
rect 1460 14909 1494 14943
rect 1869 14909 1903 14943
rect 4169 14909 4203 14943
rect 5089 14909 5123 14943
rect 6285 14909 6319 14943
rect 6837 14909 6871 14943
rect 21189 15045 21223 15079
rect 15669 14977 15703 15011
rect 16865 14977 16899 15011
rect 17877 14977 17911 15011
rect 19349 14977 19383 15011
rect 20545 14977 20579 15011
rect 21741 14977 21775 15011
rect 23765 14977 23799 15011
rect 24041 14977 24075 15011
rect 24777 14977 24811 15011
rect 12541 14909 12575 14943
rect 14289 14909 14323 14943
rect 14749 14909 14783 14943
rect 18388 14909 18422 14943
rect 19257 14909 19291 14943
rect 23397 14909 23431 14943
rect 25288 14909 25322 14943
rect 1547 14841 1581 14875
rect 2789 14841 2823 14875
rect 3709 14841 3743 14875
rect 6653 14841 6687 14875
rect 7199 14841 7233 14875
rect 8861 14841 8895 14875
rect 9315 14841 9349 14875
rect 10885 14841 10919 14875
rect 12449 14841 12483 14875
rect 12862 14841 12896 14875
rect 15209 14841 15243 14875
rect 15577 14841 15611 14875
rect 16031 14841 16065 14875
rect 18475 14841 18509 14875
rect 19711 14841 19745 14875
rect 23857 14841 23891 14875
rect 25375 14841 25409 14875
rect 2329 14773 2363 14807
rect 4537 14773 4571 14807
rect 10517 14773 10551 14807
rect 14473 14773 14507 14807
rect 16589 14773 16623 14807
rect 18889 14773 18923 14807
rect 21649 14773 21683 14807
rect 22109 14773 22143 14807
rect 25789 14773 25823 14807
rect 2973 14569 3007 14603
rect 3525 14569 3559 14603
rect 4537 14569 4571 14603
rect 6469 14569 6503 14603
rect 7665 14569 7699 14603
rect 8953 14569 8987 14603
rect 10609 14569 10643 14603
rect 10885 14569 10919 14603
rect 13093 14569 13127 14603
rect 13645 14569 13679 14603
rect 18981 14569 19015 14603
rect 19993 14569 20027 14603
rect 20637 14569 20671 14603
rect 2053 14501 2087 14535
rect 2605 14501 2639 14535
rect 7941 14501 7975 14535
rect 8033 14501 8067 14535
rect 10051 14501 10085 14535
rect 12173 14501 12207 14535
rect 15939 14501 15973 14535
rect 17509 14501 17543 14535
rect 21005 14501 21039 14535
rect 21097 14501 21131 14535
rect 23305 14501 23339 14535
rect 23857 14501 23891 14535
rect 24869 14501 24903 14535
rect 4169 14433 4203 14467
rect 7021 14433 7055 14467
rect 13829 14433 13863 14467
rect 14013 14433 14047 14467
rect 15577 14433 15611 14467
rect 18889 14433 18923 14467
rect 19349 14433 19383 14467
rect 1777 14365 1811 14399
rect 1961 14365 1995 14399
rect 6101 14365 6135 14399
rect 8217 14365 8251 14399
rect 9413 14365 9447 14399
rect 9689 14365 9723 14399
rect 12081 14365 12115 14399
rect 12725 14365 12759 14399
rect 17417 14365 17451 14399
rect 17693 14365 17727 14399
rect 21373 14365 21407 14399
rect 23029 14365 23063 14399
rect 23213 14365 23247 14399
rect 24777 14365 24811 14399
rect 25053 14365 25087 14399
rect 3893 14297 3927 14331
rect 5089 14297 5123 14331
rect 5641 14229 5675 14263
rect 7297 14229 7331 14263
rect 11253 14229 11287 14263
rect 16497 14229 16531 14263
rect 18337 14229 18371 14263
rect 22661 14229 22695 14263
rect 24225 14229 24259 14263
rect 1777 14025 1811 14059
rect 7849 14025 7883 14059
rect 8585 14025 8619 14059
rect 9873 14025 9907 14059
rect 11897 14025 11931 14059
rect 12173 14025 12207 14059
rect 15853 14025 15887 14059
rect 17693 14025 17727 14059
rect 18889 14025 18923 14059
rect 20085 14025 20119 14059
rect 21833 14025 21867 14059
rect 22707 14025 22741 14059
rect 24777 14025 24811 14059
rect 25375 14025 25409 14059
rect 2881 13957 2915 13991
rect 13553 13957 13587 13991
rect 18245 13957 18279 13991
rect 2605 13889 2639 13923
rect 3801 13889 3835 13923
rect 5917 13889 5951 13923
rect 9505 13889 9539 13923
rect 10149 13889 10183 13923
rect 12817 13889 12851 13923
rect 15485 13889 15519 13923
rect 17049 13889 17083 13923
rect 19257 13889 19291 13923
rect 5089 13821 5123 13855
rect 5365 13821 5399 13855
rect 5641 13821 5675 13855
rect 6837 13821 6871 13855
rect 7297 13821 7331 13855
rect 8217 13821 8251 13855
rect 8769 13821 8803 13855
rect 9229 13821 9263 13855
rect 9597 13821 9631 13855
rect 10701 13821 10735 13855
rect 10977 13821 11011 13855
rect 11253 13821 11287 13855
rect 14013 13821 14047 13855
rect 14749 13821 14783 13855
rect 15209 13821 15243 13855
rect 18061 13821 18095 13855
rect 18521 13821 18555 13855
rect 19901 13821 19935 13855
rect 1961 13753 1995 13787
rect 2053 13753 2087 13787
rect 3525 13753 3559 13787
rect 3617 13753 3651 13787
rect 11529 13753 11563 13787
rect 12541 13753 12575 13787
rect 12633 13753 12667 13787
rect 14565 13753 14599 13787
rect 16405 13753 16439 13787
rect 16497 13753 16531 13787
rect 19349 13753 19383 13787
rect 20637 13957 20671 13991
rect 21373 13957 21407 13991
rect 22109 13957 22143 13991
rect 23029 13957 23063 13991
rect 20821 13889 20855 13923
rect 23765 13889 23799 13923
rect 24041 13889 24075 13923
rect 25053 13889 25087 13923
rect 22569 13821 22603 13855
rect 25288 13821 25322 13855
rect 20177 13753 20211 13787
rect 20913 13753 20947 13787
rect 23397 13753 23431 13787
rect 23857 13753 23891 13787
rect 25789 13753 25823 13787
rect 3341 13685 3375 13719
rect 4537 13685 4571 13719
rect 6193 13685 6227 13719
rect 6561 13685 6595 13719
rect 6929 13685 6963 13719
rect 9597 13685 9631 13719
rect 16221 13685 16255 13719
rect 17417 13685 17451 13719
rect 20085 13685 20119 13719
rect 1961 13481 1995 13515
rect 3525 13481 3559 13515
rect 3893 13481 3927 13515
rect 5181 13481 5215 13515
rect 6101 13481 6135 13515
rect 7941 13481 7975 13515
rect 9781 13481 9815 13515
rect 12173 13481 12207 13515
rect 14749 13481 14783 13515
rect 16313 13481 16347 13515
rect 16681 13481 16715 13515
rect 18981 13481 19015 13515
rect 20637 13481 20671 13515
rect 23765 13481 23799 13515
rect 2421 13413 2455 13447
rect 4261 13413 4295 13447
rect 6653 13413 6687 13447
rect 8217 13413 8251 13447
rect 11615 13413 11649 13447
rect 14381 13413 14415 13447
rect 19441 13413 19475 13447
rect 19993 13413 20027 13447
rect 21005 13413 21039 13447
rect 21097 13413 21131 13447
rect 22753 13413 22787 13447
rect 24317 13413 24351 13447
rect 9873 13345 9907 13379
rect 10149 13345 10183 13379
rect 12449 13345 12483 13379
rect 13645 13345 13679 13379
rect 14105 13345 14139 13379
rect 15945 13345 15979 13379
rect 17877 13345 17911 13379
rect 18153 13345 18187 13379
rect 2329 13277 2363 13311
rect 2973 13277 3007 13311
rect 4169 13277 4203 13311
rect 4537 13277 4571 13311
rect 6561 13277 6595 13311
rect 8125 13277 8159 13311
rect 8401 13277 8435 13311
rect 11253 13277 11287 13311
rect 18429 13277 18463 13311
rect 19349 13277 19383 13311
rect 21281 13277 21315 13311
rect 21925 13277 21959 13311
rect 22661 13277 22695 13311
rect 24225 13277 24259 13311
rect 24501 13277 24535 13311
rect 7113 13209 7147 13243
rect 12817 13209 12851 13243
rect 23213 13209 23247 13243
rect 7481 13141 7515 13175
rect 10885 13141 10919 13175
rect 15577 13141 15611 13175
rect 4721 12937 4755 12971
rect 5917 12937 5951 12971
rect 10149 12937 10183 12971
rect 11897 12937 11931 12971
rect 13737 12937 13771 12971
rect 14013 12937 14047 12971
rect 17785 12937 17819 12971
rect 19625 12937 19659 12971
rect 20085 12937 20119 12971
rect 21373 12937 21407 12971
rect 23489 12937 23523 12971
rect 24685 12937 24719 12971
rect 1777 12869 1811 12903
rect 2881 12869 2915 12903
rect 9873 12869 9907 12903
rect 10701 12869 10735 12903
rect 16405 12869 16439 12903
rect 19349 12869 19383 12903
rect 1961 12801 1995 12835
rect 3801 12801 3835 12835
rect 5089 12801 5123 12835
rect 12817 12801 12851 12835
rect 14565 12801 14599 12835
rect 15853 12801 15887 12835
rect 22017 12801 22051 12835
rect 22661 12801 22695 12835
rect 24041 12801 24075 12835
rect 25237 12801 25271 12835
rect 5733 12733 5767 12767
rect 6193 12733 6227 12767
rect 7573 12733 7607 12767
rect 8585 12733 8619 12767
rect 10977 12733 11011 12767
rect 11253 12733 11287 12767
rect 18245 12733 18279 12767
rect 18705 12733 18739 12767
rect 20177 12733 20211 12767
rect 21097 12733 21131 12767
rect 21741 12733 21775 12767
rect 2053 12665 2087 12699
rect 2605 12665 2639 12699
rect 3617 12665 3651 12699
rect 3886 12665 3920 12699
rect 4445 12665 4479 12699
rect 6929 12665 6963 12699
rect 7021 12665 7055 12699
rect 8493 12665 8527 12699
rect 8947 12665 8981 12699
rect 11529 12665 11563 12699
rect 12541 12665 12575 12699
rect 12633 12665 12667 12699
rect 14289 12665 14323 12699
rect 14381 12665 14415 12699
rect 15945 12665 15979 12699
rect 18981 12665 19015 12699
rect 20498 12665 20532 12699
rect 22109 12665 22143 12699
rect 23765 12665 23799 12699
rect 23857 12665 23891 12699
rect 5549 12597 5583 12631
rect 6653 12597 6687 12631
rect 8033 12597 8067 12631
rect 9505 12597 9539 12631
rect 12265 12597 12299 12631
rect 15209 12597 15243 12631
rect 15577 12597 15611 12631
rect 17141 12597 17175 12631
rect 17509 12597 17543 12631
rect 22937 12597 22971 12631
rect 1685 12393 1719 12427
rect 2053 12393 2087 12427
rect 3801 12393 3835 12427
rect 5089 12393 5123 12427
rect 6929 12393 6963 12427
rect 7205 12393 7239 12427
rect 7941 12393 7975 12427
rect 11437 12393 11471 12427
rect 11989 12393 12023 12427
rect 12541 12393 12575 12427
rect 15025 12393 15059 12427
rect 16313 12393 16347 12427
rect 19625 12393 19659 12427
rect 20729 12393 20763 12427
rect 21557 12393 21591 12427
rect 22109 12393 22143 12427
rect 23765 12393 23799 12427
rect 2329 12325 2363 12359
rect 4490 12325 4524 12359
rect 6330 12325 6364 12359
rect 8217 12325 8251 12359
rect 13829 12325 13863 12359
rect 14381 12325 14415 12359
rect 15485 12325 15519 12359
rect 16037 12325 16071 12359
rect 19026 12325 19060 12359
rect 24317 12325 24351 12359
rect 24869 12325 24903 12359
rect 10149 12257 10183 12291
rect 16957 12257 16991 12291
rect 18705 12257 18739 12291
rect 21189 12257 21223 12291
rect 2237 12189 2271 12223
rect 2605 12189 2639 12223
rect 4169 12189 4203 12223
rect 6009 12189 6043 12223
rect 8125 12189 8159 12223
rect 11621 12189 11655 12223
rect 13737 12189 13771 12223
rect 15393 12189 15427 12223
rect 16865 12189 16899 12223
rect 22937 12189 22971 12223
rect 24225 12189 24259 12223
rect 8677 12121 8711 12155
rect 18337 12121 18371 12155
rect 9045 12053 9079 12087
rect 10517 12053 10551 12087
rect 11069 12053 11103 12087
rect 12909 12053 12943 12087
rect 13553 12053 13587 12087
rect 14749 12053 14783 12087
rect 20269 12053 20303 12087
rect 22661 12053 22695 12087
rect 3341 11849 3375 11883
rect 5181 11849 5215 11883
rect 5457 11849 5491 11883
rect 7251 11849 7285 11883
rect 9413 11849 9447 11883
rect 9689 11849 9723 11883
rect 10609 11849 10643 11883
rect 11897 11849 11931 11883
rect 12817 11849 12851 11883
rect 14565 11849 14599 11883
rect 14933 11849 14967 11883
rect 17877 11849 17911 11883
rect 19809 11849 19843 11883
rect 21281 11849 21315 11883
rect 21649 11849 21683 11883
rect 22753 11849 22787 11883
rect 25053 11849 25087 11883
rect 2605 11781 2639 11815
rect 9045 11781 9079 11815
rect 16865 11781 16899 11815
rect 17141 11781 17175 11815
rect 8125 11713 8159 11747
rect 11161 11713 11195 11747
rect 13185 11713 13219 11747
rect 15485 11713 15519 11747
rect 15761 11713 15795 11747
rect 16497 11713 16531 11747
rect 18429 11713 18463 11747
rect 18889 11713 18923 11747
rect 23489 11713 23523 11747
rect 24133 11713 24167 11747
rect 24777 11713 24811 11747
rect 3801 11645 3835 11679
rect 4261 11645 4295 11679
rect 7148 11645 7182 11679
rect 7573 11645 7607 11679
rect 12265 11645 12299 11679
rect 12633 11645 12667 11679
rect 13645 11645 13679 11679
rect 16957 11645 16991 11679
rect 20637 11645 20671 11679
rect 21833 11645 21867 11679
rect 23857 11645 23891 11679
rect 25640 11645 25674 11679
rect 26065 11645 26099 11679
rect 2053 11577 2087 11611
rect 2145 11577 2179 11611
rect 4169 11577 4203 11611
rect 4623 11577 4657 11611
rect 6101 11577 6135 11611
rect 8033 11577 8067 11611
rect 8487 11577 8521 11611
rect 10885 11577 10919 11611
rect 10977 11577 11011 11611
rect 13461 11577 13495 11611
rect 13966 11577 14000 11611
rect 15577 11577 15611 11611
rect 19210 11577 19244 11611
rect 22154 11577 22188 11611
rect 24225 11577 24259 11611
rect 1777 11509 1811 11543
rect 3065 11509 3099 11543
rect 6469 11509 6503 11543
rect 10241 11509 10275 11543
rect 15301 11509 15335 11543
rect 17509 11509 17543 11543
rect 18797 11509 18831 11543
rect 20453 11509 20487 11543
rect 20821 11509 20855 11543
rect 25743 11509 25777 11543
rect 4537 11305 4571 11339
rect 7021 11305 7055 11339
rect 7941 11305 7975 11339
rect 10149 11305 10183 11339
rect 11621 11305 11655 11339
rect 12495 11305 12529 11339
rect 14933 11305 14967 11339
rect 19993 11305 20027 11339
rect 21005 11305 21039 11339
rect 24731 11305 24765 11339
rect 2237 11237 2271 11271
rect 2789 11237 2823 11271
rect 4353 11237 4387 11271
rect 6422 11237 6456 11271
rect 8769 11237 8803 11271
rect 10517 11237 10551 11271
rect 11069 11237 11103 11271
rect 13731 11237 13765 11271
rect 15485 11237 15519 11271
rect 19394 11237 19428 11271
rect 21925 11237 21959 11271
rect 23213 11237 23247 11271
rect 24133 11237 24167 11271
rect 4445 11169 4479 11203
rect 4997 11169 5031 11203
rect 8309 11169 8343 11203
rect 8585 11169 8619 11203
rect 12392 11169 12426 11203
rect 14289 11169 14323 11203
rect 17785 11169 17819 11203
rect 17969 11169 18003 11203
rect 18245 11169 18279 11203
rect 21005 11169 21039 11203
rect 21373 11169 21407 11203
rect 24660 11169 24694 11203
rect 2145 11101 2179 11135
rect 6101 11101 6135 11135
rect 10425 11101 10459 11135
rect 13369 11101 13403 11135
rect 14565 11101 14599 11135
rect 15393 11101 15427 11135
rect 15761 11101 15795 11135
rect 16681 11101 16715 11135
rect 19073 11101 19107 11135
rect 20637 11101 20671 11135
rect 23121 11101 23155 11135
rect 23673 11033 23707 11067
rect 1869 10965 1903 10999
rect 9413 10965 9447 10999
rect 12909 10965 12943 10999
rect 16405 10965 16439 10999
rect 18889 10965 18923 10999
rect 1777 10761 1811 10795
rect 2053 10761 2087 10795
rect 4261 10761 4295 10795
rect 5457 10761 5491 10795
rect 6193 10761 6227 10795
rect 7941 10761 7975 10795
rect 9873 10761 9907 10795
rect 11253 10761 11287 10795
rect 12633 10761 12667 10795
rect 13737 10761 13771 10795
rect 17141 10761 17175 10795
rect 17601 10761 17635 10795
rect 22753 10761 22787 10795
rect 23489 10761 23523 10795
rect 25421 10761 25455 10795
rect 7205 10693 7239 10727
rect 15025 10693 15059 10727
rect 15209 10693 15243 10727
rect 16221 10693 16255 10727
rect 20085 10693 20119 10727
rect 2973 10625 3007 10659
rect 5181 10625 5215 10659
rect 7573 10625 7607 10659
rect 13461 10625 13495 10659
rect 21281 10625 21315 10659
rect 23121 10625 23155 10659
rect 24041 10625 24075 10659
rect 4721 10557 4755 10591
rect 4997 10557 5031 10591
rect 7021 10557 7055 10591
rect 8677 10557 8711 10591
rect 9045 10557 9079 10591
rect 9505 10557 9539 10591
rect 10333 10557 10367 10591
rect 13093 10557 13127 10591
rect 14841 10557 14875 10591
rect 15117 10557 15151 10591
rect 15393 10557 15427 10591
rect 16957 10557 16991 10591
rect 18981 10557 19015 10591
rect 19441 10557 19475 10591
rect 25237 10557 25271 10591
rect 2329 10489 2363 10523
rect 2421 10489 2455 10523
rect 3617 10489 3651 10523
rect 3893 10489 3927 10523
rect 6653 10489 6687 10523
rect 10241 10489 10275 10523
rect 10695 10489 10729 10523
rect 12173 10489 12207 10523
rect 12909 10489 12943 10523
rect 14289 10489 14323 10523
rect 18521 10489 18555 10523
rect 19717 10489 19751 10523
rect 21373 10489 21407 10523
rect 21925 10489 21959 10523
rect 23765 10489 23799 10523
rect 23857 10489 23891 10523
rect 25697 10489 25731 10523
rect 8309 10421 8343 10455
rect 11529 10421 11563 10455
rect 14565 10421 14599 10455
rect 14841 10421 14875 10455
rect 15577 10421 15611 10455
rect 16865 10421 16899 10455
rect 18797 10421 18831 10455
rect 20545 10421 20579 10455
rect 21005 10421 21039 10455
rect 22201 10421 22235 10455
rect 24777 10421 24811 10455
rect 1547 10217 1581 10251
rect 2559 10217 2593 10251
rect 4445 10217 4479 10251
rect 6193 10217 6227 10251
rect 6929 10217 6963 10251
rect 10793 10217 10827 10251
rect 13921 10217 13955 10251
rect 22109 10217 22143 10251
rect 22753 10217 22787 10251
rect 23765 10217 23799 10251
rect 24363 10217 24397 10251
rect 25375 10217 25409 10251
rect 8217 10149 8251 10183
rect 10609 10149 10643 10183
rect 17278 10149 17312 10183
rect 21189 10149 21223 10183
rect 1444 10081 1478 10115
rect 2488 10081 2522 10115
rect 4629 10081 4663 10115
rect 4905 10081 4939 10115
rect 6193 10081 6227 10115
rect 6469 10081 6503 10115
rect 9740 10081 9774 10115
rect 10701 10081 10735 10115
rect 11161 10081 11195 10115
rect 11621 10081 11655 10115
rect 11897 10081 11931 10115
rect 13001 10081 13035 10115
rect 13461 10081 13495 10115
rect 13783 10081 13817 10115
rect 14933 10081 14967 10115
rect 15209 10081 15243 10115
rect 15393 10081 15427 10115
rect 15577 10081 15611 10115
rect 19257 10081 19291 10115
rect 19717 10081 19751 10115
rect 22937 10081 22971 10115
rect 23121 10081 23155 10115
rect 24260 10081 24294 10115
rect 25237 10081 25271 10115
rect 8125 10013 8159 10047
rect 9827 10013 9861 10047
rect 10241 10013 10275 10047
rect 14749 10013 14783 10047
rect 8677 9945 8711 9979
rect 16037 10013 16071 10047
rect 16957 10013 16991 10047
rect 19993 10013 20027 10047
rect 20913 10013 20947 10047
rect 18153 9945 18187 9979
rect 2237 9877 2271 9911
rect 2881 9877 2915 9911
rect 9137 9877 9171 9911
rect 9505 9877 9539 9911
rect 12725 9877 12759 9911
rect 14933 9877 14967 9911
rect 15025 9877 15059 9911
rect 16313 9877 16347 9911
rect 17877 9877 17911 9911
rect 18981 9877 19015 9911
rect 20729 9877 20763 9911
rect 21833 9877 21867 9911
rect 1869 9673 1903 9707
rect 3341 9673 3375 9707
rect 3985 9673 4019 9707
rect 4353 9673 4387 9707
rect 5871 9673 5905 9707
rect 6561 9673 6595 9707
rect 7757 9673 7791 9707
rect 9137 9673 9171 9707
rect 9781 9673 9815 9707
rect 13829 9673 13863 9707
rect 15393 9673 15427 9707
rect 17509 9673 17543 9707
rect 19625 9673 19659 9707
rect 21097 9673 21131 9707
rect 23305 9673 23339 9707
rect 24133 9673 24167 9707
rect 24593 9673 24627 9707
rect 24869 9673 24903 9707
rect 1547 9605 1581 9639
rect 4583 9605 4617 9639
rect 6285 9605 6319 9639
rect 25329 9605 25363 9639
rect 2237 9537 2271 9571
rect 3433 9537 3467 9571
rect 7205 9537 7239 9571
rect 11529 9537 11563 9571
rect 14197 9537 14231 9571
rect 16589 9537 16623 9571
rect 18613 9537 18647 9571
rect 19901 9537 19935 9571
rect 19993 9537 20027 9571
rect 20177 9537 20211 9571
rect 22017 9537 22051 9571
rect 22293 9537 22327 9571
rect 1476 9469 1510 9503
rect 2456 9469 2490 9503
rect 2881 9469 2915 9503
rect 4512 9469 4546 9503
rect 5800 9469 5834 9503
rect 8217 9469 8251 9503
rect 10793 9469 10827 9503
rect 10885 9469 10919 9503
rect 11069 9469 11103 9503
rect 12725 9469 12759 9503
rect 13553 9469 13587 9503
rect 13737 9469 13771 9503
rect 14841 9469 14875 9503
rect 15853 9469 15887 9503
rect 16313 9469 16347 9503
rect 2559 9401 2593 9435
rect 5641 9401 5675 9435
rect 8125 9401 8159 9435
rect 8579 9401 8613 9435
rect 17785 9401 17819 9435
rect 18153 9401 18187 9435
rect 18245 9401 18279 9435
rect 19901 9401 19935 9435
rect 20498 9401 20532 9435
rect 21741 9401 21775 9435
rect 22109 9401 22143 9435
rect 4997 9333 5031 9367
rect 10333 9333 10367 9367
rect 10701 9333 10735 9367
rect 11897 9333 11931 9367
rect 12265 9333 12299 9367
rect 14473 9333 14507 9367
rect 15025 9333 15059 9367
rect 15761 9333 15795 9367
rect 16957 9333 16991 9367
rect 19257 9333 19291 9367
rect 21373 9333 21407 9367
rect 22937 9333 22971 9367
rect 23673 9333 23707 9367
rect 2421 9129 2455 9163
rect 7941 9129 7975 9163
rect 10793 9129 10827 9163
rect 14473 9129 14507 9163
rect 15577 9129 15611 9163
rect 16957 9129 16991 9163
rect 20177 9129 20211 9163
rect 21833 9129 21867 9163
rect 22109 9129 22143 9163
rect 23811 9129 23845 9163
rect 6561 9061 6595 9095
rect 8217 9061 8251 9095
rect 8769 9061 8803 9095
rect 9137 9061 9171 9095
rect 13829 9061 13863 9095
rect 19625 9061 19659 9095
rect 21234 9061 21268 9095
rect 22799 9061 22833 9095
rect 1444 8993 1478 9027
rect 6009 8993 6043 9027
rect 6285 8993 6319 9027
rect 9505 8993 9539 9027
rect 9689 8993 9723 9027
rect 10701 8993 10735 9027
rect 11437 8993 11471 9027
rect 11621 8993 11655 9027
rect 12081 8993 12115 9027
rect 13001 8993 13035 9027
rect 13185 8993 13219 9027
rect 15669 8993 15703 9027
rect 17325 8993 17359 9027
rect 17785 8993 17819 9027
rect 19165 8993 19199 9027
rect 19349 8993 19383 9027
rect 20913 8993 20947 9027
rect 22661 8993 22695 9027
rect 23740 8993 23774 9027
rect 8125 8925 8159 8959
rect 18061 8925 18095 8959
rect 18337 8925 18371 8959
rect 1547 8857 1581 8891
rect 12817 8857 12851 8891
rect 9873 8789 9907 8823
rect 10333 8789 10367 8823
rect 13277 8789 13311 8823
rect 14749 8789 14783 8823
rect 16313 8789 16347 8823
rect 1593 8585 1627 8619
rect 2007 8585 2041 8619
rect 3019 8585 3053 8619
rect 5917 8585 5951 8619
rect 6285 8585 6319 8619
rect 6975 8585 7009 8619
rect 7849 8585 7883 8619
rect 8953 8585 8987 8619
rect 9321 8585 9355 8619
rect 10701 8585 10735 8619
rect 11713 8585 11747 8619
rect 12725 8585 12759 8619
rect 14013 8585 14047 8619
rect 17325 8585 17359 8619
rect 19625 8585 19659 8619
rect 19993 8585 20027 8619
rect 20729 8585 20763 8619
rect 21005 8585 21039 8619
rect 22201 8585 22235 8619
rect 23857 8585 23891 8619
rect 10517 8517 10551 8551
rect 14841 8517 14875 8551
rect 19257 8517 19291 8551
rect 7389 8449 7423 8483
rect 8585 8449 8619 8483
rect 9045 8449 9079 8483
rect 9965 8449 9999 8483
rect 10609 8449 10643 8483
rect 11253 8449 11287 8483
rect 13645 8449 13679 8483
rect 16405 8449 16439 8483
rect 17785 8449 17819 8483
rect 18061 8449 18095 8483
rect 21925 8449 21959 8483
rect 1904 8381 1938 8415
rect 2329 8381 2363 8415
rect 2916 8381 2950 8415
rect 3341 8381 3375 8415
rect 6904 8381 6938 8415
rect 8217 8381 8251 8415
rect 8824 8381 8858 8415
rect 8677 8313 8711 8347
rect 10388 8381 10422 8415
rect 12633 8381 12667 8415
rect 14749 8381 14783 8415
rect 15025 8381 15059 8415
rect 16313 8381 16347 8415
rect 16589 8381 16623 8415
rect 20244 8381 20278 8415
rect 10241 8313 10275 8347
rect 12449 8313 12483 8347
rect 18382 8313 18416 8347
rect 21281 8313 21315 8347
rect 21373 8313 21407 8347
rect 9689 8245 9723 8279
rect 9965 8245 9999 8279
rect 10057 8245 10091 8279
rect 12173 8245 12207 8279
rect 13369 8245 13403 8279
rect 14565 8245 14599 8279
rect 15209 8245 15243 8279
rect 15761 8245 15795 8279
rect 16129 8245 16163 8279
rect 16773 8245 16807 8279
rect 18981 8245 19015 8279
rect 20315 8245 20349 8279
rect 22661 8245 22695 8279
rect 1547 8041 1581 8075
rect 9045 8041 9079 8075
rect 11805 8041 11839 8075
rect 12449 8041 12483 8075
rect 12725 8041 12759 8075
rect 13093 8041 13127 8075
rect 14841 8041 14875 8075
rect 17049 8041 17083 8075
rect 19763 8041 19797 8075
rect 20637 8041 20671 8075
rect 2559 7973 2593 8007
rect 8033 7973 8067 8007
rect 9781 7973 9815 8007
rect 10793 7973 10827 8007
rect 18245 7973 18279 8007
rect 21234 7973 21268 8007
rect 1476 7905 1510 7939
rect 2421 7905 2455 7939
rect 8585 7905 8619 7939
rect 9928 7905 9962 7939
rect 11345 7905 11379 7939
rect 11621 7905 11655 7939
rect 14289 7905 14323 7939
rect 15301 7905 15335 7939
rect 15577 7905 15611 7939
rect 16865 7905 16899 7939
rect 19692 7905 19726 7939
rect 20085 7905 20119 7939
rect 10149 7837 10183 7871
rect 14381 7837 14415 7871
rect 15393 7837 15427 7871
rect 15761 7837 15795 7871
rect 18153 7837 18187 7871
rect 18613 7837 18647 7871
rect 20913 7837 20947 7871
rect 10241 7769 10275 7803
rect 11437 7769 11471 7803
rect 16313 7769 16347 7803
rect 8769 7701 8803 7735
rect 9505 7701 9539 7735
rect 10057 7701 10091 7735
rect 11253 7701 11287 7735
rect 16681 7701 16715 7735
rect 17325 7701 17359 7735
rect 17877 7701 17911 7735
rect 19073 7701 19107 7735
rect 21833 7701 21867 7735
rect 1547 7497 1581 7531
rect 1869 7497 1903 7531
rect 8677 7497 8711 7531
rect 9413 7497 9447 7531
rect 9689 7497 9723 7531
rect 16129 7497 16163 7531
rect 17417 7497 17451 7531
rect 17877 7497 17911 7531
rect 19073 7497 19107 7531
rect 19441 7497 19475 7531
rect 21005 7497 21039 7531
rect 14197 7429 14231 7463
rect 14841 7429 14875 7463
rect 11621 7361 11655 7395
rect 13001 7361 13035 7395
rect 13185 7361 13219 7395
rect 17141 7361 17175 7395
rect 18153 7361 18187 7395
rect 18797 7361 18831 7395
rect 21925 7361 21959 7395
rect 1476 7293 1510 7327
rect 9531 7293 9565 7327
rect 10057 7293 10091 7327
rect 10425 7293 10459 7327
rect 11161 7293 11195 7327
rect 13093 7293 13127 7327
rect 13369 7293 13403 7327
rect 14749 7293 14783 7327
rect 15025 7293 15059 7327
rect 15761 7293 15795 7327
rect 19625 7293 19659 7327
rect 20085 7293 20119 7327
rect 9045 7225 9079 7259
rect 11253 7225 11287 7259
rect 13829 7225 13863 7259
rect 15485 7225 15519 7259
rect 16497 7225 16531 7259
rect 16589 7225 16623 7259
rect 18245 7225 18279 7259
rect 20361 7225 20395 7259
rect 21465 7225 21499 7259
rect 21557 7225 21591 7259
rect 2513 7157 2547 7191
rect 11989 7157 12023 7191
rect 14565 7157 14599 7191
rect 22385 7157 22419 7191
rect 1593 6953 1627 6987
rect 9413 6953 9447 6987
rect 14841 6953 14875 6987
rect 15485 6953 15519 6987
rect 16129 6953 16163 6987
rect 17693 6953 17727 6987
rect 19855 6953 19889 6987
rect 21465 6953 21499 6987
rect 9689 6885 9723 6919
rect 15761 6885 15795 6919
rect 16767 6885 16801 6919
rect 18337 6885 18371 6919
rect 21741 6885 21775 6919
rect 10333 6817 10367 6851
rect 11345 6817 11379 6851
rect 13277 6817 13311 6851
rect 14105 6817 14139 6851
rect 14289 6817 14323 6851
rect 15301 6817 15335 6851
rect 19752 6817 19786 6851
rect 11989 6749 12023 6783
rect 14381 6749 14415 6783
rect 16405 6749 16439 6783
rect 18245 6749 18279 6783
rect 17325 6681 17359 6715
rect 18797 6681 18831 6715
rect 10885 6613 10919 6647
rect 13185 6613 13219 6647
rect 18061 6613 18095 6647
rect 9689 6409 9723 6443
rect 10333 6409 10367 6443
rect 12633 6409 12667 6443
rect 13461 6409 13495 6443
rect 16497 6409 16531 6443
rect 16865 6409 16899 6443
rect 19717 6409 19751 6443
rect 10885 6341 10919 6375
rect 11805 6341 11839 6375
rect 15485 6341 15519 6375
rect 11253 6273 11287 6307
rect 14565 6273 14599 6307
rect 15025 6273 15059 6307
rect 17877 6273 17911 6307
rect 18061 6273 18095 6307
rect 9321 6205 9355 6239
rect 9597 6205 9631 6239
rect 10793 6205 10827 6239
rect 11069 6205 11103 6239
rect 12173 6205 12207 6239
rect 12449 6205 12483 6239
rect 12909 6205 12943 6239
rect 13645 6205 13679 6239
rect 14473 6205 14507 6239
rect 14749 6205 14783 6239
rect 15577 6205 15611 6239
rect 17509 6205 17543 6239
rect 18153 6205 18187 6239
rect 9413 6137 9447 6171
rect 15898 6137 15932 6171
rect 10701 6069 10735 6103
rect 9413 5865 9447 5899
rect 13001 5865 13035 5899
rect 13461 5865 13495 5899
rect 14381 5865 14415 5899
rect 15485 5865 15519 5899
rect 16221 5865 16255 5899
rect 16589 5865 16623 5899
rect 18245 5865 18279 5899
rect 18337 5865 18371 5899
rect 11897 5797 11931 5831
rect 13185 5797 13219 5831
rect 14013 5797 14047 5831
rect 16957 5797 16991 5831
rect 17509 5797 17543 5831
rect 10885 5729 10919 5763
rect 11069 5729 11103 5763
rect 11437 5729 11471 5763
rect 13369 5729 13403 5763
rect 15761 5729 15795 5763
rect 16865 5661 16899 5695
rect 15945 5525 15979 5559
rect 11805 5321 11839 5355
rect 13277 5321 13311 5355
rect 13553 5321 13587 5355
rect 14013 5321 14047 5355
rect 16129 5321 16163 5355
rect 14473 5253 14507 5287
rect 11161 5185 11195 5219
rect 17049 5185 17083 5219
rect 17325 5185 17359 5219
rect 9873 5117 9907 5151
rect 10241 5117 10275 5151
rect 10517 5117 10551 5151
rect 14289 5117 14323 5151
rect 14749 5117 14783 5151
rect 15301 5117 15335 5151
rect 15761 5117 15795 5151
rect 16681 5117 16715 5151
rect 11529 4981 11563 5015
rect 15485 4981 15519 5015
rect 10977 4777 11011 4811
rect 16635 4777 16669 4811
rect 16957 4777 16991 4811
rect 21971 4777 22005 4811
rect 10885 4641 10919 4675
rect 16564 4641 16598 4675
rect 21741 4641 21775 4675
rect 16405 4573 16439 4607
rect 16589 4233 16623 4267
rect 21925 4233 21959 4267
rect 10793 3893 10827 3927
rect 1444 3553 1478 3587
rect 1547 3485 1581 3519
rect 1593 3145 1627 3179
rect 24731 2601 24765 2635
rect 24660 2465 24694 2499
rect 25145 2261 25179 2295
<< metal1 >>
rect 4798 27480 4804 27532
rect 4856 27520 4862 27532
rect 6454 27520 6460 27532
rect 4856 27492 6460 27520
rect 4856 27480 4862 27492
rect 6454 27480 6460 27492
rect 6512 27480 6518 27532
rect 9674 27480 9680 27532
rect 9732 27520 9738 27532
rect 10410 27520 10416 27532
rect 9732 27492 10416 27520
rect 9732 27480 9738 27492
rect 10410 27480 10416 27492
rect 10468 27480 10474 27532
rect 13630 27480 13636 27532
rect 13688 27520 13694 27532
rect 16022 27520 16028 27532
rect 13688 27492 16028 27520
rect 13688 27480 13694 27492
rect 16022 27480 16028 27492
rect 16080 27480 16086 27532
rect 2038 27072 2044 27124
rect 2096 27112 2102 27124
rect 5994 27112 6000 27124
rect 2096 27084 6000 27112
rect 2096 27072 2102 27084
rect 5994 27072 6000 27084
rect 6052 27072 6058 27124
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 3418 25100 3424 25152
rect 3476 25140 3482 25152
rect 6914 25140 6920 25152
rect 3476 25112 6920 25140
rect 3476 25100 3482 25112
rect 6914 25100 6920 25112
rect 6972 25100 6978 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 24762 24868 24768 24880
rect 24723 24840 24768 24868
rect 24762 24828 24768 24840
rect 24820 24828 24826 24880
rect 24026 24692 24032 24744
rect 24084 24732 24090 24744
rect 24581 24735 24639 24741
rect 24581 24732 24593 24735
rect 24084 24704 24593 24732
rect 24084 24692 24090 24704
rect 24581 24701 24593 24704
rect 24627 24732 24639 24735
rect 25133 24735 25191 24741
rect 25133 24732 25145 24735
rect 24627 24704 25145 24732
rect 24627 24701 24639 24704
rect 24581 24695 24639 24701
rect 25133 24701 25145 24704
rect 25179 24701 25191 24735
rect 25133 24695 25191 24701
rect 658 24556 664 24608
rect 716 24596 722 24608
rect 6270 24596 6276 24608
rect 716 24568 6276 24596
rect 716 24556 722 24568
rect 6270 24556 6276 24568
rect 6328 24556 6334 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1578 24392 1584 24404
rect 1539 24364 1584 24392
rect 1578 24352 1584 24364
rect 1636 24352 1642 24404
rect 17773 24395 17831 24401
rect 17773 24361 17785 24395
rect 17819 24392 17831 24395
rect 18782 24392 18788 24404
rect 17819 24364 18788 24392
rect 17819 24361 17831 24364
rect 17773 24355 17831 24361
rect 18782 24352 18788 24364
rect 18840 24352 18846 24404
rect 24765 24395 24823 24401
rect 24765 24361 24777 24395
rect 24811 24392 24823 24395
rect 25498 24392 25504 24404
rect 24811 24364 25504 24392
rect 24811 24361 24823 24364
rect 24765 24355 24823 24361
rect 25498 24352 25504 24364
rect 25556 24352 25562 24404
rect 1394 24256 1400 24268
rect 1355 24228 1400 24256
rect 1394 24216 1400 24228
rect 1452 24216 1458 24268
rect 17586 24256 17592 24268
rect 17547 24228 17592 24256
rect 17586 24216 17592 24228
rect 17644 24216 17650 24268
rect 23474 24216 23480 24268
rect 23532 24256 23538 24268
rect 24581 24259 24639 24265
rect 23532 24228 23577 24256
rect 23532 24216 23538 24228
rect 24581 24225 24593 24259
rect 24627 24256 24639 24259
rect 24670 24256 24676 24268
rect 24627 24228 24676 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 24670 24216 24676 24228
rect 24728 24216 24734 24268
rect 23661 24123 23719 24129
rect 23661 24089 23673 24123
rect 23707 24120 23719 24123
rect 25774 24120 25780 24132
rect 23707 24092 25780 24120
rect 23707 24089 23719 24092
rect 23661 24083 23719 24089
rect 25774 24080 25780 24092
rect 25832 24080 25838 24132
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1394 23808 1400 23860
rect 1452 23848 1458 23860
rect 1949 23851 2007 23857
rect 1949 23848 1961 23851
rect 1452 23820 1961 23848
rect 1452 23808 1458 23820
rect 1949 23817 1961 23820
rect 1995 23848 2007 23851
rect 2038 23848 2044 23860
rect 1995 23820 2044 23848
rect 1995 23817 2007 23820
rect 1949 23811 2007 23817
rect 2038 23808 2044 23820
rect 2096 23808 2102 23860
rect 12986 23848 12992 23860
rect 12947 23820 12992 23848
rect 12986 23808 12992 23820
rect 13044 23808 13050 23860
rect 14550 23848 14556 23860
rect 14511 23820 14556 23848
rect 14550 23808 14556 23820
rect 14608 23808 14614 23860
rect 16577 23851 16635 23857
rect 16577 23817 16589 23851
rect 16623 23848 16635 23851
rect 17402 23848 17408 23860
rect 16623 23820 17408 23848
rect 16623 23817 16635 23820
rect 16577 23811 16635 23817
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 17586 23848 17592 23860
rect 17547 23820 17592 23848
rect 17586 23808 17592 23820
rect 17644 23808 17650 23860
rect 19981 23851 20039 23857
rect 19981 23817 19993 23851
rect 20027 23848 20039 23851
rect 21634 23848 21640 23860
rect 20027 23820 21640 23848
rect 20027 23817 20039 23820
rect 19981 23811 20039 23817
rect 21634 23808 21640 23820
rect 21692 23808 21698 23860
rect 22005 23851 22063 23857
rect 22005 23817 22017 23851
rect 22051 23848 22063 23851
rect 23014 23848 23020 23860
rect 22051 23820 23020 23848
rect 22051 23817 22063 23820
rect 22005 23811 22063 23817
rect 23014 23808 23020 23820
rect 23072 23808 23078 23860
rect 23474 23808 23480 23860
rect 23532 23848 23538 23860
rect 23842 23848 23848 23860
rect 23532 23820 23848 23848
rect 23532 23808 23538 23820
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 24765 23851 24823 23857
rect 24765 23817 24777 23851
rect 24811 23848 24823 23851
rect 27154 23848 27160 23860
rect 24811 23820 27160 23848
rect 24811 23817 24823 23820
rect 24765 23811 24823 23817
rect 27154 23808 27160 23820
rect 27212 23808 27218 23860
rect 1486 23740 1492 23792
rect 1544 23780 1550 23792
rect 1581 23783 1639 23789
rect 1581 23780 1593 23783
rect 1544 23752 1593 23780
rect 1544 23740 1550 23752
rect 1581 23749 1593 23752
rect 1627 23749 1639 23783
rect 1581 23743 1639 23749
rect 18877 23783 18935 23789
rect 18877 23749 18889 23783
rect 18923 23780 18935 23783
rect 20162 23780 20168 23792
rect 18923 23752 20168 23780
rect 18923 23749 18935 23752
rect 18877 23743 18935 23749
rect 20162 23740 20168 23752
rect 20220 23740 20226 23792
rect 23474 23672 23480 23724
rect 23532 23712 23538 23724
rect 24670 23712 24676 23724
rect 23532 23684 24676 23712
rect 23532 23672 23538 23684
rect 24670 23672 24676 23684
rect 24728 23712 24734 23724
rect 25133 23715 25191 23721
rect 25133 23712 25145 23715
rect 24728 23684 25145 23712
rect 24728 23672 24734 23684
rect 25133 23681 25145 23684
rect 25179 23681 25191 23715
rect 25133 23675 25191 23681
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 12504 23647 12562 23653
rect 1443 23616 2452 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 2424 23517 2452 23616
rect 12504 23613 12516 23647
rect 12550 23644 12562 23647
rect 12986 23644 12992 23656
rect 12550 23616 12992 23644
rect 12550 23613 12562 23616
rect 12504 23607 12562 23613
rect 12986 23604 12992 23616
rect 13044 23604 13050 23656
rect 14068 23647 14126 23653
rect 14068 23613 14080 23647
rect 14114 23644 14126 23647
rect 14550 23644 14556 23656
rect 14114 23616 14556 23644
rect 14114 23613 14126 23616
rect 14068 23607 14126 23613
rect 14550 23604 14556 23616
rect 14608 23604 14614 23656
rect 16390 23644 16396 23656
rect 16303 23616 16396 23644
rect 16390 23604 16396 23616
rect 16448 23644 16454 23656
rect 16945 23647 17003 23653
rect 16945 23644 16957 23647
rect 16448 23616 16957 23644
rect 16448 23604 16454 23616
rect 16945 23613 16957 23616
rect 16991 23613 17003 23647
rect 16945 23607 17003 23613
rect 18693 23647 18751 23653
rect 18693 23613 18705 23647
rect 18739 23644 18751 23647
rect 19242 23644 19248 23656
rect 18739 23616 19248 23644
rect 18739 23613 18751 23616
rect 18693 23607 18751 23613
rect 19242 23604 19248 23616
rect 19300 23604 19306 23656
rect 19518 23604 19524 23656
rect 19576 23644 19582 23656
rect 19797 23647 19855 23653
rect 19797 23644 19809 23647
rect 19576 23616 19809 23644
rect 19576 23604 19582 23616
rect 19797 23613 19809 23616
rect 19843 23644 19855 23647
rect 20349 23647 20407 23653
rect 20349 23644 20361 23647
rect 19843 23616 20361 23644
rect 19843 23613 19855 23616
rect 19797 23607 19855 23613
rect 20349 23613 20361 23616
rect 20395 23613 20407 23647
rect 20349 23607 20407 23613
rect 21821 23647 21879 23653
rect 21821 23613 21833 23647
rect 21867 23613 21879 23647
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 21821 23607 21879 23613
rect 24412 23616 24593 23644
rect 20254 23536 20260 23588
rect 20312 23576 20318 23588
rect 21836 23576 21864 23607
rect 22373 23579 22431 23585
rect 22373 23576 22385 23579
rect 20312 23548 22385 23576
rect 20312 23536 20318 23548
rect 22373 23545 22385 23548
rect 22419 23576 22431 23579
rect 24026 23576 24032 23588
rect 22419 23548 24032 23576
rect 22419 23545 22431 23548
rect 22373 23539 22431 23545
rect 24026 23536 24032 23548
rect 24084 23536 24090 23588
rect 2409 23511 2467 23517
rect 2409 23477 2421 23511
rect 2455 23508 2467 23511
rect 2958 23508 2964 23520
rect 2455 23480 2964 23508
rect 2455 23477 2467 23480
rect 2409 23471 2467 23477
rect 2958 23468 2964 23480
rect 3016 23468 3022 23520
rect 12342 23468 12348 23520
rect 12400 23508 12406 23520
rect 12575 23511 12633 23517
rect 12575 23508 12587 23511
rect 12400 23480 12587 23508
rect 12400 23468 12406 23480
rect 12575 23477 12587 23480
rect 12621 23477 12633 23511
rect 12575 23471 12633 23477
rect 13538 23468 13544 23520
rect 13596 23508 13602 23520
rect 14139 23511 14197 23517
rect 14139 23508 14151 23511
rect 13596 23480 14151 23508
rect 13596 23468 13602 23480
rect 14139 23477 14151 23480
rect 14185 23477 14197 23511
rect 14139 23471 14197 23477
rect 24210 23468 24216 23520
rect 24268 23508 24274 23520
rect 24412 23517 24440 23616
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 24268 23480 24409 23508
rect 24268 23468 24274 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24397 23471 24455 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1578 23304 1584 23316
rect 1539 23276 1584 23304
rect 1578 23264 1584 23276
rect 1636 23264 1642 23316
rect 11655 23307 11713 23313
rect 11655 23273 11667 23307
rect 11701 23304 11713 23307
rect 15102 23304 15108 23316
rect 11701 23276 15108 23304
rect 11701 23273 11713 23276
rect 11655 23267 11713 23273
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 15427 23307 15485 23313
rect 15427 23273 15439 23307
rect 15473 23304 15485 23307
rect 16390 23304 16396 23316
rect 15473 23276 16396 23304
rect 15473 23273 15485 23276
rect 15427 23267 15485 23273
rect 16390 23264 16396 23276
rect 16448 23264 16454 23316
rect 23477 23307 23535 23313
rect 23477 23273 23489 23307
rect 23523 23304 23535 23307
rect 24118 23304 24124 23316
rect 23523 23276 24124 23304
rect 23523 23273 23535 23276
rect 23477 23267 23535 23273
rect 24118 23264 24124 23276
rect 24176 23264 24182 23316
rect 24765 23307 24823 23313
rect 24765 23273 24777 23307
rect 24811 23304 24823 23307
rect 25222 23304 25228 23316
rect 24811 23276 25228 23304
rect 24811 23273 24823 23276
rect 24765 23267 24823 23273
rect 25222 23264 25228 23276
rect 25280 23264 25286 23316
rect 1394 23168 1400 23180
rect 1355 23140 1400 23168
rect 1394 23128 1400 23140
rect 1452 23128 1458 23180
rect 11146 23128 11152 23180
rect 11204 23168 11210 23180
rect 11552 23171 11610 23177
rect 11552 23168 11564 23171
rect 11204 23140 11564 23168
rect 11204 23128 11210 23140
rect 11552 23137 11564 23140
rect 11598 23137 11610 23171
rect 11552 23131 11610 23137
rect 15197 23171 15255 23177
rect 15197 23137 15209 23171
rect 15243 23168 15255 23171
rect 15286 23168 15292 23180
rect 15243 23140 15292 23168
rect 15243 23137 15255 23140
rect 15197 23131 15255 23137
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 23290 23168 23296 23180
rect 23251 23140 23296 23168
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 24118 23128 24124 23180
rect 24176 23168 24182 23180
rect 24581 23171 24639 23177
rect 24581 23168 24593 23171
rect 24176 23140 24593 23168
rect 24176 23128 24182 23140
rect 24581 23137 24593 23140
rect 24627 23137 24639 23171
rect 24581 23131 24639 23137
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 23290 22760 23296 22772
rect 23251 22732 23296 22760
rect 23290 22720 23296 22732
rect 23348 22720 23354 22772
rect 24762 22760 24768 22772
rect 24723 22732 24768 22760
rect 24762 22720 24768 22732
rect 24820 22720 24826 22772
rect 23382 22516 23388 22568
rect 23440 22556 23446 22568
rect 24118 22556 24124 22568
rect 23440 22528 24124 22556
rect 23440 22516 23446 22528
rect 24118 22516 24124 22528
rect 24176 22556 24182 22568
rect 24397 22559 24455 22565
rect 24397 22556 24409 22559
rect 24176 22528 24409 22556
rect 24176 22516 24182 22528
rect 24397 22525 24409 22528
rect 24443 22525 24455 22559
rect 24397 22519 24455 22525
rect 24581 22559 24639 22565
rect 24581 22525 24593 22559
rect 24627 22525 24639 22559
rect 24581 22519 24639 22525
rect 24596 22488 24624 22519
rect 25133 22491 25191 22497
rect 25133 22488 25145 22491
rect 24044 22460 25145 22488
rect 24044 22432 24072 22460
rect 25133 22457 25145 22460
rect 25179 22457 25191 22491
rect 25133 22451 25191 22457
rect 1394 22380 1400 22432
rect 1452 22420 1458 22432
rect 1673 22423 1731 22429
rect 1673 22420 1685 22423
rect 1452 22392 1685 22420
rect 1452 22380 1458 22392
rect 1673 22389 1685 22392
rect 1719 22420 1731 22423
rect 9030 22420 9036 22432
rect 1719 22392 9036 22420
rect 1719 22389 1731 22392
rect 1673 22383 1731 22389
rect 9030 22380 9036 22392
rect 9088 22380 9094 22432
rect 11146 22380 11152 22432
rect 11204 22420 11210 22432
rect 11517 22423 11575 22429
rect 11517 22420 11529 22423
rect 11204 22392 11529 22420
rect 11204 22380 11210 22392
rect 11517 22389 11529 22392
rect 11563 22389 11575 22423
rect 11517 22383 11575 22389
rect 13906 22380 13912 22432
rect 13964 22420 13970 22432
rect 15286 22420 15292 22432
rect 13964 22392 15292 22420
rect 13964 22380 13970 22392
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 23290 22380 23296 22432
rect 23348 22420 23354 22432
rect 24026 22420 24032 22432
rect 23348 22392 24032 22420
rect 23348 22380 23354 22392
rect 24026 22380 24032 22392
rect 24084 22380 24090 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1464 22083 1522 22089
rect 1464 22049 1476 22083
rect 1510 22080 1522 22083
rect 1946 22080 1952 22092
rect 1510 22052 1952 22080
rect 1510 22049 1522 22052
rect 1464 22043 1522 22049
rect 1946 22040 1952 22052
rect 2004 22040 2010 22092
rect 2038 22040 2044 22092
rect 2096 22080 2102 22092
rect 2476 22083 2534 22089
rect 2476 22080 2488 22083
rect 2096 22052 2488 22080
rect 2096 22040 2102 22052
rect 2476 22049 2488 22052
rect 2522 22080 2534 22083
rect 3050 22080 3056 22092
rect 2522 22052 3056 22080
rect 2522 22049 2534 22052
rect 2476 22043 2534 22049
rect 3050 22040 3056 22052
rect 3108 22040 3114 22092
rect 1535 21947 1593 21953
rect 1535 21913 1547 21947
rect 1581 21944 1593 21947
rect 3510 21944 3516 21956
rect 1581 21916 3516 21944
rect 1581 21913 1593 21916
rect 1535 21907 1593 21913
rect 3510 21904 3516 21916
rect 3568 21904 3574 21956
rect 1762 21836 1768 21888
rect 1820 21876 1826 21888
rect 2547 21879 2605 21885
rect 2547 21876 2559 21879
rect 1820 21848 2559 21876
rect 1820 21836 1826 21848
rect 2547 21845 2559 21848
rect 2593 21845 2605 21879
rect 2547 21839 2605 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1486 21632 1492 21684
rect 1544 21672 1550 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1544 21644 1593 21672
rect 1544 21632 1550 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 1581 21635 1639 21641
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 3050 21536 3056 21548
rect 3011 21508 3056 21536
rect 3050 21496 3056 21508
rect 3108 21496 3114 21548
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21437 1455 21471
rect 1397 21431 1455 21437
rect 24581 21471 24639 21477
rect 24581 21437 24593 21471
rect 24627 21468 24639 21471
rect 24670 21468 24676 21480
rect 24627 21440 24676 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 1412 21400 1440 21431
rect 24670 21428 24676 21440
rect 24728 21468 24734 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24728 21440 25145 21468
rect 24728 21428 24734 21440
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 2409 21403 2467 21409
rect 2409 21400 2421 21403
rect 1412 21372 2421 21400
rect 2409 21369 2421 21372
rect 2455 21400 2467 21403
rect 4982 21400 4988 21412
rect 2455 21372 4988 21400
rect 2455 21369 2467 21372
rect 2409 21363 2467 21369
rect 4982 21360 4988 21372
rect 5040 21360 5046 21412
rect 1946 21332 1952 21344
rect 1907 21304 1952 21332
rect 1946 21292 1952 21304
rect 2004 21292 2010 21344
rect 2498 21332 2504 21344
rect 2459 21304 2504 21332
rect 2498 21292 2504 21304
rect 2556 21292 2562 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1578 21128 1584 21140
rect 1539 21100 1584 21128
rect 1578 21088 1584 21100
rect 1636 21088 1642 21140
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 2038 20992 2044 21004
rect 1443 20964 2044 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 2038 20952 2044 20964
rect 2096 20952 2102 21004
rect 2547 20995 2605 21001
rect 2547 20961 2559 20995
rect 2593 20961 2605 20995
rect 2547 20955 2605 20961
rect 1210 20884 1216 20936
rect 1268 20924 1274 20936
rect 2562 20924 2590 20955
rect 3326 20924 3332 20936
rect 1268 20896 3332 20924
rect 1268 20884 1274 20896
rect 3326 20884 3332 20896
rect 3384 20884 3390 20936
rect 2130 20748 2136 20800
rect 2188 20788 2194 20800
rect 2639 20791 2697 20797
rect 2639 20788 2651 20791
rect 2188 20760 2651 20788
rect 2188 20748 2194 20760
rect 2639 20757 2651 20760
rect 2685 20757 2697 20791
rect 2639 20751 2697 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1302 20544 1308 20596
rect 1360 20584 1366 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 1360 20556 1593 20584
rect 1360 20544 1366 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 3326 20584 3332 20596
rect 3287 20556 3332 20584
rect 1581 20547 1639 20553
rect 3326 20544 3332 20556
rect 3384 20544 3390 20596
rect 24765 20587 24823 20593
rect 24765 20553 24777 20587
rect 24811 20584 24823 20587
rect 24854 20584 24860 20596
rect 24811 20556 24860 20584
rect 24811 20553 24823 20556
rect 24765 20547 24823 20553
rect 24854 20544 24860 20556
rect 24912 20544 24918 20596
rect 3053 20451 3111 20457
rect 3053 20417 3065 20451
rect 3099 20448 3111 20451
rect 3786 20448 3792 20460
rect 3099 20420 3792 20448
rect 3099 20417 3111 20420
rect 3053 20411 3111 20417
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 2568 20383 2626 20389
rect 1443 20352 2452 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 2424 20256 2452 20352
rect 2568 20349 2580 20383
rect 2614 20380 2626 20383
rect 2958 20380 2964 20392
rect 2614 20352 2964 20380
rect 2614 20349 2626 20352
rect 2568 20343 2626 20349
rect 2958 20340 2964 20352
rect 3016 20380 3022 20392
rect 3068 20380 3096 20411
rect 3786 20408 3792 20420
rect 3844 20408 3850 20460
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 9732 20420 13814 20448
rect 9732 20408 9738 20420
rect 3016 20352 3096 20380
rect 3564 20383 3622 20389
rect 3016 20340 3022 20352
rect 3564 20349 3576 20383
rect 3610 20380 3622 20383
rect 3970 20380 3976 20392
rect 3610 20352 3976 20380
rect 3610 20349 3622 20352
rect 3564 20343 3622 20349
rect 3970 20340 3976 20352
rect 4028 20340 4034 20392
rect 9585 20383 9643 20389
rect 9585 20349 9597 20383
rect 9631 20380 9643 20383
rect 13786 20380 13814 20420
rect 15048 20383 15106 20389
rect 15048 20380 15060 20383
rect 9631 20352 9996 20380
rect 13786 20352 15060 20380
rect 9631 20349 9643 20352
rect 9585 20343 9643 20349
rect 3142 20272 3148 20324
rect 3200 20312 3206 20324
rect 3651 20315 3709 20321
rect 3651 20312 3663 20315
rect 3200 20284 3663 20312
rect 3200 20272 3206 20284
rect 3651 20281 3663 20284
rect 3697 20281 3709 20315
rect 3651 20275 3709 20281
rect 9968 20256 9996 20352
rect 15048 20349 15060 20352
rect 15094 20380 15106 20383
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 15094 20352 15485 20380
rect 15094 20349 15106 20352
rect 15048 20343 15106 20349
rect 15473 20349 15485 20352
rect 15519 20349 15531 20383
rect 15473 20343 15531 20349
rect 24118 20340 24124 20392
rect 24176 20380 24182 20392
rect 24581 20383 24639 20389
rect 24581 20380 24593 20383
rect 24176 20352 24593 20380
rect 24176 20340 24182 20352
rect 24581 20349 24593 20352
rect 24627 20380 24639 20383
rect 25133 20383 25191 20389
rect 25133 20380 25145 20383
rect 24627 20352 25145 20380
rect 24627 20349 24639 20352
rect 24581 20343 24639 20349
rect 25133 20349 25145 20352
rect 25179 20349 25191 20383
rect 25133 20343 25191 20349
rect 2038 20244 2044 20256
rect 1999 20216 2044 20244
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 2406 20244 2412 20256
rect 2367 20216 2412 20244
rect 2406 20204 2412 20216
rect 2464 20204 2470 20256
rect 2639 20247 2697 20253
rect 2639 20213 2651 20247
rect 2685 20244 2697 20247
rect 2866 20244 2872 20256
rect 2685 20216 2872 20244
rect 2685 20213 2697 20216
rect 2639 20207 2697 20213
rect 2866 20204 2872 20216
rect 2924 20204 2930 20256
rect 9769 20247 9827 20253
rect 9769 20213 9781 20247
rect 9815 20244 9827 20247
rect 9858 20244 9864 20256
rect 9815 20216 9864 20244
rect 9815 20213 9827 20216
rect 9769 20207 9827 20213
rect 9858 20204 9864 20216
rect 9916 20204 9922 20256
rect 9950 20204 9956 20256
rect 10008 20244 10014 20256
rect 10045 20247 10103 20253
rect 10045 20244 10057 20247
rect 10008 20216 10057 20244
rect 10008 20204 10014 20216
rect 10045 20213 10057 20216
rect 10091 20213 10103 20247
rect 10045 20207 10103 20213
rect 15151 20247 15209 20253
rect 15151 20213 15163 20247
rect 15197 20244 15209 20247
rect 16298 20244 16304 20256
rect 15197 20216 16304 20244
rect 15197 20213 15209 20216
rect 15151 20207 15209 20213
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 198 20000 204 20052
rect 256 20040 262 20052
rect 1581 20043 1639 20049
rect 1581 20040 1593 20043
rect 256 20012 1593 20040
rect 256 20000 262 20012
rect 1581 20009 1593 20012
rect 1627 20009 1639 20043
rect 1581 20003 1639 20009
rect 2406 20000 2412 20052
rect 2464 20040 2470 20052
rect 4203 20043 4261 20049
rect 4203 20040 4215 20043
rect 2464 20012 4215 20040
rect 2464 20000 2470 20012
rect 4203 20009 4215 20012
rect 4249 20009 4261 20043
rect 4203 20003 4261 20009
rect 4982 20000 4988 20052
rect 5040 20040 5046 20052
rect 5215 20043 5273 20049
rect 5215 20040 5227 20043
rect 5040 20012 5227 20040
rect 5040 20000 5046 20012
rect 5215 20009 5227 20012
rect 5261 20009 5273 20043
rect 5215 20003 5273 20009
rect 19242 19932 19248 19984
rect 19300 19972 19306 19984
rect 22462 19972 22468 19984
rect 19300 19944 22468 19972
rect 19300 19932 19306 19944
rect 22462 19932 22468 19944
rect 22520 19932 22526 19984
rect 1394 19904 1400 19916
rect 1355 19876 1400 19904
rect 1394 19864 1400 19876
rect 1452 19864 1458 19916
rect 2501 19907 2559 19913
rect 2501 19873 2513 19907
rect 2547 19904 2559 19907
rect 2774 19904 2780 19916
rect 2547 19876 2780 19904
rect 2547 19873 2559 19876
rect 2501 19867 2559 19873
rect 2774 19864 2780 19876
rect 2832 19864 2838 19916
rect 4132 19907 4190 19913
rect 4132 19873 4144 19907
rect 4178 19904 4190 19907
rect 4614 19904 4620 19916
rect 4178 19876 4620 19904
rect 4178 19873 4190 19876
rect 4132 19867 4190 19873
rect 4614 19864 4620 19876
rect 4672 19864 4678 19916
rect 5144 19907 5202 19913
rect 5144 19873 5156 19907
rect 5190 19904 5202 19907
rect 5350 19904 5356 19916
rect 5190 19876 5356 19904
rect 5190 19873 5202 19876
rect 5144 19867 5202 19873
rect 5350 19864 5356 19876
rect 5408 19864 5414 19916
rect 6086 19864 6092 19916
rect 6144 19904 6150 19916
rect 6952 19907 7010 19913
rect 6952 19904 6964 19907
rect 6144 19876 6964 19904
rect 6144 19864 6150 19876
rect 6952 19873 6964 19876
rect 6998 19904 7010 19907
rect 7650 19904 7656 19916
rect 6998 19876 7656 19904
rect 6998 19873 7010 19876
rect 6952 19867 7010 19873
rect 7650 19864 7656 19876
rect 7708 19864 7714 19916
rect 7929 19907 7987 19913
rect 7929 19873 7941 19907
rect 7975 19904 7987 19907
rect 8018 19904 8024 19916
rect 7975 19876 8024 19904
rect 7975 19873 7987 19876
rect 7929 19867 7987 19873
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 8938 19864 8944 19916
rect 8996 19904 9002 19916
rect 9712 19907 9770 19913
rect 9712 19904 9724 19907
rect 8996 19876 9724 19904
rect 8996 19864 9002 19876
rect 9712 19873 9724 19876
rect 9758 19873 9770 19907
rect 9712 19867 9770 19873
rect 10756 19907 10814 19913
rect 10756 19873 10768 19907
rect 10802 19904 10814 19907
rect 11422 19904 11428 19916
rect 10802 19876 11428 19904
rect 10802 19873 10814 19876
rect 10756 19867 10814 19873
rect 11422 19864 11428 19876
rect 11480 19864 11486 19916
rect 13998 19864 14004 19916
rect 14056 19904 14062 19916
rect 14220 19907 14278 19913
rect 14220 19904 14232 19907
rect 14056 19876 14232 19904
rect 14056 19864 14062 19876
rect 14220 19873 14232 19876
rect 14266 19873 14278 19907
rect 14220 19867 14278 19873
rect 15356 19907 15414 19913
rect 15356 19873 15368 19907
rect 15402 19904 15414 19907
rect 15562 19904 15568 19916
rect 15402 19876 15568 19904
rect 15402 19873 15414 19876
rect 15356 19867 15414 19873
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 18046 19904 18052 19916
rect 18007 19876 18052 19904
rect 18046 19864 18052 19876
rect 18104 19864 18110 19916
rect 18598 19904 18604 19916
rect 18559 19876 18604 19904
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 19648 19907 19706 19913
rect 19648 19904 19660 19907
rect 19484 19876 19660 19904
rect 19484 19864 19490 19876
rect 19648 19873 19660 19876
rect 19694 19873 19706 19907
rect 19648 19867 19706 19873
rect 18782 19836 18788 19848
rect 18743 19808 18788 19836
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 2682 19768 2688 19780
rect 2643 19740 2688 19768
rect 2682 19728 2688 19740
rect 2740 19728 2746 19780
rect 13722 19728 13728 19780
rect 13780 19768 13786 19780
rect 14645 19771 14703 19777
rect 14645 19768 14657 19771
rect 13780 19740 14657 19768
rect 13780 19728 13786 19740
rect 14645 19737 14657 19740
rect 14691 19737 14703 19771
rect 14645 19731 14703 19737
rect 15427 19771 15485 19777
rect 15427 19737 15439 19771
rect 15473 19768 15485 19771
rect 17862 19768 17868 19780
rect 15473 19740 17868 19768
rect 15473 19737 15485 19740
rect 15427 19731 15485 19737
rect 17862 19728 17868 19740
rect 17920 19728 17926 19780
rect 19242 19728 19248 19780
rect 19300 19768 19306 19780
rect 20073 19771 20131 19777
rect 20073 19768 20085 19771
rect 19300 19740 20085 19768
rect 19300 19728 19306 19740
rect 20073 19737 20085 19740
rect 20119 19737 20131 19771
rect 20073 19731 20131 19737
rect 4614 19700 4620 19712
rect 4575 19672 4620 19700
rect 4614 19660 4620 19672
rect 4672 19660 4678 19712
rect 7055 19703 7113 19709
rect 7055 19669 7067 19703
rect 7101 19700 7113 19703
rect 7926 19700 7932 19712
rect 7101 19672 7932 19700
rect 7101 19669 7113 19672
rect 7055 19663 7113 19669
rect 7926 19660 7932 19672
rect 7984 19660 7990 19712
rect 8067 19703 8125 19709
rect 8067 19669 8079 19703
rect 8113 19700 8125 19703
rect 8478 19700 8484 19712
rect 8113 19672 8484 19700
rect 8113 19669 8125 19672
rect 8067 19663 8125 19669
rect 8478 19660 8484 19672
rect 8536 19660 8542 19712
rect 9815 19703 9873 19709
rect 9815 19669 9827 19703
rect 9861 19700 9873 19703
rect 10134 19700 10140 19712
rect 9861 19672 10140 19700
rect 9861 19669 9873 19672
rect 9815 19663 9873 19669
rect 10134 19660 10140 19672
rect 10192 19660 10198 19712
rect 10827 19703 10885 19709
rect 10827 19669 10839 19703
rect 10873 19700 10885 19703
rect 10962 19700 10968 19712
rect 10873 19672 10968 19700
rect 10873 19669 10885 19672
rect 10827 19663 10885 19669
rect 10962 19660 10968 19672
rect 11020 19660 11026 19712
rect 14182 19660 14188 19712
rect 14240 19700 14246 19712
rect 14323 19703 14381 19709
rect 14323 19700 14335 19703
rect 14240 19672 14335 19700
rect 14240 19660 14246 19672
rect 14323 19669 14335 19672
rect 14369 19669 14381 19703
rect 16206 19700 16212 19712
rect 16167 19672 16212 19700
rect 14323 19663 14381 19669
rect 16206 19660 16212 19672
rect 16264 19660 16270 19712
rect 19751 19703 19809 19709
rect 19751 19669 19763 19703
rect 19797 19700 19809 19703
rect 19978 19700 19984 19712
rect 19797 19672 19984 19700
rect 19797 19669 19809 19672
rect 19751 19663 19809 19669
rect 19978 19660 19984 19672
rect 20036 19660 20042 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 7650 19496 7656 19508
rect 7611 19468 7656 19496
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 8018 19456 8024 19508
rect 8076 19496 8082 19508
rect 8573 19499 8631 19505
rect 8573 19496 8585 19499
rect 8076 19468 8585 19496
rect 8076 19456 8082 19468
rect 8573 19465 8585 19468
rect 8619 19465 8631 19499
rect 8938 19496 8944 19508
rect 8899 19468 8944 19496
rect 8573 19459 8631 19465
rect 8938 19456 8944 19468
rect 8996 19496 9002 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 8996 19468 10241 19496
rect 8996 19456 9002 19468
rect 10229 19465 10241 19468
rect 10275 19465 10287 19499
rect 13630 19496 13636 19508
rect 13591 19468 13636 19496
rect 10229 19459 10287 19465
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 15746 19456 15752 19508
rect 15804 19496 15810 19508
rect 17865 19499 17923 19505
rect 17865 19496 17877 19499
rect 15804 19468 17877 19496
rect 15804 19456 15810 19468
rect 17865 19465 17877 19468
rect 17911 19496 17923 19499
rect 18046 19496 18052 19508
rect 17911 19468 18052 19496
rect 17911 19465 17923 19468
rect 17865 19459 17923 19465
rect 18046 19456 18052 19468
rect 18104 19456 18110 19508
rect 24762 19496 24768 19508
rect 24723 19468 24768 19496
rect 24762 19456 24768 19468
rect 24820 19456 24826 19508
rect 4706 19360 4712 19372
rect 4632 19332 4712 19360
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 1670 19292 1676 19304
rect 1443 19264 1676 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 2038 19252 2044 19304
rect 2096 19292 2102 19304
rect 4632 19301 4660 19332
rect 4706 19320 4712 19332
rect 4764 19320 4770 19372
rect 6914 19360 6920 19372
rect 6827 19332 6920 19360
rect 6907 19320 6920 19332
rect 6972 19360 6978 19372
rect 7374 19360 7380 19372
rect 6972 19332 7380 19360
rect 6972 19320 6978 19332
rect 7374 19320 7380 19332
rect 7432 19320 7438 19372
rect 19426 19360 19432 19372
rect 19387 19332 19432 19360
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 6907 19306 6960 19320
rect 2568 19295 2626 19301
rect 2568 19292 2580 19295
rect 2096 19264 2580 19292
rect 2096 19252 2102 19264
rect 2568 19261 2580 19264
rect 2614 19292 2626 19295
rect 2869 19295 2927 19301
rect 2869 19292 2881 19295
rect 2614 19264 2881 19292
rect 2614 19261 2626 19264
rect 2568 19255 2626 19261
rect 2869 19261 2881 19264
rect 2915 19261 2927 19295
rect 2869 19255 2927 19261
rect 4249 19295 4307 19301
rect 4249 19261 4261 19295
rect 4295 19292 4307 19295
rect 4617 19295 4675 19301
rect 4617 19292 4629 19295
rect 4295 19264 4629 19292
rect 4295 19261 4307 19264
rect 4249 19255 4307 19261
rect 4617 19261 4629 19264
rect 4663 19261 4675 19295
rect 4617 19255 4675 19261
rect 4893 19295 4951 19301
rect 4893 19261 4905 19295
rect 4939 19261 4951 19295
rect 4893 19255 4951 19261
rect 1486 19184 1492 19236
rect 1544 19224 1550 19236
rect 1949 19227 2007 19233
rect 1949 19224 1961 19227
rect 1544 19196 1961 19224
rect 1544 19184 1550 19196
rect 1949 19193 1961 19196
rect 1995 19193 2007 19227
rect 1949 19187 2007 19193
rect 2774 19184 2780 19236
rect 2832 19224 2838 19236
rect 2961 19227 3019 19233
rect 2961 19224 2973 19227
rect 2832 19196 2973 19224
rect 2832 19184 2838 19196
rect 2961 19193 2973 19196
rect 3007 19224 3019 19227
rect 4908 19224 4936 19255
rect 4982 19224 4988 19236
rect 3007 19196 4752 19224
rect 4908 19196 4988 19224
rect 3007 19193 3019 19196
rect 2961 19187 3019 19193
rect 198 19116 204 19168
rect 256 19156 262 19168
rect 1581 19159 1639 19165
rect 1581 19156 1593 19159
rect 256 19128 1593 19156
rect 256 19116 262 19128
rect 1581 19125 1593 19128
rect 1627 19125 1639 19159
rect 1581 19119 1639 19125
rect 2406 19116 2412 19168
rect 2464 19156 2470 19168
rect 2639 19159 2697 19165
rect 2639 19156 2651 19159
rect 2464 19128 2651 19156
rect 2464 19116 2470 19128
rect 2639 19125 2651 19128
rect 2685 19125 2697 19159
rect 2639 19119 2697 19125
rect 2869 19159 2927 19165
rect 2869 19125 2881 19159
rect 2915 19156 2927 19159
rect 3421 19159 3479 19165
rect 3421 19156 3433 19159
rect 2915 19128 3433 19156
rect 2915 19125 2927 19128
rect 2869 19119 2927 19125
rect 3421 19125 3433 19128
rect 3467 19156 3479 19159
rect 3694 19156 3700 19168
rect 3467 19128 3700 19156
rect 3467 19125 3479 19128
rect 3421 19119 3479 19125
rect 3694 19116 3700 19128
rect 3752 19116 3758 19168
rect 3878 19156 3884 19168
rect 3839 19128 3884 19156
rect 3878 19116 3884 19128
rect 3936 19116 3942 19168
rect 4338 19116 4344 19168
rect 4396 19156 4402 19168
rect 4433 19159 4491 19165
rect 4433 19156 4445 19159
rect 4396 19128 4445 19156
rect 4396 19116 4402 19128
rect 4433 19125 4445 19128
rect 4479 19125 4491 19159
rect 4724 19156 4752 19196
rect 4982 19184 4988 19196
rect 5040 19184 5046 19236
rect 6641 19227 6699 19233
rect 6641 19193 6653 19227
rect 6687 19224 6699 19227
rect 6932 19224 6960 19306
rect 8180 19295 8238 19301
rect 8180 19261 8192 19295
rect 8226 19292 8238 19295
rect 8938 19292 8944 19304
rect 8226 19264 8944 19292
rect 8226 19261 8238 19264
rect 8180 19255 8238 19261
rect 8938 19252 8944 19264
rect 8996 19252 9002 19304
rect 11422 19301 11428 19304
rect 9769 19295 9827 19301
rect 9769 19292 9781 19295
rect 9600 19264 9781 19292
rect 6687 19196 6960 19224
rect 6687 19193 6699 19196
rect 6641 19187 6699 19193
rect 4798 19156 4804 19168
rect 4724 19128 4804 19156
rect 4433 19119 4491 19125
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 5350 19156 5356 19168
rect 5311 19128 5356 19156
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 6963 19159 7021 19165
rect 6963 19125 6975 19159
rect 7009 19156 7021 19159
rect 7190 19156 7196 19168
rect 7009 19128 7196 19156
rect 7009 19125 7021 19128
rect 6963 19119 7021 19125
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 8110 19116 8116 19168
rect 8168 19156 8174 19168
rect 8251 19159 8309 19165
rect 8251 19156 8263 19159
rect 8168 19128 8263 19156
rect 8168 19116 8174 19128
rect 8251 19125 8263 19128
rect 8297 19125 8309 19159
rect 8251 19119 8309 19125
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 9600 19165 9628 19264
rect 9769 19261 9781 19264
rect 9815 19261 9827 19295
rect 9769 19255 9827 19261
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19292 10839 19295
rect 11400 19295 11428 19301
rect 11400 19292 11412 19295
rect 10827 19264 11412 19292
rect 10827 19261 10839 19264
rect 10781 19255 10839 19261
rect 11400 19261 11412 19264
rect 11480 19292 11486 19304
rect 11793 19295 11851 19301
rect 11793 19292 11805 19295
rect 11480 19264 11805 19292
rect 11400 19255 11428 19261
rect 11422 19252 11428 19255
rect 11480 19252 11486 19264
rect 11793 19261 11805 19264
rect 11839 19261 11851 19295
rect 11793 19255 11851 19261
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19261 13507 19295
rect 13449 19255 13507 19261
rect 13464 19168 13492 19255
rect 13722 19252 13728 19304
rect 13780 19292 13786 19304
rect 14366 19292 14372 19304
rect 13780 19264 14372 19292
rect 13780 19252 13786 19264
rect 14366 19252 14372 19264
rect 14424 19292 14430 19304
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 14424 19264 14565 19292
rect 14424 19252 14430 19264
rect 14553 19261 14565 19264
rect 14599 19261 14611 19295
rect 14553 19255 14611 19261
rect 14642 19252 14648 19304
rect 14700 19292 14706 19304
rect 15013 19295 15071 19301
rect 15013 19292 15025 19295
rect 14700 19264 15025 19292
rect 14700 19252 14706 19264
rect 15013 19261 15025 19264
rect 15059 19261 15071 19295
rect 15013 19255 15071 19261
rect 17494 19252 17500 19304
rect 17552 19292 17558 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17552 19264 18061 19292
rect 17552 19252 17558 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18598 19292 18604 19304
rect 18511 19264 18604 19292
rect 18049 19255 18107 19261
rect 18598 19252 18604 19264
rect 18656 19252 18662 19304
rect 19242 19252 19248 19304
rect 19300 19292 19306 19304
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 19300 19264 19625 19292
rect 19300 19252 19306 19264
rect 19613 19261 19625 19264
rect 19659 19261 19671 19295
rect 20070 19292 20076 19304
rect 20031 19264 20076 19292
rect 19613 19255 19671 19261
rect 20070 19252 20076 19264
rect 20128 19252 20134 19304
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 24581 19295 24639 19301
rect 24581 19292 24593 19295
rect 20772 19264 24593 19292
rect 20772 19252 20778 19264
rect 24581 19261 24593 19264
rect 24627 19292 24639 19295
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 24627 19264 25145 19292
rect 24627 19261 24639 19264
rect 24581 19255 24639 19261
rect 25133 19261 25145 19264
rect 25179 19261 25191 19295
rect 25133 19255 25191 19261
rect 15286 19224 15292 19236
rect 15247 19196 15292 19224
rect 15286 19184 15292 19196
rect 15344 19184 15350 19236
rect 16206 19224 16212 19236
rect 16167 19196 16212 19224
rect 16206 19184 16212 19196
rect 16264 19184 16270 19236
rect 16301 19227 16359 19233
rect 16301 19193 16313 19227
rect 16347 19224 16359 19227
rect 16482 19224 16488 19236
rect 16347 19196 16488 19224
rect 16347 19193 16359 19196
rect 16301 19187 16359 19193
rect 9585 19159 9643 19165
rect 9585 19156 9597 19159
rect 9364 19128 9597 19156
rect 9364 19116 9370 19128
rect 9585 19125 9597 19128
rect 9631 19125 9643 19159
rect 9585 19119 9643 19125
rect 9766 19116 9772 19168
rect 9824 19156 9830 19168
rect 9953 19159 10011 19165
rect 9953 19156 9965 19159
rect 9824 19128 9965 19156
rect 9824 19116 9830 19128
rect 9953 19125 9965 19128
rect 9999 19125 10011 19159
rect 9953 19119 10011 19125
rect 11471 19159 11529 19165
rect 11471 19125 11483 19159
rect 11517 19156 11529 19159
rect 12986 19156 12992 19168
rect 11517 19128 12992 19156
rect 11517 19125 11529 19128
rect 11471 19119 11529 19125
rect 12986 19116 12992 19128
rect 13044 19116 13050 19168
rect 13357 19159 13415 19165
rect 13357 19125 13369 19159
rect 13403 19156 13415 19159
rect 13446 19156 13452 19168
rect 13403 19128 13452 19156
rect 13403 19125 13415 19128
rect 13357 19119 13415 19125
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 13998 19116 14004 19168
rect 14056 19156 14062 19168
rect 14185 19159 14243 19165
rect 14185 19156 14197 19159
rect 14056 19128 14197 19156
rect 14056 19116 14062 19128
rect 14185 19125 14197 19128
rect 14231 19125 14243 19159
rect 15562 19156 15568 19168
rect 15523 19128 15568 19156
rect 14185 19119 14243 19125
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 16025 19159 16083 19165
rect 16025 19125 16037 19159
rect 16071 19156 16083 19159
rect 16316 19156 16344 19187
rect 16482 19184 16488 19196
rect 16540 19184 16546 19236
rect 16853 19227 16911 19233
rect 16853 19193 16865 19227
rect 16899 19224 16911 19227
rect 16942 19224 16948 19236
rect 16899 19196 16948 19224
rect 16899 19193 16911 19196
rect 16853 19187 16911 19193
rect 16942 19184 16948 19196
rect 17000 19184 17006 19236
rect 17034 19184 17040 19236
rect 17092 19224 17098 19236
rect 18616 19224 18644 19252
rect 17092 19196 18644 19224
rect 17092 19184 17098 19196
rect 17494 19156 17500 19168
rect 16071 19128 16344 19156
rect 17455 19128 17500 19156
rect 16071 19125 16083 19128
rect 16025 19119 16083 19125
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 18138 19156 18144 19168
rect 18099 19128 18144 19156
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 18616 19156 18644 19196
rect 18966 19184 18972 19236
rect 19024 19224 19030 19236
rect 19024 19196 19748 19224
rect 19024 19184 19030 19196
rect 19058 19156 19064 19168
rect 18616 19128 19064 19156
rect 19058 19116 19064 19128
rect 19116 19116 19122 19168
rect 19720 19165 19748 19196
rect 19705 19159 19763 19165
rect 19705 19125 19717 19159
rect 19751 19125 19763 19159
rect 19705 19119 19763 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 3878 18912 3884 18964
rect 3936 18952 3942 18964
rect 4982 18952 4988 18964
rect 3936 18924 4988 18952
rect 3936 18912 3942 18924
rect 4982 18912 4988 18924
rect 5040 18912 5046 18964
rect 6270 18912 6276 18964
rect 6328 18952 6334 18964
rect 7650 18952 7656 18964
rect 6328 18924 7656 18952
rect 6328 18912 6334 18924
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 12342 18912 12348 18964
rect 12400 18952 12406 18964
rect 12437 18955 12495 18961
rect 12437 18952 12449 18955
rect 12400 18924 12449 18952
rect 12400 18912 12406 18924
rect 12437 18921 12449 18924
rect 12483 18921 12495 18955
rect 18414 18952 18420 18964
rect 12437 18915 12495 18921
rect 16960 18924 18420 18952
rect 16960 18896 16988 18924
rect 18414 18912 18420 18924
rect 18472 18952 18478 18964
rect 18877 18955 18935 18961
rect 18472 18924 18552 18952
rect 18472 18912 18478 18924
rect 2222 18844 2228 18896
rect 2280 18884 2286 18896
rect 2501 18887 2559 18893
rect 2501 18884 2513 18887
rect 2280 18856 2513 18884
rect 2280 18844 2286 18856
rect 2501 18853 2513 18856
rect 2547 18884 2559 18887
rect 3418 18884 3424 18896
rect 2547 18856 3424 18884
rect 2547 18853 2559 18856
rect 2501 18847 2559 18853
rect 3418 18844 3424 18856
rect 3476 18844 3482 18896
rect 4249 18887 4307 18893
rect 4249 18853 4261 18887
rect 4295 18884 4307 18887
rect 4890 18884 4896 18896
rect 4295 18856 4896 18884
rect 4295 18853 4307 18856
rect 4249 18847 4307 18853
rect 4890 18844 4896 18856
rect 4948 18844 4954 18896
rect 6546 18844 6552 18896
rect 6604 18884 6610 18896
rect 6917 18887 6975 18893
rect 6917 18884 6929 18887
rect 6604 18856 6929 18884
rect 6604 18844 6610 18856
rect 6917 18853 6929 18856
rect 6963 18853 6975 18887
rect 16298 18884 16304 18896
rect 16259 18856 16304 18884
rect 6917 18847 6975 18853
rect 16298 18844 16304 18856
rect 16356 18844 16362 18896
rect 16390 18844 16396 18896
rect 16448 18884 16454 18896
rect 16942 18884 16948 18896
rect 16448 18856 16493 18884
rect 16903 18856 16948 18884
rect 16448 18844 16454 18856
rect 16942 18844 16948 18856
rect 17000 18844 17006 18896
rect 17862 18884 17868 18896
rect 17823 18856 17868 18884
rect 17862 18844 17868 18856
rect 17920 18844 17926 18896
rect 17957 18887 18015 18893
rect 17957 18853 17969 18887
rect 18003 18884 18015 18887
rect 18046 18884 18052 18896
rect 18003 18856 18052 18884
rect 18003 18853 18015 18856
rect 17957 18847 18015 18853
rect 18046 18844 18052 18856
rect 18104 18844 18110 18896
rect 18524 18893 18552 18924
rect 18877 18921 18889 18955
rect 18923 18952 18935 18955
rect 19058 18952 19064 18964
rect 18923 18924 19064 18952
rect 18923 18921 18935 18924
rect 18877 18915 18935 18921
rect 19058 18912 19064 18924
rect 19116 18952 19122 18964
rect 19705 18955 19763 18961
rect 19705 18952 19717 18955
rect 19116 18924 19717 18952
rect 19116 18912 19122 18924
rect 19705 18921 19717 18924
rect 19751 18952 19763 18955
rect 20070 18952 20076 18964
rect 19751 18924 20076 18952
rect 19751 18921 19763 18924
rect 19705 18915 19763 18921
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 23247 18955 23305 18961
rect 23247 18921 23259 18955
rect 23293 18952 23305 18955
rect 23382 18952 23388 18964
rect 23293 18924 23388 18952
rect 23293 18921 23305 18924
rect 23247 18915 23305 18921
rect 23382 18912 23388 18924
rect 23440 18912 23446 18964
rect 18509 18887 18567 18893
rect 18509 18853 18521 18887
rect 18555 18853 18567 18887
rect 21082 18884 21088 18896
rect 21043 18856 21088 18884
rect 18509 18847 18567 18853
rect 21082 18844 21088 18856
rect 21140 18844 21146 18896
rect 5772 18819 5830 18825
rect 5772 18785 5784 18819
rect 5818 18816 5830 18819
rect 6086 18816 6092 18828
rect 5818 18788 6092 18816
rect 5818 18785 5830 18788
rect 5772 18779 5830 18785
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 8018 18776 8024 18828
rect 8076 18816 8082 18828
rect 8332 18819 8390 18825
rect 8332 18816 8344 18819
rect 8076 18788 8344 18816
rect 8076 18776 8082 18788
rect 8332 18785 8344 18788
rect 8378 18785 8390 18819
rect 8332 18779 8390 18785
rect 9585 18819 9643 18825
rect 9585 18785 9597 18819
rect 9631 18816 9643 18819
rect 9674 18816 9680 18828
rect 9631 18788 9680 18816
rect 9631 18785 9643 18788
rect 9585 18779 9643 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 11584 18819 11642 18825
rect 11584 18785 11596 18819
rect 11630 18816 11642 18819
rect 11698 18816 11704 18828
rect 11630 18788 11704 18816
rect 11630 18785 11642 18788
rect 11584 18779 11642 18785
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 12158 18776 12164 18828
rect 12216 18816 12222 18828
rect 12621 18819 12679 18825
rect 12621 18816 12633 18819
rect 12216 18788 12633 18816
rect 12216 18776 12222 18788
rect 12621 18785 12633 18788
rect 12667 18785 12679 18819
rect 12621 18779 12679 18785
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 14185 18819 14243 18825
rect 13872 18788 13917 18816
rect 13872 18776 13878 18788
rect 14185 18785 14197 18819
rect 14231 18816 14243 18819
rect 14550 18816 14556 18828
rect 14231 18788 14556 18816
rect 14231 18785 14243 18788
rect 14185 18779 14243 18785
rect 14550 18776 14556 18788
rect 14608 18776 14614 18828
rect 19797 18819 19855 18825
rect 19797 18785 19809 18819
rect 19843 18816 19855 18819
rect 19886 18816 19892 18828
rect 19843 18788 19892 18816
rect 19843 18785 19855 18788
rect 19797 18779 19855 18785
rect 19886 18776 19892 18788
rect 19944 18776 19950 18828
rect 23106 18816 23112 18828
rect 23067 18788 23112 18816
rect 23106 18776 23112 18788
rect 23164 18776 23170 18828
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18748 2467 18751
rect 2498 18748 2504 18760
rect 2455 18720 2504 18748
rect 2455 18717 2467 18720
rect 2409 18711 2467 18717
rect 2498 18708 2504 18720
rect 2556 18708 2562 18760
rect 2590 18708 2596 18760
rect 2648 18748 2654 18760
rect 2685 18751 2743 18757
rect 2685 18748 2697 18751
rect 2648 18720 2697 18748
rect 2648 18708 2654 18720
rect 2685 18717 2697 18720
rect 2731 18717 2743 18751
rect 2685 18711 2743 18717
rect 3050 18708 3056 18760
rect 3108 18748 3114 18760
rect 4154 18748 4160 18760
rect 3108 18720 4160 18748
rect 3108 18708 3114 18720
rect 4154 18708 4160 18720
rect 4212 18748 4218 18760
rect 4614 18748 4620 18760
rect 4212 18720 4257 18748
rect 4575 18720 4620 18748
rect 4212 18708 4218 18720
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 5859 18751 5917 18757
rect 5859 18717 5871 18751
rect 5905 18748 5917 18751
rect 6273 18751 6331 18757
rect 6273 18748 6285 18751
rect 5905 18720 6285 18748
rect 5905 18717 5917 18720
rect 5859 18711 5917 18717
rect 6273 18717 6285 18720
rect 6319 18748 6331 18751
rect 6825 18751 6883 18757
rect 6825 18748 6837 18751
rect 6319 18720 6837 18748
rect 6319 18717 6331 18720
rect 6273 18711 6331 18717
rect 6825 18717 6837 18720
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18748 7527 18751
rect 7558 18748 7564 18760
rect 7515 18720 7564 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 14369 18751 14427 18757
rect 14369 18717 14381 18751
rect 14415 18748 14427 18751
rect 14826 18748 14832 18760
rect 14415 18720 14832 18748
rect 14415 18717 14427 18720
rect 14369 18711 14427 18717
rect 14826 18708 14832 18720
rect 14884 18708 14890 18760
rect 8294 18640 8300 18692
rect 8352 18680 8358 18692
rect 8757 18683 8815 18689
rect 8757 18680 8769 18683
rect 8352 18652 8769 18680
rect 8352 18640 8358 18652
rect 8757 18649 8769 18652
rect 8803 18649 8815 18683
rect 19904 18680 19932 18776
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 20993 18751 21051 18757
rect 20993 18748 21005 18751
rect 20864 18720 21005 18748
rect 20864 18708 20870 18720
rect 20993 18717 21005 18720
rect 21039 18717 21051 18751
rect 21266 18748 21272 18760
rect 21227 18720 21272 18748
rect 20993 18711 21051 18717
rect 21266 18708 21272 18720
rect 21324 18708 21330 18760
rect 24118 18680 24124 18692
rect 19904 18652 24124 18680
rect 8757 18643 8815 18649
rect 24118 18640 24124 18652
rect 24176 18640 24182 18692
rect 1670 18612 1676 18624
rect 1583 18584 1676 18612
rect 1670 18572 1676 18584
rect 1728 18612 1734 18624
rect 2314 18612 2320 18624
rect 1728 18584 2320 18612
rect 1728 18572 1734 18584
rect 2314 18572 2320 18584
rect 2372 18572 2378 18624
rect 6546 18612 6552 18624
rect 6507 18584 6552 18612
rect 6546 18572 6552 18584
rect 6604 18572 6610 18624
rect 7282 18572 7288 18624
rect 7340 18612 7346 18624
rect 8435 18615 8493 18621
rect 8435 18612 8447 18615
rect 7340 18584 8447 18612
rect 7340 18572 7346 18584
rect 8435 18581 8447 18584
rect 8481 18581 8493 18615
rect 8435 18575 8493 18581
rect 9815 18615 9873 18621
rect 9815 18581 9827 18615
rect 9861 18612 9873 18615
rect 10229 18615 10287 18621
rect 10229 18612 10241 18615
rect 9861 18584 10241 18612
rect 9861 18581 9873 18584
rect 9815 18575 9873 18581
rect 10229 18581 10241 18584
rect 10275 18612 10287 18615
rect 10318 18612 10324 18624
rect 10275 18584 10324 18612
rect 10275 18581 10287 18584
rect 10229 18575 10287 18581
rect 10318 18572 10324 18584
rect 10376 18572 10382 18624
rect 10870 18572 10876 18624
rect 10928 18612 10934 18624
rect 11655 18615 11713 18621
rect 11655 18612 11667 18615
rect 10928 18584 11667 18612
rect 10928 18572 10934 18584
rect 11655 18581 11667 18584
rect 11701 18581 11713 18615
rect 11655 18575 11713 18581
rect 12805 18615 12863 18621
rect 12805 18581 12817 18615
rect 12851 18612 12863 18615
rect 14458 18612 14464 18624
rect 12851 18584 14464 18612
rect 12851 18581 12863 18584
rect 12805 18575 12863 18581
rect 14458 18572 14464 18584
rect 14516 18572 14522 18624
rect 14550 18572 14556 18624
rect 14608 18612 14614 18624
rect 14645 18615 14703 18621
rect 14645 18612 14657 18615
rect 14608 18584 14657 18612
rect 14608 18572 14614 18584
rect 14645 18581 14657 18584
rect 14691 18581 14703 18615
rect 14645 18575 14703 18581
rect 15654 18572 15660 18624
rect 15712 18612 15718 18624
rect 15749 18615 15807 18621
rect 15749 18612 15761 18615
rect 15712 18584 15761 18612
rect 15712 18572 15718 18584
rect 15749 18581 15761 18584
rect 15795 18581 15807 18615
rect 15749 18575 15807 18581
rect 19935 18615 19993 18621
rect 19935 18581 19947 18615
rect 19981 18612 19993 18615
rect 20162 18612 20168 18624
rect 19981 18584 20168 18612
rect 19981 18581 19993 18584
rect 19935 18575 19993 18581
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2225 18411 2283 18417
rect 2225 18377 2237 18411
rect 2271 18408 2283 18411
rect 2498 18408 2504 18420
rect 2271 18380 2504 18408
rect 2271 18377 2283 18380
rect 2225 18371 2283 18377
rect 2498 18368 2504 18380
rect 2556 18368 2562 18420
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 5261 18411 5319 18417
rect 5261 18408 5273 18411
rect 4212 18380 5273 18408
rect 4212 18368 4218 18380
rect 5261 18377 5273 18380
rect 5307 18377 5319 18411
rect 5261 18371 5319 18377
rect 6086 18368 6092 18420
rect 6144 18408 6150 18420
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 6144 18380 6561 18408
rect 6144 18368 6150 18380
rect 6549 18377 6561 18380
rect 6595 18377 6607 18411
rect 6549 18371 6607 18377
rect 8018 18368 8024 18420
rect 8076 18408 8082 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 8076 18380 8309 18408
rect 8076 18368 8082 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 9674 18408 9680 18420
rect 9635 18380 9680 18408
rect 8297 18371 8355 18377
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 16390 18368 16396 18420
rect 16448 18408 16454 18420
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 16448 18380 16681 18408
rect 16448 18368 16454 18380
rect 16669 18377 16681 18380
rect 16715 18408 16727 18411
rect 16945 18411 17003 18417
rect 16945 18408 16957 18411
rect 16715 18380 16957 18408
rect 16715 18377 16727 18380
rect 16669 18371 16727 18377
rect 16945 18377 16957 18380
rect 16991 18377 17003 18411
rect 16945 18371 17003 18377
rect 17497 18411 17555 18417
rect 17497 18377 17509 18411
rect 17543 18408 17555 18411
rect 17862 18408 17868 18420
rect 17543 18380 17868 18408
rect 17543 18377 17555 18380
rect 17497 18371 17555 18377
rect 3418 18340 3424 18352
rect 3331 18312 3424 18340
rect 3418 18300 3424 18312
rect 3476 18340 3482 18352
rect 4890 18340 4896 18352
rect 3476 18312 4752 18340
rect 4851 18312 4896 18340
rect 3476 18300 3482 18312
rect 2406 18272 2412 18284
rect 2367 18244 2412 18272
rect 2406 18232 2412 18244
rect 2464 18232 2470 18284
rect 3050 18272 3056 18284
rect 3011 18244 3056 18272
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 4724 18272 4752 18312
rect 4890 18300 4896 18312
rect 4948 18300 4954 18352
rect 6454 18300 6460 18352
rect 6512 18340 6518 18352
rect 7834 18340 7840 18352
rect 6512 18312 7840 18340
rect 6512 18300 6518 18312
rect 7834 18300 7840 18312
rect 7892 18300 7898 18352
rect 16960 18340 16988 18371
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 17954 18368 17960 18420
rect 18012 18408 18018 18420
rect 20993 18411 21051 18417
rect 20993 18408 21005 18411
rect 18012 18380 21005 18408
rect 18012 18368 18018 18380
rect 20993 18377 21005 18380
rect 21039 18408 21051 18411
rect 21082 18408 21088 18420
rect 21039 18380 21088 18408
rect 21039 18377 21051 18380
rect 20993 18371 21051 18377
rect 21082 18368 21088 18380
rect 21140 18408 21146 18420
rect 22738 18408 22744 18420
rect 21140 18380 22744 18408
rect 21140 18368 21146 18380
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 24765 18411 24823 18417
rect 24765 18377 24777 18411
rect 24811 18408 24823 18411
rect 24854 18408 24860 18420
rect 24811 18380 24860 18408
rect 24811 18377 24823 18380
rect 24765 18371 24823 18377
rect 24854 18368 24860 18380
rect 24912 18368 24918 18420
rect 20438 18340 20444 18352
rect 16960 18312 20444 18340
rect 20438 18300 20444 18312
rect 20496 18300 20502 18352
rect 20806 18300 20812 18352
rect 20864 18340 20870 18352
rect 22097 18343 22155 18349
rect 22097 18340 22109 18343
rect 20864 18312 22109 18340
rect 20864 18300 20870 18312
rect 22097 18309 22109 18312
rect 22143 18309 22155 18343
rect 22097 18303 22155 18309
rect 10318 18272 10324 18284
rect 3160 18244 4660 18272
rect 4724 18244 9444 18272
rect 10279 18244 10324 18272
rect 1854 18136 1860 18148
rect 1767 18108 1860 18136
rect 1854 18096 1860 18108
rect 1912 18136 1918 18148
rect 2501 18139 2559 18145
rect 2501 18136 2513 18139
rect 1912 18108 2513 18136
rect 1912 18096 1918 18108
rect 2501 18105 2513 18108
rect 2547 18136 2559 18139
rect 3160 18136 3188 18244
rect 4632 18204 4660 18244
rect 5772 18207 5830 18213
rect 4632 18176 5672 18204
rect 3970 18136 3976 18148
rect 2547 18108 3188 18136
rect 3931 18108 3976 18136
rect 2547 18105 2559 18108
rect 2501 18099 2559 18105
rect 3970 18096 3976 18108
rect 4028 18096 4034 18148
rect 4062 18096 4068 18148
rect 4120 18136 4126 18148
rect 4614 18136 4620 18148
rect 4120 18108 4165 18136
rect 4575 18108 4620 18136
rect 4120 18096 4126 18108
rect 4614 18096 4620 18108
rect 4672 18096 4678 18148
rect 3789 18071 3847 18077
rect 3789 18037 3801 18071
rect 3835 18068 3847 18071
rect 3878 18068 3884 18080
rect 3835 18040 3884 18068
rect 3835 18037 3847 18040
rect 3789 18031 3847 18037
rect 3878 18028 3884 18040
rect 3936 18028 3942 18080
rect 5644 18068 5672 18176
rect 5772 18173 5784 18207
rect 5818 18204 5830 18207
rect 5994 18204 6000 18216
rect 5818 18176 6000 18204
rect 5818 18173 5830 18176
rect 5772 18167 5830 18173
rect 5994 18164 6000 18176
rect 6052 18204 6058 18216
rect 6270 18204 6276 18216
rect 6052 18176 6276 18204
rect 6052 18164 6058 18176
rect 6270 18164 6276 18176
rect 6328 18164 6334 18216
rect 8294 18164 8300 18216
rect 8352 18204 8358 18216
rect 9416 18213 9444 18244
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 10686 18272 10692 18284
rect 10647 18244 10692 18272
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 12342 18232 12348 18284
rect 12400 18272 12406 18284
rect 12529 18275 12587 18281
rect 12529 18272 12541 18275
rect 12400 18244 12541 18272
rect 12400 18232 12406 18244
rect 12529 18241 12541 18244
rect 12575 18241 12587 18275
rect 15838 18272 15844 18284
rect 12529 18235 12587 18241
rect 14752 18244 15844 18272
rect 8481 18207 8539 18213
rect 8481 18204 8493 18207
rect 8352 18176 8493 18204
rect 8352 18164 8358 18176
rect 8481 18173 8493 18176
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 9401 18207 9459 18213
rect 9401 18173 9413 18207
rect 9447 18204 9459 18207
rect 10045 18207 10103 18213
rect 10045 18204 10057 18207
rect 9447 18176 10057 18204
rect 9447 18173 9459 18176
rect 9401 18167 9459 18173
rect 10045 18173 10057 18176
rect 10091 18173 10103 18207
rect 10045 18167 10103 18173
rect 5859 18139 5917 18145
rect 5859 18105 5871 18139
rect 5905 18136 5917 18139
rect 6914 18136 6920 18148
rect 5905 18108 6920 18136
rect 5905 18105 5917 18108
rect 5859 18099 5917 18105
rect 6914 18096 6920 18108
rect 6972 18096 6978 18148
rect 7009 18139 7067 18145
rect 7009 18105 7021 18139
rect 7055 18105 7067 18139
rect 7558 18136 7564 18148
rect 7519 18108 7564 18136
rect 7009 18099 7067 18105
rect 7024 18068 7052 18099
rect 7558 18096 7564 18108
rect 7616 18096 7622 18148
rect 8802 18139 8860 18145
rect 8802 18105 8814 18139
rect 8848 18105 8860 18139
rect 10060 18136 10088 18167
rect 11606 18164 11612 18216
rect 11664 18204 11670 18216
rect 12158 18204 12164 18216
rect 11664 18176 12164 18204
rect 11664 18164 11670 18176
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 13262 18164 13268 18216
rect 13320 18204 13326 18216
rect 14093 18207 14151 18213
rect 14093 18204 14105 18207
rect 13320 18176 14105 18204
rect 13320 18164 13326 18176
rect 14093 18173 14105 18176
rect 14139 18204 14151 18207
rect 14366 18204 14372 18216
rect 14139 18176 14372 18204
rect 14139 18173 14151 18176
rect 14093 18167 14151 18173
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 14458 18164 14464 18216
rect 14516 18204 14522 18216
rect 14752 18213 14780 18244
rect 15838 18232 15844 18244
rect 15896 18272 15902 18284
rect 17034 18272 17040 18284
rect 15896 18244 17040 18272
rect 15896 18232 15902 18244
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 18414 18272 18420 18284
rect 18375 18244 18420 18272
rect 18414 18232 18420 18244
rect 18472 18272 18478 18284
rect 19337 18275 19395 18281
rect 19337 18272 19349 18275
rect 18472 18244 19349 18272
rect 18472 18232 18478 18244
rect 19337 18241 19349 18244
rect 19383 18241 19395 18275
rect 21450 18272 21456 18284
rect 19337 18235 19395 18241
rect 20916 18244 21456 18272
rect 14737 18207 14795 18213
rect 14737 18204 14749 18207
rect 14516 18176 14749 18204
rect 14516 18164 14522 18176
rect 14737 18173 14749 18176
rect 14783 18173 14795 18207
rect 14737 18167 14795 18173
rect 15654 18164 15660 18216
rect 15712 18204 15718 18216
rect 15749 18207 15807 18213
rect 15749 18204 15761 18207
rect 15712 18176 15761 18204
rect 15712 18164 15718 18176
rect 15749 18173 15761 18176
rect 15795 18173 15807 18207
rect 15749 18167 15807 18173
rect 19061 18207 19119 18213
rect 19061 18173 19073 18207
rect 19107 18204 19119 18207
rect 20916 18204 20944 18244
rect 21450 18232 21456 18244
rect 21508 18272 21514 18284
rect 23106 18272 23112 18284
rect 21508 18244 23112 18272
rect 21508 18232 21514 18244
rect 23106 18232 23112 18244
rect 23164 18232 23170 18284
rect 19107 18176 20944 18204
rect 19107 18173 19119 18176
rect 19061 18167 19119 18173
rect 23566 18164 23572 18216
rect 23624 18204 23630 18216
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 23624 18176 24593 18204
rect 23624 18164 23630 18176
rect 24581 18173 24593 18176
rect 24627 18204 24639 18207
rect 25133 18207 25191 18213
rect 25133 18204 25145 18207
rect 24627 18176 25145 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 25133 18173 25145 18176
rect 25179 18173 25191 18207
rect 25133 18167 25191 18173
rect 10413 18139 10471 18145
rect 10413 18136 10425 18139
rect 10060 18108 10425 18136
rect 8802 18099 8860 18105
rect 10413 18105 10425 18108
rect 10459 18105 10471 18139
rect 10413 18099 10471 18105
rect 7098 18068 7104 18080
rect 5644 18040 7104 18068
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 7926 18068 7932 18080
rect 7887 18040 7932 18068
rect 7926 18028 7932 18040
rect 7984 18068 7990 18080
rect 8817 18068 8845 18099
rect 12526 18096 12532 18148
rect 12584 18136 12590 18148
rect 12621 18139 12679 18145
rect 12621 18136 12633 18139
rect 12584 18108 12633 18136
rect 12584 18096 12590 18108
rect 12621 18105 12633 18108
rect 12667 18105 12679 18139
rect 12621 18099 12679 18105
rect 13173 18139 13231 18145
rect 13173 18105 13185 18139
rect 13219 18136 13231 18139
rect 13354 18136 13360 18148
rect 13219 18108 13360 18136
rect 13219 18105 13231 18108
rect 13173 18099 13231 18105
rect 13354 18096 13360 18108
rect 13412 18096 13418 18148
rect 13725 18139 13783 18145
rect 13725 18105 13737 18139
rect 13771 18136 13783 18139
rect 14550 18136 14556 18148
rect 13771 18108 14556 18136
rect 13771 18105 13783 18108
rect 13725 18099 13783 18105
rect 14550 18096 14556 18108
rect 14608 18096 14614 18148
rect 14921 18139 14979 18145
rect 14921 18105 14933 18139
rect 14967 18136 14979 18139
rect 15470 18136 15476 18148
rect 14967 18108 15476 18136
rect 14967 18105 14979 18108
rect 14921 18099 14979 18105
rect 15470 18096 15476 18108
rect 15528 18096 15534 18148
rect 16070 18139 16128 18145
rect 16070 18136 16082 18139
rect 15580 18108 16082 18136
rect 15580 18080 15608 18108
rect 16070 18105 16082 18108
rect 16116 18105 16128 18139
rect 16070 18099 16128 18105
rect 18506 18096 18512 18148
rect 18564 18136 18570 18148
rect 19886 18136 19892 18148
rect 18564 18108 18609 18136
rect 19799 18108 19892 18136
rect 18564 18096 18570 18108
rect 19886 18096 19892 18108
rect 19944 18136 19950 18148
rect 20346 18136 20352 18148
rect 19944 18108 20352 18136
rect 19944 18096 19950 18108
rect 20346 18096 20352 18108
rect 20404 18096 20410 18148
rect 21174 18136 21180 18148
rect 21135 18108 21180 18136
rect 21174 18096 21180 18108
rect 21232 18096 21238 18148
rect 21269 18139 21327 18145
rect 21269 18105 21281 18139
rect 21315 18105 21327 18139
rect 21269 18099 21327 18105
rect 7984 18040 8845 18068
rect 11609 18071 11667 18077
rect 7984 18028 7990 18040
rect 11609 18037 11621 18071
rect 11655 18068 11667 18071
rect 11698 18068 11704 18080
rect 11655 18040 11704 18068
rect 11655 18037 11667 18040
rect 11609 18031 11667 18037
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 15562 18068 15568 18080
rect 15523 18040 15568 18068
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 17218 18028 17224 18080
rect 17276 18068 17282 18080
rect 17773 18071 17831 18077
rect 17773 18068 17785 18071
rect 17276 18040 17785 18068
rect 17276 18028 17282 18040
rect 17773 18037 17785 18040
rect 17819 18068 17831 18071
rect 18046 18068 18052 18080
rect 17819 18040 18052 18068
rect 17819 18037 17831 18040
rect 17773 18031 17831 18037
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 20070 18068 20076 18080
rect 20031 18040 20076 18068
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 20530 18068 20536 18080
rect 20491 18040 20536 18068
rect 20530 18028 20536 18040
rect 20588 18068 20594 18080
rect 21284 18068 21312 18099
rect 20588 18040 21312 18068
rect 20588 18028 20594 18040
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2406 17824 2412 17876
rect 2464 17864 2470 17876
rect 2961 17867 3019 17873
rect 2961 17864 2973 17867
rect 2464 17836 2973 17864
rect 2464 17824 2470 17836
rect 2961 17833 2973 17836
rect 3007 17833 3019 17867
rect 2961 17827 3019 17833
rect 3878 17824 3884 17876
rect 3936 17864 3942 17876
rect 4062 17864 4068 17876
rect 3936 17836 4068 17864
rect 3936 17824 3942 17836
rect 4062 17824 4068 17836
rect 4120 17864 4126 17876
rect 5169 17867 5227 17873
rect 5169 17864 5181 17867
rect 4120 17836 5181 17864
rect 4120 17824 4126 17836
rect 5169 17833 5181 17836
rect 5215 17833 5227 17867
rect 6454 17864 6460 17876
rect 6415 17836 6460 17864
rect 5169 17827 5227 17833
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 6972 17836 7665 17864
rect 6972 17824 6978 17836
rect 7653 17833 7665 17836
rect 7699 17833 7711 17867
rect 9766 17864 9772 17876
rect 9727 17836 9772 17864
rect 7653 17827 7711 17833
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 10870 17864 10876 17876
rect 10831 17836 10876 17864
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 14458 17864 14464 17876
rect 14419 17836 14464 17864
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 16298 17824 16304 17876
rect 16356 17864 16362 17876
rect 16577 17867 16635 17873
rect 16577 17864 16589 17867
rect 16356 17836 16589 17864
rect 16356 17824 16362 17836
rect 16577 17833 16589 17836
rect 16623 17833 16635 17867
rect 17678 17864 17684 17876
rect 17639 17836 17684 17864
rect 16577 17827 16635 17833
rect 17678 17824 17684 17836
rect 17736 17824 17742 17876
rect 18233 17867 18291 17873
rect 18233 17833 18245 17867
rect 18279 17864 18291 17867
rect 18506 17864 18512 17876
rect 18279 17836 18512 17864
rect 18279 17833 18291 17836
rect 18233 17827 18291 17833
rect 18506 17824 18512 17836
rect 18564 17824 18570 17876
rect 18966 17864 18972 17876
rect 18927 17836 18972 17864
rect 18966 17824 18972 17836
rect 19024 17864 19030 17876
rect 19426 17864 19432 17876
rect 19024 17836 19104 17864
rect 19387 17836 19432 17864
rect 19024 17824 19030 17836
rect 2038 17756 2044 17808
rect 2096 17796 2102 17808
rect 2133 17799 2191 17805
rect 2133 17796 2145 17799
rect 2096 17768 2145 17796
rect 2096 17756 2102 17768
rect 2133 17765 2145 17768
rect 2179 17796 2191 17799
rect 2179 17768 2728 17796
rect 2179 17765 2191 17768
rect 2133 17759 2191 17765
rect 2700 17728 2728 17768
rect 4154 17756 4160 17808
rect 4212 17796 4218 17808
rect 4570 17799 4628 17805
rect 4570 17796 4582 17799
rect 4212 17768 4582 17796
rect 4212 17756 4218 17768
rect 4570 17765 4582 17768
rect 4616 17765 4628 17799
rect 4570 17759 4628 17765
rect 7098 17756 7104 17808
rect 7156 17796 7162 17808
rect 7285 17799 7343 17805
rect 7285 17796 7297 17799
rect 7156 17768 7297 17796
rect 7156 17756 7162 17768
rect 7285 17765 7297 17768
rect 7331 17765 7343 17799
rect 8202 17796 8208 17808
rect 8163 17768 8208 17796
rect 7285 17759 7343 17765
rect 8202 17756 8208 17768
rect 8260 17756 8266 17808
rect 10042 17796 10048 17808
rect 9784 17768 10048 17796
rect 6546 17728 6552 17740
rect 2700 17700 6552 17728
rect 6546 17688 6552 17700
rect 6604 17728 6610 17740
rect 9784 17737 9812 17768
rect 10042 17756 10048 17768
rect 10100 17756 10106 17808
rect 11603 17799 11661 17805
rect 11603 17765 11615 17799
rect 11649 17796 11661 17799
rect 11882 17796 11888 17808
rect 11649 17768 11888 17796
rect 11649 17765 11661 17768
rect 11603 17759 11661 17765
rect 11882 17756 11888 17768
rect 11940 17756 11946 17808
rect 13170 17796 13176 17808
rect 13131 17768 13176 17796
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 15562 17756 15568 17808
rect 15620 17796 15626 17808
rect 15743 17799 15801 17805
rect 15743 17796 15755 17799
rect 15620 17768 15755 17796
rect 15620 17756 15626 17768
rect 15743 17765 15755 17768
rect 15789 17796 15801 17799
rect 17696 17796 17724 17824
rect 15789 17768 17724 17796
rect 15789 17765 15801 17768
rect 15743 17759 15801 17765
rect 7009 17731 7067 17737
rect 7009 17728 7021 17731
rect 6604 17700 7021 17728
rect 6604 17688 6610 17700
rect 7009 17697 7021 17700
rect 7055 17697 7067 17731
rect 7009 17691 7067 17697
rect 9769 17731 9827 17737
rect 9769 17697 9781 17731
rect 9815 17697 9827 17731
rect 9769 17691 9827 17697
rect 9858 17688 9864 17740
rect 9916 17728 9922 17740
rect 10137 17731 10195 17737
rect 10137 17728 10149 17731
rect 9916 17700 10149 17728
rect 9916 17688 9922 17700
rect 10137 17697 10149 17700
rect 10183 17697 10195 17731
rect 10137 17691 10195 17697
rect 16301 17731 16359 17737
rect 16301 17697 16313 17731
rect 16347 17728 16359 17731
rect 17218 17728 17224 17740
rect 16347 17700 17224 17728
rect 16347 17697 16359 17700
rect 16301 17691 16359 17697
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 17313 17731 17371 17737
rect 17313 17697 17325 17731
rect 17359 17728 17371 17731
rect 18138 17728 18144 17740
rect 17359 17700 18144 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 18138 17688 18144 17700
rect 18196 17688 18202 17740
rect 19076 17737 19104 17836
rect 19426 17824 19432 17836
rect 19484 17824 19490 17876
rect 21174 17824 21180 17876
rect 21232 17864 21238 17876
rect 21913 17867 21971 17873
rect 21913 17864 21925 17867
rect 21232 17836 21925 17864
rect 21232 17824 21238 17836
rect 21913 17833 21925 17836
rect 21959 17864 21971 17867
rect 24762 17864 24768 17876
rect 21959 17836 23244 17864
rect 24723 17836 24768 17864
rect 21959 17833 21971 17836
rect 21913 17827 21971 17833
rect 23216 17808 23244 17836
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 21082 17796 21088 17808
rect 19996 17768 21088 17796
rect 19996 17737 20024 17768
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 22370 17756 22376 17808
rect 22428 17796 22434 17808
rect 22649 17799 22707 17805
rect 22649 17796 22661 17799
rect 22428 17768 22661 17796
rect 22428 17756 22434 17768
rect 22649 17765 22661 17768
rect 22695 17765 22707 17799
rect 23198 17796 23204 17808
rect 23111 17768 23204 17796
rect 22649 17759 22707 17765
rect 23198 17756 23204 17768
rect 23256 17756 23262 17808
rect 19061 17731 19119 17737
rect 19061 17697 19073 17731
rect 19107 17697 19119 17731
rect 19061 17691 19119 17697
rect 19981 17731 20039 17737
rect 19981 17697 19993 17731
rect 20027 17697 20039 17731
rect 19981 17691 20039 17697
rect 24118 17688 24124 17740
rect 24176 17728 24182 17740
rect 24581 17731 24639 17737
rect 24581 17728 24593 17731
rect 24176 17700 24593 17728
rect 24176 17688 24182 17700
rect 24581 17697 24593 17700
rect 24627 17697 24639 17731
rect 24581 17691 24639 17697
rect 1857 17663 1915 17669
rect 1857 17629 1869 17663
rect 1903 17660 1915 17663
rect 2041 17663 2099 17669
rect 2041 17660 2053 17663
rect 1903 17632 2053 17660
rect 1903 17629 1915 17632
rect 1857 17623 1915 17629
rect 2041 17629 2053 17632
rect 2087 17660 2099 17663
rect 3142 17660 3148 17672
rect 2087 17632 3148 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 3142 17620 3148 17632
rect 3200 17620 3206 17672
rect 3418 17620 3424 17672
rect 3476 17660 3482 17672
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 3476 17632 4261 17660
rect 3476 17620 3482 17632
rect 4249 17629 4261 17632
rect 4295 17660 4307 17663
rect 5166 17660 5172 17672
rect 4295 17632 5172 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 5994 17620 6000 17672
rect 6052 17660 6058 17672
rect 6089 17663 6147 17669
rect 6089 17660 6101 17663
rect 6052 17632 6101 17660
rect 6052 17620 6058 17632
rect 6089 17629 6101 17632
rect 6135 17629 6147 17663
rect 6089 17623 6147 17629
rect 7558 17620 7564 17672
rect 7616 17660 7622 17672
rect 8113 17663 8171 17669
rect 8113 17660 8125 17663
rect 7616 17632 8125 17660
rect 7616 17620 7622 17632
rect 8113 17629 8125 17632
rect 8159 17660 8171 17663
rect 10686 17660 10692 17672
rect 8159 17632 10692 17660
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 10686 17620 10692 17632
rect 10744 17620 10750 17672
rect 11238 17660 11244 17672
rect 11199 17632 11244 17660
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13354 17660 13360 17672
rect 13127 17632 13360 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 13722 17660 13728 17672
rect 13683 17632 13728 17660
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 15378 17660 15384 17672
rect 15339 17632 15384 17660
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 20993 17663 21051 17669
rect 20993 17629 21005 17663
rect 21039 17660 21051 17663
rect 21266 17660 21272 17672
rect 21039 17632 21272 17660
rect 21039 17629 21051 17632
rect 20993 17623 21051 17629
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 21450 17660 21456 17672
rect 21411 17632 21456 17660
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 22554 17660 22560 17672
rect 22515 17632 22560 17660
rect 22554 17620 22560 17632
rect 22612 17620 22618 17672
rect 2590 17592 2596 17604
rect 2551 17564 2596 17592
rect 2590 17552 2596 17564
rect 2648 17592 2654 17604
rect 3789 17595 3847 17601
rect 3789 17592 3801 17595
rect 2648 17564 3801 17592
rect 2648 17552 2654 17564
rect 3789 17561 3801 17564
rect 3835 17592 3847 17595
rect 3970 17592 3976 17604
rect 3835 17564 3976 17592
rect 3835 17561 3847 17564
rect 3789 17555 3847 17561
rect 3970 17552 3976 17564
rect 4028 17552 4034 17604
rect 4614 17552 4620 17604
rect 4672 17592 4678 17604
rect 8665 17595 8723 17601
rect 8665 17592 8677 17595
rect 4672 17564 8677 17592
rect 4672 17552 4678 17564
rect 8665 17561 8677 17564
rect 8711 17561 8723 17595
rect 8665 17555 8723 17561
rect 11054 17552 11060 17604
rect 11112 17592 11118 17604
rect 13814 17592 13820 17604
rect 11112 17564 13820 17592
rect 11112 17552 11118 17564
rect 13786 17552 13820 17564
rect 13872 17552 13878 17604
rect 20622 17552 20628 17604
rect 20680 17592 20686 17604
rect 23474 17592 23480 17604
rect 20680 17564 23480 17592
rect 20680 17552 20686 17564
rect 23474 17552 23480 17564
rect 23532 17552 23538 17604
rect 11330 17484 11336 17536
rect 11388 17524 11394 17536
rect 12161 17527 12219 17533
rect 12161 17524 12173 17527
rect 11388 17496 12173 17524
rect 11388 17484 11394 17496
rect 12161 17493 12173 17496
rect 12207 17524 12219 17527
rect 12437 17527 12495 17533
rect 12437 17524 12449 17527
rect 12207 17496 12449 17524
rect 12207 17493 12219 17496
rect 12161 17487 12219 17493
rect 12437 17493 12449 17496
rect 12483 17524 12495 17527
rect 12526 17524 12532 17536
rect 12483 17496 12532 17524
rect 12483 17493 12495 17496
rect 12437 17487 12495 17493
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 12805 17527 12863 17533
rect 12805 17524 12817 17527
rect 12676 17496 12817 17524
rect 12676 17484 12682 17496
rect 12805 17493 12817 17496
rect 12851 17493 12863 17527
rect 13786 17524 13814 17552
rect 14093 17527 14151 17533
rect 14093 17524 14105 17527
rect 13786 17496 14105 17524
rect 12805 17487 12863 17493
rect 14093 17493 14105 17496
rect 14139 17524 14151 17527
rect 15562 17524 15568 17536
rect 14139 17496 15568 17524
rect 14139 17493 14151 17496
rect 14093 17487 14151 17493
rect 15562 17484 15568 17496
rect 15620 17484 15626 17536
rect 18046 17484 18052 17536
rect 18104 17524 18110 17536
rect 20898 17524 20904 17536
rect 18104 17496 20904 17524
rect 18104 17484 18110 17496
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 2038 17320 2044 17332
rect 1719 17292 2044 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 2038 17280 2044 17292
rect 2096 17280 2102 17332
rect 3418 17320 3424 17332
rect 3379 17292 3424 17320
rect 3418 17280 3424 17292
rect 3476 17280 3482 17332
rect 4890 17280 4896 17332
rect 4948 17320 4954 17332
rect 5169 17323 5227 17329
rect 5169 17320 5181 17323
rect 4948 17292 5181 17320
rect 4948 17280 4954 17292
rect 5169 17289 5181 17292
rect 5215 17289 5227 17323
rect 5169 17283 5227 17289
rect 7098 17280 7104 17332
rect 7156 17320 7162 17332
rect 7745 17323 7803 17329
rect 7745 17320 7757 17323
rect 7156 17292 7757 17320
rect 7156 17280 7162 17292
rect 7745 17289 7757 17292
rect 7791 17289 7803 17323
rect 7745 17283 7803 17289
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 10137 17323 10195 17329
rect 10137 17320 10149 17323
rect 9916 17292 10149 17320
rect 9916 17280 9922 17292
rect 10137 17289 10149 17292
rect 10183 17289 10195 17323
rect 10137 17283 10195 17289
rect 13170 17280 13176 17332
rect 13228 17320 13234 17332
rect 13357 17323 13415 17329
rect 13357 17320 13369 17323
rect 13228 17292 13369 17320
rect 13228 17280 13234 17292
rect 13357 17289 13369 17292
rect 13403 17320 13415 17323
rect 13633 17323 13691 17329
rect 13633 17320 13645 17323
rect 13403 17292 13645 17320
rect 13403 17289 13415 17292
rect 13357 17283 13415 17289
rect 13633 17289 13645 17292
rect 13679 17289 13691 17323
rect 13633 17283 13691 17289
rect 16393 17323 16451 17329
rect 16393 17289 16405 17323
rect 16439 17320 16451 17323
rect 16482 17320 16488 17332
rect 16439 17292 16488 17320
rect 16439 17289 16451 17292
rect 16393 17283 16451 17289
rect 16482 17280 16488 17292
rect 16540 17320 16546 17332
rect 17773 17323 17831 17329
rect 16540 17292 17356 17320
rect 16540 17280 16546 17292
rect 8113 17255 8171 17261
rect 8113 17221 8125 17255
rect 8159 17252 8171 17255
rect 8202 17252 8208 17264
rect 8159 17224 8208 17252
rect 8159 17221 8171 17224
rect 8113 17215 8171 17221
rect 8202 17212 8208 17224
rect 8260 17252 8266 17264
rect 9493 17255 9551 17261
rect 9493 17252 9505 17255
rect 8260 17224 9505 17252
rect 8260 17212 8266 17224
rect 9493 17221 9505 17224
rect 9539 17221 9551 17255
rect 9493 17215 9551 17221
rect 10013 17224 11008 17252
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17184 2467 17187
rect 2866 17184 2872 17196
rect 2455 17156 2872 17184
rect 2455 17153 2467 17156
rect 2409 17147 2467 17153
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 3050 17184 3056 17196
rect 3011 17156 3056 17184
rect 3050 17144 3056 17156
rect 3108 17144 3114 17196
rect 6089 17187 6147 17193
rect 6089 17184 6101 17187
rect 4515 17156 6101 17184
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17116 3847 17119
rect 4246 17116 4252 17128
rect 3835 17088 4252 17116
rect 3835 17085 3847 17088
rect 3789 17079 3847 17085
rect 4246 17076 4252 17088
rect 4304 17076 4310 17128
rect 4515 17057 4543 17156
rect 6089 17153 6101 17156
rect 6135 17184 6147 17187
rect 6454 17184 6460 17196
rect 6135 17156 6460 17184
rect 6135 17153 6147 17156
rect 6089 17147 6147 17153
rect 6454 17144 6460 17156
rect 6512 17184 6518 17196
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 6512 17156 6561 17184
rect 6512 17144 6518 17156
rect 6549 17153 6561 17156
rect 6595 17184 6607 17187
rect 6595 17156 7052 17184
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 6822 17116 6828 17128
rect 6783 17088 6828 17116
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 2501 17051 2559 17057
rect 2501 17017 2513 17051
rect 2547 17017 2559 17051
rect 2501 17011 2559 17017
rect 4500 17051 4558 17057
rect 4500 17017 4512 17051
rect 4546 17017 4558 17051
rect 4500 17011 4558 17017
rect 5813 17051 5871 17057
rect 5813 17017 5825 17051
rect 5859 17048 5871 17051
rect 5994 17048 6000 17060
rect 5859 17020 6000 17048
rect 5859 17017 5871 17020
rect 5813 17011 5871 17017
rect 2038 16940 2044 16992
rect 2096 16980 2102 16992
rect 2516 16980 2544 17011
rect 4154 16980 4160 16992
rect 2096 16952 2544 16980
rect 4115 16952 4160 16980
rect 2096 16940 2102 16952
rect 4154 16940 4160 16952
rect 4212 16980 4218 16992
rect 4515 16980 4543 17011
rect 5994 17008 6000 17020
rect 6052 17048 6058 17060
rect 6914 17048 6920 17060
rect 6052 17020 6920 17048
rect 6052 17008 6058 17020
rect 6914 17008 6920 17020
rect 6972 17008 6978 17060
rect 7024 17048 7052 17156
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 10013 17184 10041 17224
rect 10870 17184 10876 17196
rect 7708 17156 10041 17184
rect 10831 17156 10876 17184
rect 7708 17144 7714 17156
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 10980 17184 11008 17224
rect 13446 17212 13452 17264
rect 13504 17252 13510 17264
rect 14323 17255 14381 17261
rect 14323 17252 14335 17255
rect 13504 17224 14335 17252
rect 13504 17212 13510 17224
rect 14323 17221 14335 17224
rect 14369 17221 14381 17255
rect 17328 17252 17356 17292
rect 17773 17289 17785 17323
rect 17819 17320 17831 17323
rect 18138 17320 18144 17332
rect 17819 17292 18144 17320
rect 17819 17289 17831 17292
rect 17773 17283 17831 17289
rect 18138 17280 18144 17292
rect 18196 17280 18202 17332
rect 20070 17280 20076 17332
rect 20128 17320 20134 17332
rect 20809 17323 20867 17329
rect 20809 17320 20821 17323
rect 20128 17292 20821 17320
rect 20128 17280 20134 17292
rect 20809 17289 20821 17292
rect 20855 17289 20867 17323
rect 20809 17283 20867 17289
rect 17954 17252 17960 17264
rect 14323 17215 14381 17221
rect 15304 17224 16804 17252
rect 17328 17224 17960 17252
rect 15304 17184 15332 17224
rect 10980 17156 15332 17184
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15436 17156 16681 17184
rect 15436 17144 15442 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 9766 17116 9772 17128
rect 8619 17088 9772 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12032 17088 12449 17116
rect 12032 17076 12038 17088
rect 12437 17085 12449 17088
rect 12483 17116 12495 17119
rect 12618 17116 12624 17128
rect 12483 17088 12624 17116
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 15470 17116 15476 17128
rect 13786 17088 14136 17116
rect 15431 17088 15476 17116
rect 7146 17051 7204 17057
rect 7146 17048 7158 17051
rect 7024 17020 7158 17048
rect 7146 17017 7158 17020
rect 7192 17048 7204 17051
rect 7926 17048 7932 17060
rect 7192 17020 7932 17048
rect 7192 17017 7204 17020
rect 7146 17011 7204 17017
rect 7926 17008 7932 17020
rect 7984 17048 7990 17060
rect 8389 17051 8447 17057
rect 8389 17048 8401 17051
rect 7984 17020 8401 17048
rect 7984 17008 7990 17020
rect 8389 17017 8401 17020
rect 8435 17048 8447 17051
rect 8894 17051 8952 17057
rect 8894 17048 8906 17051
rect 8435 17020 8906 17048
rect 8435 17017 8447 17020
rect 8389 17011 8447 17017
rect 8894 17017 8906 17020
rect 8940 17048 8952 17051
rect 10689 17051 10747 17057
rect 8940 17020 10640 17048
rect 8940 17017 8952 17020
rect 8894 17011 8952 17017
rect 4212 16952 4543 16980
rect 9861 16983 9919 16989
rect 4212 16940 4218 16952
rect 9861 16949 9873 16983
rect 9907 16980 9919 16983
rect 10042 16980 10048 16992
rect 9907 16952 10048 16980
rect 9907 16949 9919 16952
rect 9861 16943 9919 16949
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10612 16980 10640 17020
rect 10689 17017 10701 17051
rect 10735 17048 10747 17051
rect 10965 17051 11023 17057
rect 10965 17048 10977 17051
rect 10735 17020 10977 17048
rect 10735 17017 10747 17020
rect 10689 17011 10747 17017
rect 10965 17017 10977 17020
rect 11011 17048 11023 17051
rect 11330 17048 11336 17060
rect 11011 17020 11336 17048
rect 11011 17017 11023 17020
rect 10965 17011 11023 17017
rect 11330 17008 11336 17020
rect 11388 17008 11394 17060
rect 11514 17048 11520 17060
rect 11475 17020 11520 17048
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 11882 17048 11888 17060
rect 11795 17020 11888 17048
rect 11882 17008 11888 17020
rect 11940 17048 11946 17060
rect 12253 17051 12311 17057
rect 12253 17048 12265 17051
rect 11940 17020 12265 17048
rect 11940 17008 11946 17020
rect 12253 17017 12265 17020
rect 12299 17048 12311 17051
rect 12799 17051 12857 17057
rect 12799 17048 12811 17051
rect 12299 17020 12811 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12799 17017 12811 17020
rect 12845 17048 12857 17051
rect 13786 17048 13814 17088
rect 12845 17020 13814 17048
rect 14108 17048 14136 17088
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 16776 17116 16804 17224
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 20165 17255 20223 17261
rect 20165 17221 20177 17255
rect 20211 17252 20223 17255
rect 20530 17252 20536 17264
rect 20211 17224 20536 17252
rect 20211 17221 20223 17224
rect 20165 17215 20223 17221
rect 20530 17212 20536 17224
rect 20588 17212 20594 17264
rect 18782 17144 18788 17196
rect 18840 17184 18846 17196
rect 19245 17187 19303 17193
rect 19245 17184 19257 17187
rect 18840 17156 19257 17184
rect 18840 17144 18846 17156
rect 19245 17153 19257 17156
rect 19291 17184 19303 17187
rect 20070 17184 20076 17196
rect 19291 17156 20076 17184
rect 19291 17153 19303 17156
rect 19245 17147 19303 17153
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 20438 17184 20444 17196
rect 20399 17156 20444 17184
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 20824 17184 20852 17283
rect 21082 17280 21088 17332
rect 21140 17320 21146 17332
rect 22005 17323 22063 17329
rect 22005 17320 22017 17323
rect 21140 17292 22017 17320
rect 21140 17280 21146 17292
rect 22005 17289 22017 17292
rect 22051 17289 22063 17323
rect 23106 17320 23112 17332
rect 23067 17292 23112 17320
rect 22005 17283 22063 17289
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 20898 17212 20904 17264
rect 20956 17252 20962 17264
rect 23385 17255 23443 17261
rect 23385 17252 23397 17255
rect 20956 17224 23397 17252
rect 20956 17212 20962 17224
rect 23385 17221 23397 17224
rect 23431 17252 23443 17255
rect 23842 17252 23848 17264
rect 23431 17224 23848 17252
rect 23431 17221 23443 17224
rect 23385 17215 23443 17221
rect 23842 17212 23848 17224
rect 23900 17212 23906 17264
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 20824 17156 21097 17184
rect 21085 17153 21097 17156
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 21266 17144 21272 17196
rect 21324 17184 21330 17196
rect 21361 17187 21419 17193
rect 21361 17184 21373 17187
rect 21324 17156 21373 17184
rect 21324 17144 21330 17156
rect 21361 17153 21373 17156
rect 21407 17153 21419 17187
rect 21361 17147 21419 17153
rect 23198 17144 23204 17196
rect 23256 17184 23262 17196
rect 24029 17187 24087 17193
rect 24029 17184 24041 17187
rect 23256 17156 24041 17184
rect 23256 17144 23262 17156
rect 24029 17153 24041 17156
rect 24075 17153 24087 17187
rect 24029 17147 24087 17153
rect 18084 17119 18142 17125
rect 18084 17116 18096 17119
rect 16776 17088 18096 17116
rect 18084 17085 18096 17088
rect 18130 17116 18142 17119
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 18130 17088 18521 17116
rect 18130 17085 18142 17088
rect 18084 17079 18142 17085
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 15013 17051 15071 17057
rect 15013 17048 15025 17051
rect 14108 17020 15025 17048
rect 12845 17017 12857 17020
rect 12799 17011 12857 17017
rect 15013 17017 15025 17020
rect 15059 17048 15071 17051
rect 15381 17051 15439 17057
rect 15381 17048 15393 17051
rect 15059 17020 15393 17048
rect 15059 17017 15071 17020
rect 15013 17011 15071 17017
rect 15381 17017 15393 17020
rect 15427 17048 15439 17051
rect 15835 17051 15893 17057
rect 15835 17048 15847 17051
rect 15427 17020 15847 17048
rect 15427 17017 15439 17020
rect 15381 17011 15439 17017
rect 15835 17017 15847 17020
rect 15881 17048 15893 17051
rect 17405 17051 17463 17057
rect 17405 17048 17417 17051
rect 15881 17020 17417 17048
rect 15881 17017 15893 17020
rect 15835 17011 15893 17017
rect 17405 17017 17417 17020
rect 17451 17048 17463 17051
rect 17678 17048 17684 17060
rect 17451 17020 17684 17048
rect 17451 17017 17463 17020
rect 17405 17011 17463 17017
rect 17678 17008 17684 17020
rect 17736 17048 17742 17060
rect 19426 17048 19432 17060
rect 17736 17020 19432 17048
rect 17736 17008 17742 17020
rect 11900 16980 11928 17008
rect 19076 16992 19104 17020
rect 19426 17008 19432 17020
rect 19484 17048 19490 17060
rect 19566 17051 19624 17057
rect 19566 17048 19578 17051
rect 19484 17020 19578 17048
rect 19484 17008 19490 17020
rect 19566 17017 19578 17020
rect 19612 17017 19624 17051
rect 20456 17048 20484 17144
rect 22624 17119 22682 17125
rect 22624 17085 22636 17119
rect 22670 17116 22682 17119
rect 23106 17116 23112 17128
rect 22670 17088 23112 17116
rect 22670 17085 22682 17088
rect 22624 17079 22682 17085
rect 23106 17076 23112 17088
rect 23164 17076 23170 17128
rect 21177 17051 21235 17057
rect 21177 17048 21189 17051
rect 20456 17020 21189 17048
rect 19566 17011 19624 17017
rect 21177 17017 21189 17020
rect 21223 17048 21235 17051
rect 22370 17048 22376 17060
rect 21223 17020 22376 17048
rect 21223 17017 21235 17020
rect 21177 17011 21235 17017
rect 22370 17008 22376 17020
rect 22428 17008 22434 17060
rect 23750 17048 23756 17060
rect 23711 17020 23756 17048
rect 23750 17008 23756 17020
rect 23808 17008 23814 17060
rect 23842 17008 23848 17060
rect 23900 17048 23906 17060
rect 23900 17020 23945 17048
rect 23900 17008 23906 17020
rect 10612 16952 11928 16980
rect 13446 16940 13452 16992
rect 13504 16980 13510 16992
rect 13722 16980 13728 16992
rect 13504 16952 13728 16980
rect 13504 16940 13510 16952
rect 13722 16940 13728 16952
rect 13780 16980 13786 16992
rect 14001 16983 14059 16989
rect 14001 16980 14013 16983
rect 13780 16952 14013 16980
rect 13780 16940 13786 16952
rect 14001 16949 14013 16952
rect 14047 16949 14059 16983
rect 14001 16943 14059 16949
rect 17770 16940 17776 16992
rect 17828 16980 17834 16992
rect 18187 16983 18245 16989
rect 18187 16980 18199 16983
rect 17828 16952 18199 16980
rect 17828 16940 17834 16952
rect 18187 16949 18199 16952
rect 18233 16949 18245 16983
rect 19058 16980 19064 16992
rect 19019 16952 19064 16980
rect 18187 16943 18245 16949
rect 19058 16940 19064 16952
rect 19116 16940 19122 16992
rect 22554 16940 22560 16992
rect 22612 16980 22618 16992
rect 22695 16983 22753 16989
rect 22695 16980 22707 16983
rect 22612 16952 22707 16980
rect 22612 16940 22618 16952
rect 22695 16949 22707 16952
rect 22741 16949 22753 16983
rect 22695 16943 22753 16949
rect 24118 16940 24124 16992
rect 24176 16980 24182 16992
rect 24673 16983 24731 16989
rect 24673 16980 24685 16983
rect 24176 16952 24685 16980
rect 24176 16940 24182 16952
rect 24673 16949 24685 16952
rect 24719 16949 24731 16983
rect 24673 16943 24731 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3145 16779 3203 16785
rect 3145 16776 3157 16779
rect 2924 16748 3157 16776
rect 2924 16736 2930 16748
rect 3145 16745 3157 16748
rect 3191 16745 3203 16779
rect 3510 16776 3516 16788
rect 3471 16748 3516 16776
rect 3145 16739 3203 16745
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 4246 16736 4252 16788
rect 4304 16776 4310 16788
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 4304 16748 4537 16776
rect 4304 16736 4310 16748
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 7558 16736 7564 16788
rect 7616 16776 7622 16788
rect 7837 16779 7895 16785
rect 7837 16776 7849 16779
rect 7616 16748 7849 16776
rect 7616 16736 7622 16748
rect 7837 16745 7849 16748
rect 7883 16745 7895 16779
rect 8294 16776 8300 16788
rect 8255 16748 8300 16776
rect 7837 16739 7895 16745
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 9125 16779 9183 16785
rect 9125 16745 9137 16779
rect 9171 16776 9183 16779
rect 9766 16776 9772 16788
rect 9171 16748 9772 16776
rect 9171 16745 9183 16748
rect 9125 16739 9183 16745
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 11238 16776 11244 16788
rect 11199 16748 11244 16776
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 11514 16736 11520 16788
rect 11572 16776 11578 16788
rect 12710 16776 12716 16788
rect 11572 16748 12716 16776
rect 11572 16736 11578 16748
rect 12710 16736 12716 16748
rect 12768 16776 12774 16788
rect 12989 16779 13047 16785
rect 12989 16776 13001 16779
rect 12768 16748 13001 16776
rect 12768 16736 12774 16748
rect 12989 16745 13001 16748
rect 13035 16745 13047 16779
rect 15378 16776 15384 16788
rect 15339 16748 15384 16776
rect 12989 16739 13047 16745
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 15470 16736 15476 16788
rect 15528 16776 15534 16788
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 15528 16748 16313 16776
rect 15528 16736 15534 16748
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 16301 16739 16359 16745
rect 16482 16736 16488 16788
rect 16540 16776 16546 16788
rect 16761 16779 16819 16785
rect 16761 16776 16773 16779
rect 16540 16748 16773 16776
rect 16540 16736 16546 16748
rect 16761 16745 16773 16748
rect 16807 16776 16819 16779
rect 17770 16776 17776 16788
rect 16807 16748 17776 16776
rect 16807 16745 16819 16748
rect 16761 16739 16819 16745
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 19935 16779 19993 16785
rect 19935 16745 19947 16779
rect 19981 16776 19993 16779
rect 20806 16776 20812 16788
rect 19981 16748 20812 16776
rect 19981 16745 19993 16748
rect 19935 16739 19993 16745
rect 20806 16736 20812 16748
rect 20864 16736 20870 16788
rect 20898 16736 20904 16788
rect 20956 16776 20962 16788
rect 22373 16779 22431 16785
rect 20956 16748 21128 16776
rect 20956 16736 20962 16748
rect 2222 16708 2228 16720
rect 2183 16680 2228 16708
rect 2222 16668 2228 16680
rect 2280 16668 2286 16720
rect 2777 16711 2835 16717
rect 2777 16677 2789 16711
rect 2823 16708 2835 16711
rect 3050 16708 3056 16720
rect 2823 16680 3056 16708
rect 2823 16677 2835 16680
rect 2777 16671 2835 16677
rect 3050 16668 3056 16680
rect 3108 16668 3114 16720
rect 6733 16711 6791 16717
rect 6733 16677 6745 16711
rect 6779 16708 6791 16711
rect 6822 16708 6828 16720
rect 6779 16680 6828 16708
rect 6779 16677 6791 16680
rect 6733 16671 6791 16677
rect 6822 16668 6828 16680
rect 6880 16708 6886 16720
rect 7009 16711 7067 16717
rect 7009 16708 7021 16711
rect 6880 16680 7021 16708
rect 6880 16668 6886 16680
rect 7009 16677 7021 16680
rect 7055 16677 7067 16711
rect 7009 16671 7067 16677
rect 10965 16711 11023 16717
rect 10965 16677 10977 16711
rect 11011 16708 11023 16711
rect 11974 16708 11980 16720
rect 11011 16680 11980 16708
rect 11011 16677 11023 16680
rect 10965 16671 11023 16677
rect 11974 16668 11980 16680
rect 12032 16668 12038 16720
rect 12155 16711 12213 16717
rect 12155 16677 12167 16711
rect 12201 16677 12213 16711
rect 12155 16671 12213 16677
rect 14369 16711 14427 16717
rect 14369 16677 14381 16711
rect 14415 16708 14427 16711
rect 15654 16708 15660 16720
rect 14415 16680 15660 16708
rect 14415 16677 14427 16680
rect 14369 16671 14427 16677
rect 4614 16640 4620 16652
rect 4575 16612 4620 16640
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 4982 16640 4988 16652
rect 4943 16612 4988 16640
rect 4982 16600 4988 16612
rect 5040 16600 5046 16652
rect 6181 16643 6239 16649
rect 6181 16609 6193 16643
rect 6227 16609 6239 16643
rect 6181 16603 6239 16609
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 7098 16640 7104 16652
rect 6595 16612 7104 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 2133 16575 2191 16581
rect 2133 16572 2145 16575
rect 1872 16544 2145 16572
rect 1578 16396 1584 16448
rect 1636 16436 1642 16448
rect 1872 16445 1900 16544
rect 2133 16541 2145 16544
rect 2179 16541 2191 16575
rect 2133 16535 2191 16541
rect 6086 16464 6092 16516
rect 6144 16504 6150 16516
rect 6196 16504 6224 16603
rect 7098 16600 7104 16612
rect 7156 16600 7162 16652
rect 8018 16640 8024 16652
rect 7979 16612 8024 16640
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 8573 16643 8631 16649
rect 8573 16640 8585 16643
rect 8352 16612 8585 16640
rect 8352 16600 8358 16612
rect 8573 16609 8585 16612
rect 8619 16640 8631 16643
rect 9858 16640 9864 16652
rect 8619 16612 9864 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10042 16600 10048 16652
rect 10100 16640 10106 16652
rect 10226 16640 10232 16652
rect 10100 16612 10232 16640
rect 10100 16600 10106 16612
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 10778 16640 10784 16652
rect 10739 16612 10784 16640
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 11882 16600 11888 16652
rect 11940 16640 11946 16652
rect 12170 16640 12198 16671
rect 15654 16668 15660 16680
rect 15712 16668 15718 16720
rect 19242 16708 19248 16720
rect 18156 16680 19248 16708
rect 13906 16640 13912 16652
rect 11940 16612 12198 16640
rect 13867 16612 13912 16640
rect 11940 16600 11946 16612
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 14185 16643 14243 16649
rect 14185 16609 14197 16643
rect 14231 16640 14243 16643
rect 14458 16640 14464 16652
rect 14231 16612 14464 16640
rect 14231 16609 14243 16612
rect 14185 16603 14243 16609
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 15470 16640 15476 16652
rect 15431 16612 15476 16640
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 15838 16640 15844 16652
rect 15799 16612 15844 16640
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 17770 16600 17776 16652
rect 17828 16640 17834 16652
rect 18156 16649 18184 16680
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 19705 16711 19763 16717
rect 19705 16677 19717 16711
rect 19751 16708 19763 16711
rect 20070 16708 20076 16720
rect 19751 16680 20076 16708
rect 19751 16677 19763 16680
rect 19705 16671 19763 16677
rect 20070 16668 20076 16680
rect 20128 16668 20134 16720
rect 20162 16668 20168 16720
rect 20220 16708 20226 16720
rect 21100 16717 21128 16748
rect 22373 16745 22385 16779
rect 22419 16776 22431 16779
rect 22554 16776 22560 16788
rect 22419 16748 22560 16776
rect 22419 16745 22431 16748
rect 22373 16739 22431 16745
rect 22554 16736 22560 16748
rect 22612 16736 22618 16788
rect 24167 16779 24225 16785
rect 24167 16745 24179 16779
rect 24213 16776 24225 16779
rect 24670 16776 24676 16788
rect 24213 16748 24676 16776
rect 24213 16745 24225 16748
rect 24167 16739 24225 16745
rect 24670 16736 24676 16748
rect 24728 16736 24734 16788
rect 20993 16711 21051 16717
rect 20993 16708 21005 16711
rect 20220 16680 21005 16708
rect 20220 16668 20226 16680
rect 20993 16677 21005 16680
rect 21039 16677 21051 16711
rect 20993 16671 21051 16677
rect 21085 16711 21143 16717
rect 21085 16677 21097 16711
rect 21131 16677 21143 16711
rect 21085 16671 21143 16677
rect 22649 16711 22707 16717
rect 22649 16677 22661 16711
rect 22695 16708 22707 16711
rect 22738 16708 22744 16720
rect 22695 16680 22744 16708
rect 22695 16677 22707 16680
rect 22649 16671 22707 16677
rect 22738 16668 22744 16680
rect 22796 16668 22802 16720
rect 23198 16708 23204 16720
rect 23159 16680 23204 16708
rect 23198 16668 23204 16680
rect 23256 16668 23262 16720
rect 18141 16643 18199 16649
rect 18141 16640 18153 16643
rect 17828 16612 18153 16640
rect 17828 16600 17834 16612
rect 18141 16609 18153 16612
rect 18187 16609 18199 16643
rect 18598 16640 18604 16652
rect 18559 16612 18604 16640
rect 18141 16603 18199 16609
rect 18598 16600 18604 16612
rect 18656 16600 18662 16652
rect 19794 16640 19800 16652
rect 19755 16612 19800 16640
rect 19794 16600 19800 16612
rect 19852 16640 19858 16652
rect 20622 16640 20628 16652
rect 19852 16612 20628 16640
rect 19852 16600 19858 16612
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 23934 16640 23940 16652
rect 23895 16612 23940 16640
rect 23934 16600 23940 16612
rect 23992 16600 23998 16652
rect 25092 16643 25150 16649
rect 25092 16609 25104 16643
rect 25138 16640 25150 16643
rect 25590 16640 25596 16652
rect 25138 16612 25596 16640
rect 25138 16609 25150 16612
rect 25092 16603 25150 16609
rect 25590 16600 25596 16612
rect 25648 16600 25654 16652
rect 11054 16572 11060 16584
rect 9646 16544 11060 16572
rect 9646 16504 9674 16544
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 11790 16572 11796 16584
rect 11751 16544 11796 16572
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 14274 16532 14280 16584
rect 14332 16572 14338 16584
rect 16853 16575 16911 16581
rect 16853 16572 16865 16575
rect 14332 16544 16865 16572
rect 14332 16532 14338 16544
rect 16853 16541 16865 16544
rect 16899 16541 16911 16575
rect 16853 16535 16911 16541
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19426 16572 19432 16584
rect 18923 16544 19432 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 21266 16572 21272 16584
rect 21227 16544 21272 16572
rect 21266 16532 21272 16544
rect 21324 16532 21330 16584
rect 22554 16572 22560 16584
rect 22515 16544 22560 16572
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 23750 16572 23756 16584
rect 23663 16544 23756 16572
rect 23750 16532 23756 16544
rect 23808 16572 23814 16584
rect 25179 16575 25237 16581
rect 25179 16572 25191 16575
rect 23808 16544 25191 16572
rect 23808 16532 23814 16544
rect 25179 16541 25191 16544
rect 25225 16541 25237 16575
rect 25179 16535 25237 16541
rect 6144 16476 9674 16504
rect 6144 16464 6150 16476
rect 10134 16464 10140 16516
rect 10192 16504 10198 16516
rect 17034 16504 17040 16516
rect 10192 16476 17040 16504
rect 10192 16464 10198 16476
rect 17034 16464 17040 16476
rect 17092 16464 17098 16516
rect 20717 16507 20775 16513
rect 20717 16473 20729 16507
rect 20763 16504 20775 16507
rect 21284 16504 21312 16532
rect 20763 16476 21312 16504
rect 20763 16473 20775 16476
rect 20717 16467 20775 16473
rect 1857 16439 1915 16445
rect 1857 16436 1869 16439
rect 1636 16408 1869 16436
rect 1636 16396 1642 16408
rect 1857 16405 1869 16408
rect 1903 16405 1915 16439
rect 1857 16399 1915 16405
rect 4154 16396 4160 16448
rect 4212 16436 4218 16448
rect 4341 16439 4399 16445
rect 4341 16436 4353 16439
rect 4212 16408 4353 16436
rect 4212 16396 4218 16408
rect 4341 16405 4353 16408
rect 4387 16436 4399 16439
rect 4522 16436 4528 16448
rect 4387 16408 4528 16436
rect 4387 16405 4399 16408
rect 4341 16399 4399 16405
rect 4522 16396 4528 16408
rect 4580 16396 4586 16448
rect 12713 16439 12771 16445
rect 12713 16405 12725 16439
rect 12759 16436 12771 16439
rect 12802 16436 12808 16448
rect 12759 16408 12808 16436
rect 12759 16405 12771 16408
rect 12713 16399 12771 16405
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 13354 16436 13360 16448
rect 13315 16408 13360 16436
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 17586 16396 17592 16448
rect 17644 16436 17650 16448
rect 17957 16439 18015 16445
rect 17957 16436 17969 16439
rect 17644 16408 17969 16436
rect 17644 16396 17650 16408
rect 17957 16405 17969 16408
rect 18003 16405 18015 16439
rect 17957 16399 18015 16405
rect 18230 16396 18236 16448
rect 18288 16436 18294 16448
rect 19058 16436 19064 16448
rect 18288 16408 19064 16436
rect 18288 16396 18294 16408
rect 19058 16396 19064 16408
rect 19116 16436 19122 16448
rect 19245 16439 19303 16445
rect 19245 16436 19257 16439
rect 19116 16408 19257 16436
rect 19116 16396 19122 16408
rect 19245 16405 19257 16408
rect 19291 16405 19303 16439
rect 19245 16399 19303 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1854 16232 1860 16244
rect 1815 16204 1860 16232
rect 1854 16192 1860 16204
rect 1912 16192 1918 16244
rect 2222 16192 2228 16244
rect 2280 16232 2286 16244
rect 2961 16235 3019 16241
rect 2961 16232 2973 16235
rect 2280 16204 2973 16232
rect 2280 16192 2286 16204
rect 2961 16201 2973 16204
rect 3007 16201 3019 16235
rect 6086 16232 6092 16244
rect 6047 16204 6092 16232
rect 2961 16195 3019 16201
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 8018 16232 8024 16244
rect 7979 16204 8024 16232
rect 8018 16192 8024 16204
rect 8076 16192 8082 16244
rect 11882 16232 11888 16244
rect 11843 16204 11888 16232
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 14093 16235 14151 16241
rect 14093 16201 14105 16235
rect 14139 16232 14151 16235
rect 14458 16232 14464 16244
rect 14139 16204 14464 16232
rect 14139 16201 14151 16204
rect 14093 16195 14151 16201
rect 14458 16192 14464 16204
rect 14516 16192 14522 16244
rect 20162 16232 20168 16244
rect 20123 16204 20168 16232
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 20898 16192 20904 16244
rect 20956 16232 20962 16244
rect 21729 16235 21787 16241
rect 21729 16232 21741 16235
rect 20956 16204 21741 16232
rect 20956 16192 20962 16204
rect 21729 16201 21741 16204
rect 21775 16201 21787 16235
rect 21729 16195 21787 16201
rect 22554 16192 22560 16244
rect 22612 16232 22618 16244
rect 23109 16235 23167 16241
rect 23109 16232 23121 16235
rect 22612 16204 23121 16232
rect 22612 16192 22618 16204
rect 23109 16201 23121 16204
rect 23155 16232 23167 16235
rect 23155 16204 23474 16232
rect 23155 16201 23167 16204
rect 23109 16195 23167 16201
rect 2590 16164 2596 16176
rect 2551 16136 2596 16164
rect 2590 16124 2596 16136
rect 2648 16124 2654 16176
rect 4614 16124 4620 16176
rect 4672 16164 4678 16176
rect 10686 16164 10692 16176
rect 4672 16136 10692 16164
rect 4672 16124 4678 16136
rect 10686 16124 10692 16136
rect 10744 16124 10750 16176
rect 11238 16124 11244 16176
rect 11296 16164 11302 16176
rect 18233 16167 18291 16173
rect 18233 16164 18245 16167
rect 11296 16136 11376 16164
rect 11296 16124 11302 16136
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 2130 16096 2136 16108
rect 2087 16068 2136 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 3050 16056 3056 16108
rect 3108 16096 3114 16108
rect 3881 16099 3939 16105
rect 3881 16096 3893 16099
rect 3108 16068 3893 16096
rect 3108 16056 3114 16068
rect 3881 16065 3893 16068
rect 3927 16065 3939 16099
rect 4982 16096 4988 16108
rect 4895 16068 4988 16096
rect 3881 16059 3939 16065
rect 4982 16056 4988 16068
rect 5040 16096 5046 16108
rect 10226 16096 10232 16108
rect 5040 16068 7144 16096
rect 5040 16056 5046 16068
rect 5258 16028 5264 16040
rect 5219 16000 5264 16028
rect 5258 15988 5264 16000
rect 5316 15988 5322 16040
rect 5644 16037 5672 16068
rect 7116 16040 7144 16068
rect 9048 16068 10232 16096
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 15997 5687 16031
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 5629 15991 5687 15997
rect 6564 16000 6837 16028
rect 1854 15920 1860 15972
rect 1912 15960 1918 15972
rect 2133 15963 2191 15969
rect 2133 15960 2145 15963
rect 1912 15932 2145 15960
rect 1912 15920 1918 15932
rect 2133 15929 2145 15932
rect 2179 15929 2191 15963
rect 3602 15960 3608 15972
rect 3563 15932 3608 15960
rect 2133 15923 2191 15929
rect 3602 15920 3608 15932
rect 3660 15920 3666 15972
rect 3697 15963 3755 15969
rect 3697 15929 3709 15963
rect 3743 15929 3755 15963
rect 3697 15923 3755 15929
rect 3418 15892 3424 15904
rect 3379 15864 3424 15892
rect 3418 15852 3424 15864
rect 3476 15892 3482 15904
rect 3712 15892 3740 15923
rect 4614 15892 4620 15904
rect 3476 15864 3740 15892
rect 4575 15864 4620 15892
rect 3476 15852 3482 15864
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 6564 15901 6592 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 7377 16031 7435 16037
rect 7377 16028 7389 16031
rect 7156 16000 7389 16028
rect 7156 15988 7162 16000
rect 7377 15997 7389 16000
rect 7423 16028 7435 16031
rect 8294 16028 8300 16040
rect 7423 16000 8300 16028
rect 7423 15997 7435 16000
rect 7377 15991 7435 15997
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 9048 16037 9076 16068
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 11348 16105 11376 16136
rect 15850 16136 18245 16164
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16065 11391 16099
rect 12710 16096 12716 16108
rect 12671 16068 12716 16096
rect 11333 16059 11391 16065
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 15746 16096 15752 16108
rect 15120 16068 15752 16096
rect 9033 16031 9091 16037
rect 9033 16028 9045 16031
rect 8588 16000 9045 16028
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 6420 15864 6561 15892
rect 6420 15852 6426 15864
rect 6549 15861 6561 15864
rect 6595 15861 6607 15895
rect 6914 15892 6920 15904
rect 6875 15864 6920 15892
rect 6549 15855 6607 15861
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 8588 15901 8616 16000
rect 9033 15997 9045 16000
rect 9079 15997 9091 16031
rect 9033 15991 9091 15997
rect 9309 16031 9367 16037
rect 9309 15997 9321 16031
rect 9355 16028 9367 16031
rect 9674 16028 9680 16040
rect 9355 16000 9680 16028
rect 9355 15997 9367 16000
rect 9309 15991 9367 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 16028 10747 16031
rect 11054 16028 11060 16040
rect 10735 16000 11060 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 11054 15988 11060 16000
rect 11112 15988 11118 16040
rect 11241 16031 11299 16037
rect 11241 15997 11253 16031
rect 11287 15997 11299 16031
rect 11241 15991 11299 15997
rect 11256 15960 11284 15991
rect 14918 15988 14924 16040
rect 14976 16028 14982 16040
rect 15120 16037 15148 16068
rect 15746 16056 15752 16068
rect 15804 16056 15810 16108
rect 15105 16031 15163 16037
rect 15105 16028 15117 16031
rect 14976 16000 15117 16028
rect 14976 15988 14982 16000
rect 15105 15997 15117 16000
rect 15151 15997 15163 16031
rect 15105 15991 15163 15997
rect 15289 16031 15347 16037
rect 15289 15997 15301 16031
rect 15335 16028 15347 16031
rect 15850 16028 15878 16136
rect 18233 16133 18245 16136
rect 18279 16164 18291 16167
rect 18598 16164 18604 16176
rect 18279 16136 18604 16164
rect 18279 16133 18291 16136
rect 18233 16127 18291 16133
rect 18598 16124 18604 16136
rect 18656 16124 18662 16176
rect 21358 16164 21364 16176
rect 21319 16136 21364 16164
rect 21358 16124 21364 16136
rect 21416 16124 21422 16176
rect 22738 16164 22744 16176
rect 22699 16136 22744 16164
rect 22738 16124 22744 16136
rect 22796 16124 22802 16176
rect 23446 16164 23474 16204
rect 23934 16192 23940 16244
rect 23992 16232 23998 16244
rect 24489 16235 24547 16241
rect 24489 16232 24501 16235
rect 23992 16204 24501 16232
rect 23992 16192 23998 16204
rect 24489 16201 24501 16204
rect 24535 16201 24547 16235
rect 24489 16195 24547 16201
rect 24578 16164 24584 16176
rect 23446 16136 24584 16164
rect 24578 16124 24584 16136
rect 24636 16124 24642 16176
rect 16482 16096 16488 16108
rect 16443 16068 16488 16096
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 17954 16056 17960 16108
rect 18012 16096 18018 16108
rect 19794 16096 19800 16108
rect 18012 16068 19800 16096
rect 18012 16056 18018 16068
rect 19794 16056 19800 16068
rect 19852 16056 19858 16108
rect 20806 16096 20812 16108
rect 20719 16068 20812 16096
rect 20806 16056 20812 16068
rect 20864 16096 20870 16108
rect 22097 16099 22155 16105
rect 22097 16096 22109 16099
rect 20864 16068 22109 16096
rect 20864 16056 20870 16068
rect 22097 16065 22109 16068
rect 22143 16065 22155 16099
rect 24213 16099 24271 16105
rect 24213 16096 24225 16099
rect 22097 16059 22155 16065
rect 23743 16068 24225 16096
rect 23743 16037 23771 16068
rect 24213 16065 24225 16068
rect 24259 16096 24271 16099
rect 24854 16096 24860 16108
rect 24259 16068 24860 16096
rect 24259 16065 24271 16068
rect 24213 16059 24271 16065
rect 24854 16056 24860 16068
rect 24912 16056 24918 16108
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16096 25283 16099
rect 27614 16096 27620 16108
rect 25271 16068 27620 16096
rect 25271 16065 25283 16068
rect 25225 16059 25283 16065
rect 15335 16000 15878 16028
rect 23728 16031 23786 16037
rect 15335 15997 15347 16000
rect 15289 15991 15347 15997
rect 23728 15997 23740 16031
rect 23774 15997 23786 16031
rect 23728 15991 23786 15997
rect 24740 16031 24798 16037
rect 24740 15997 24752 16031
rect 24786 16028 24798 16031
rect 25240 16028 25268 16059
rect 27614 16056 27620 16068
rect 27672 16056 27678 16108
rect 24786 16000 25268 16028
rect 24786 15997 24798 16000
rect 24740 15991 24798 15997
rect 11072 15932 11284 15960
rect 11072 15904 11100 15932
rect 12802 15920 12808 15972
rect 12860 15960 12866 15972
rect 13357 15963 13415 15969
rect 12860 15932 12905 15960
rect 12860 15920 12866 15932
rect 13357 15929 13369 15963
rect 13403 15960 13415 15963
rect 13446 15960 13452 15972
rect 13403 15932 13452 15960
rect 13403 15929 13415 15932
rect 13357 15923 13415 15929
rect 13446 15920 13452 15932
rect 13504 15920 13510 15972
rect 15304 15960 15332 15991
rect 15562 15960 15568 15972
rect 14660 15932 15332 15960
rect 15523 15932 15568 15960
rect 8573 15895 8631 15901
rect 8573 15892 8585 15895
rect 8444 15864 8585 15892
rect 8444 15852 8450 15864
rect 8573 15861 8585 15864
rect 8619 15861 8631 15895
rect 8846 15892 8852 15904
rect 8807 15864 8852 15892
rect 8573 15855 8631 15861
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 9953 15895 10011 15901
rect 9953 15861 9965 15895
rect 9999 15892 10011 15895
rect 10778 15892 10784 15904
rect 9999 15864 10784 15892
rect 9999 15861 10011 15864
rect 9953 15855 10011 15861
rect 10778 15852 10784 15864
rect 10836 15892 10842 15904
rect 11054 15892 11060 15904
rect 10836 15864 11060 15892
rect 10836 15852 10842 15864
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 12253 15895 12311 15901
rect 12253 15861 12265 15895
rect 12299 15892 12311 15895
rect 12820 15892 12848 15920
rect 12299 15864 12848 15892
rect 13725 15895 13783 15901
rect 12299 15861 12311 15864
rect 12253 15855 12311 15861
rect 13725 15861 13737 15895
rect 13771 15892 13783 15895
rect 13906 15892 13912 15904
rect 13771 15864 13912 15892
rect 13771 15861 13783 15864
rect 13725 15855 13783 15861
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 14550 15852 14556 15904
rect 14608 15892 14614 15904
rect 14660 15901 14688 15932
rect 15562 15920 15568 15932
rect 15620 15920 15626 15972
rect 16301 15963 16359 15969
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 16574 15960 16580 15972
rect 16347 15932 16580 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 17129 15963 17187 15969
rect 17129 15929 17141 15963
rect 17175 15960 17187 15963
rect 17586 15960 17592 15972
rect 17175 15932 17592 15960
rect 17175 15929 17187 15932
rect 17129 15923 17187 15929
rect 17586 15920 17592 15932
rect 17644 15960 17650 15972
rect 18601 15963 18659 15969
rect 18601 15960 18613 15963
rect 17644 15932 18613 15960
rect 17644 15920 17650 15932
rect 18601 15929 18613 15932
rect 18647 15929 18659 15963
rect 18601 15923 18659 15929
rect 18690 15920 18696 15972
rect 18748 15960 18754 15972
rect 19242 15960 19248 15972
rect 18748 15932 18793 15960
rect 19203 15932 19248 15960
rect 18748 15920 18754 15932
rect 19242 15920 19248 15932
rect 19300 15920 19306 15972
rect 20901 15963 20959 15969
rect 20901 15929 20913 15963
rect 20947 15929 20959 15963
rect 20901 15923 20959 15929
rect 14645 15895 14703 15901
rect 14645 15892 14657 15895
rect 14608 15864 14657 15892
rect 14608 15852 14614 15864
rect 14645 15861 14657 15864
rect 14691 15861 14703 15895
rect 14645 15855 14703 15861
rect 15470 15852 15476 15904
rect 15528 15892 15534 15904
rect 15930 15892 15936 15904
rect 15528 15864 15936 15892
rect 15528 15852 15534 15864
rect 15930 15852 15936 15864
rect 15988 15852 15994 15904
rect 17770 15892 17776 15904
rect 17731 15864 17776 15892
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 20530 15892 20536 15904
rect 20491 15864 20536 15892
rect 20530 15852 20536 15864
rect 20588 15892 20594 15904
rect 20916 15892 20944 15923
rect 22278 15892 22284 15904
rect 20588 15864 20944 15892
rect 22239 15864 22284 15892
rect 20588 15852 20594 15864
rect 22278 15852 22284 15864
rect 22336 15852 22342 15904
rect 23799 15895 23857 15901
rect 23799 15861 23811 15895
rect 23845 15892 23857 15895
rect 23934 15892 23940 15904
rect 23845 15864 23940 15892
rect 23845 15861 23857 15864
rect 23799 15855 23857 15861
rect 23934 15852 23940 15864
rect 23992 15852 23998 15904
rect 24670 15852 24676 15904
rect 24728 15892 24734 15904
rect 24811 15895 24869 15901
rect 24811 15892 24823 15895
rect 24728 15864 24823 15892
rect 24728 15852 24734 15864
rect 24811 15861 24823 15864
rect 24857 15861 24869 15895
rect 25590 15892 25596 15904
rect 25551 15864 25596 15892
rect 24811 15855 24869 15861
rect 25590 15852 25596 15864
rect 25648 15852 25654 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1857 15691 1915 15697
rect 1857 15657 1869 15691
rect 1903 15688 1915 15691
rect 2038 15688 2044 15700
rect 1903 15660 2044 15688
rect 1903 15657 1915 15660
rect 1857 15651 1915 15657
rect 2038 15648 2044 15660
rect 2096 15648 2102 15700
rect 3050 15688 3056 15700
rect 2700 15660 3056 15688
rect 2700 15632 2728 15660
rect 3050 15648 3056 15660
rect 3108 15648 3114 15700
rect 3418 15648 3424 15700
rect 3476 15688 3482 15700
rect 8294 15688 8300 15700
rect 3476 15660 7420 15688
rect 8255 15660 8300 15688
rect 3476 15648 3482 15660
rect 2133 15623 2191 15629
rect 2133 15589 2145 15623
rect 2179 15620 2191 15623
rect 2498 15620 2504 15632
rect 2179 15592 2504 15620
rect 2179 15589 2191 15592
rect 2133 15583 2191 15589
rect 2498 15580 2504 15592
rect 2556 15580 2562 15632
rect 2682 15620 2688 15632
rect 2595 15592 2688 15620
rect 2682 15580 2688 15592
rect 2740 15580 2746 15632
rect 3970 15580 3976 15632
rect 4028 15620 4034 15632
rect 4249 15623 4307 15629
rect 4249 15620 4261 15623
rect 4028 15592 4261 15620
rect 4028 15580 4034 15592
rect 4249 15589 4261 15592
rect 4295 15589 4307 15623
rect 4249 15583 4307 15589
rect 4982 15580 4988 15632
rect 5040 15620 5046 15632
rect 5077 15623 5135 15629
rect 5077 15620 5089 15623
rect 5040 15592 5089 15620
rect 5040 15580 5046 15592
rect 5077 15589 5089 15592
rect 5123 15589 5135 15623
rect 5077 15583 5135 15589
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 5813 15623 5871 15629
rect 5813 15620 5825 15623
rect 5500 15592 5825 15620
rect 5500 15580 5506 15592
rect 5813 15589 5825 15592
rect 5859 15589 5871 15623
rect 5813 15583 5871 15589
rect 6733 15623 6791 15629
rect 6733 15589 6745 15623
rect 6779 15620 6791 15623
rect 7098 15620 7104 15632
rect 6779 15592 7104 15620
rect 6779 15589 6791 15592
rect 6733 15583 6791 15589
rect 7098 15580 7104 15592
rect 7156 15580 7162 15632
rect 7282 15620 7288 15632
rect 7243 15592 7288 15620
rect 7282 15580 7288 15592
rect 7340 15580 7346 15632
rect 7392 15629 7420 15660
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 9674 15688 9680 15700
rect 9539 15660 9680 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 14918 15688 14924 15700
rect 14879 15660 14924 15688
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 15565 15691 15623 15697
rect 15565 15657 15577 15691
rect 15611 15688 15623 15691
rect 15838 15688 15844 15700
rect 15611 15660 15844 15688
rect 15611 15657 15623 15660
rect 15565 15651 15623 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 16114 15688 16120 15700
rect 16027 15660 16120 15688
rect 16114 15648 16120 15660
rect 16172 15688 16178 15700
rect 18230 15688 18236 15700
rect 16172 15660 18236 15688
rect 16172 15648 16178 15660
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 18690 15648 18696 15700
rect 18748 15688 18754 15700
rect 18785 15691 18843 15697
rect 18785 15688 18797 15691
rect 18748 15660 18797 15688
rect 18748 15648 18754 15660
rect 18785 15657 18797 15660
rect 18831 15688 18843 15691
rect 19061 15691 19119 15697
rect 19061 15688 19073 15691
rect 18831 15660 19073 15688
rect 18831 15657 18843 15660
rect 18785 15651 18843 15657
rect 19061 15657 19073 15660
rect 19107 15657 19119 15691
rect 19426 15688 19432 15700
rect 19387 15660 19432 15688
rect 19061 15651 19119 15657
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 19935 15691 19993 15697
rect 19935 15657 19947 15691
rect 19981 15688 19993 15691
rect 20806 15688 20812 15700
rect 19981 15660 20812 15688
rect 19981 15657 19993 15660
rect 19935 15651 19993 15657
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 23934 15688 23940 15700
rect 23895 15660 23940 15688
rect 23934 15648 23940 15660
rect 23992 15648 23998 15700
rect 24578 15648 24584 15700
rect 24636 15688 24642 15700
rect 24719 15691 24777 15697
rect 24719 15688 24731 15691
rect 24636 15660 24731 15688
rect 24636 15648 24642 15660
rect 24719 15657 24731 15660
rect 24765 15657 24777 15691
rect 24719 15651 24777 15657
rect 7377 15623 7435 15629
rect 7377 15589 7389 15623
rect 7423 15620 7435 15623
rect 7742 15620 7748 15632
rect 7423 15592 7748 15620
rect 7423 15589 7435 15592
rect 7377 15583 7435 15589
rect 7742 15580 7748 15592
rect 7800 15580 7806 15632
rect 9858 15620 9864 15632
rect 9819 15592 9864 15620
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 11054 15580 11060 15632
rect 11112 15620 11118 15632
rect 13078 15620 13084 15632
rect 11112 15592 11744 15620
rect 13039 15592 13084 15620
rect 11112 15580 11118 15592
rect 5258 15512 5264 15564
rect 5316 15552 5322 15564
rect 5316 15524 5488 15552
rect 5316 15512 5322 15524
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15484 2099 15487
rect 2406 15484 2412 15496
rect 2087 15456 2412 15484
rect 2087 15453 2099 15456
rect 2041 15447 2099 15453
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 3510 15444 3516 15496
rect 3568 15484 3574 15496
rect 5460 15493 5488 15524
rect 10686 15512 10692 15564
rect 10744 15552 10750 15564
rect 11238 15552 11244 15564
rect 10744 15524 11244 15552
rect 10744 15512 10750 15524
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11716 15561 11744 15592
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 13446 15580 13452 15632
rect 13504 15620 13510 15632
rect 13633 15623 13691 15629
rect 13633 15620 13645 15623
rect 13504 15592 13645 15620
rect 13504 15580 13510 15592
rect 13633 15589 13645 15592
rect 13679 15589 13691 15623
rect 21082 15620 21088 15632
rect 21043 15592 21088 15620
rect 13633 15583 13691 15589
rect 21082 15580 21088 15592
rect 21140 15580 21146 15632
rect 23106 15620 23112 15632
rect 23067 15592 23112 15620
rect 23106 15580 23112 15592
rect 23164 15580 23170 15632
rect 23661 15623 23719 15629
rect 23661 15589 23673 15623
rect 23707 15620 23719 15623
rect 23842 15620 23848 15632
rect 23707 15592 23848 15620
rect 23707 15589 23719 15592
rect 23661 15583 23719 15589
rect 11701 15555 11759 15561
rect 11701 15521 11713 15555
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 18046 15512 18052 15564
rect 18104 15552 18110 15564
rect 19864 15555 19922 15561
rect 19864 15552 19876 15555
rect 18104 15524 19876 15552
rect 18104 15512 18110 15524
rect 19864 15521 19876 15524
rect 19910 15552 19922 15555
rect 20254 15552 20260 15564
rect 19910 15524 20260 15552
rect 19910 15521 19922 15524
rect 19864 15515 19922 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 4157 15487 4215 15493
rect 4157 15484 4169 15487
rect 3568 15456 4169 15484
rect 3568 15444 3574 15456
rect 4157 15453 4169 15456
rect 4203 15484 4215 15487
rect 5445 15487 5503 15493
rect 4203 15456 4844 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 3326 15376 3332 15428
rect 3384 15416 3390 15428
rect 4709 15419 4767 15425
rect 4709 15416 4721 15419
rect 3384 15388 4721 15416
rect 3384 15376 3390 15388
rect 4709 15385 4721 15388
rect 4755 15385 4767 15419
rect 4816 15416 4844 15456
rect 5445 15453 5457 15487
rect 5491 15453 5503 15487
rect 5445 15447 5503 15453
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 5721 15487 5779 15493
rect 5721 15484 5733 15487
rect 5592 15456 5733 15484
rect 5592 15444 5598 15456
rect 5721 15453 5733 15456
rect 5767 15453 5779 15487
rect 5997 15487 6055 15493
rect 5997 15484 6009 15487
rect 5721 15447 5779 15453
rect 5828 15456 6009 15484
rect 5828 15416 5856 15456
rect 5997 15453 6009 15456
rect 6043 15453 6055 15487
rect 5997 15447 6055 15453
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8202 15484 8208 15496
rect 7975 15456 8208 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8202 15444 8208 15456
rect 8260 15484 8266 15496
rect 9766 15484 9772 15496
rect 8260 15456 9772 15484
rect 8260 15444 8266 15456
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 11790 15484 11796 15496
rect 11751 15456 11796 15484
rect 11790 15444 11796 15456
rect 11848 15484 11854 15496
rect 12253 15487 12311 15493
rect 12253 15484 12265 15487
rect 11848 15456 12265 15484
rect 11848 15444 11854 15456
rect 12253 15453 12265 15456
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15484 13047 15487
rect 13814 15484 13820 15496
rect 13035 15456 13820 15484
rect 13035 15453 13047 15456
rect 12989 15447 13047 15453
rect 13814 15444 13820 15456
rect 13872 15484 13878 15496
rect 14274 15484 14280 15496
rect 13872 15456 14280 15484
rect 13872 15444 13878 15456
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 14366 15444 14372 15496
rect 14424 15484 14430 15496
rect 15749 15487 15807 15493
rect 15749 15484 15761 15487
rect 14424 15456 15761 15484
rect 14424 15444 14430 15456
rect 15749 15453 15761 15456
rect 15795 15484 15807 15487
rect 17218 15484 17224 15496
rect 15795 15456 17224 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 17862 15484 17868 15496
rect 17823 15456 17868 15484
rect 17862 15444 17868 15456
rect 17920 15444 17926 15496
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15484 20775 15487
rect 20993 15487 21051 15493
rect 20993 15484 21005 15487
rect 20763 15456 21005 15484
rect 20763 15453 20775 15456
rect 20717 15447 20775 15453
rect 20993 15453 21005 15456
rect 21039 15484 21051 15487
rect 21358 15484 21364 15496
rect 21039 15456 21364 15484
rect 21039 15453 21051 15456
rect 20993 15447 21051 15453
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 22833 15487 22891 15493
rect 22833 15453 22845 15487
rect 22879 15484 22891 15487
rect 23017 15487 23075 15493
rect 23017 15484 23029 15487
rect 22879 15456 23029 15484
rect 22879 15453 22891 15456
rect 22833 15447 22891 15453
rect 23017 15453 23029 15456
rect 23063 15484 23075 15487
rect 23474 15484 23480 15496
rect 23063 15456 23480 15484
rect 23063 15453 23075 15456
rect 23017 15447 23075 15453
rect 23474 15444 23480 15456
rect 23532 15444 23538 15496
rect 10321 15419 10379 15425
rect 10321 15416 10333 15419
rect 4816 15388 5856 15416
rect 6104 15388 10333 15416
rect 4709 15379 4767 15385
rect 3881 15351 3939 15357
rect 3881 15317 3893 15351
rect 3927 15348 3939 15351
rect 4430 15348 4436 15360
rect 3927 15320 4436 15348
rect 3927 15317 3939 15320
rect 3881 15311 3939 15317
rect 4430 15308 4436 15320
rect 4488 15308 4494 15360
rect 4724 15348 4752 15379
rect 5350 15348 5356 15360
rect 4724 15320 5356 15348
rect 5350 15308 5356 15320
rect 5408 15348 5414 15360
rect 6104 15348 6132 15388
rect 10321 15385 10333 15388
rect 10367 15385 10379 15419
rect 14918 15416 14924 15428
rect 10321 15379 10379 15385
rect 13786 15388 14924 15416
rect 5408 15320 6132 15348
rect 5408 15308 5414 15320
rect 8570 15308 8576 15360
rect 8628 15348 8634 15360
rect 8757 15351 8815 15357
rect 8757 15348 8769 15351
rect 8628 15320 8769 15348
rect 8628 15308 8634 15320
rect 8757 15317 8769 15320
rect 8803 15348 8815 15351
rect 9493 15351 9551 15357
rect 9493 15348 9505 15351
rect 8803 15320 9505 15348
rect 8803 15317 8815 15320
rect 8757 15311 8815 15317
rect 9493 15317 9505 15320
rect 9539 15317 9551 15351
rect 9493 15311 9551 15317
rect 10873 15351 10931 15357
rect 10873 15317 10885 15351
rect 10919 15348 10931 15351
rect 11054 15348 11060 15360
rect 10919 15320 11060 15348
rect 10919 15317 10931 15320
rect 10873 15311 10931 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 12710 15348 12716 15360
rect 12671 15320 12716 15348
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 12894 15308 12900 15360
rect 12952 15348 12958 15360
rect 13786 15348 13814 15388
rect 14918 15376 14924 15388
rect 14976 15376 14982 15428
rect 19242 15376 19248 15428
rect 19300 15416 19306 15428
rect 21545 15419 21603 15425
rect 21545 15416 21557 15419
rect 19300 15388 21557 15416
rect 19300 15376 19306 15388
rect 21545 15385 21557 15388
rect 21591 15416 21603 15419
rect 23676 15416 23704 15583
rect 23842 15580 23848 15592
rect 23900 15580 23906 15632
rect 24648 15555 24706 15561
rect 24648 15521 24660 15555
rect 24694 15552 24706 15555
rect 24762 15552 24768 15564
rect 24694 15524 24768 15552
rect 24694 15521 24706 15524
rect 24648 15515 24706 15521
rect 24762 15512 24768 15524
rect 24820 15512 24826 15564
rect 21591 15388 23704 15416
rect 21591 15385 21603 15388
rect 21545 15379 21603 15385
rect 16666 15348 16672 15360
rect 12952 15320 13814 15348
rect 16627 15320 16672 15348
rect 12952 15308 12958 15320
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 4065 15147 4123 15153
rect 4065 15113 4077 15147
rect 4111 15144 4123 15147
rect 4522 15144 4528 15156
rect 4111 15116 4528 15144
rect 4111 15113 4123 15116
rect 4065 15107 4123 15113
rect 4522 15104 4528 15116
rect 4580 15104 4586 15156
rect 7742 15144 7748 15156
rect 7703 15116 7748 15144
rect 7742 15104 7748 15116
rect 7800 15144 7806 15156
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 7800 15116 8033 15144
rect 7800 15104 7806 15116
rect 8021 15113 8033 15116
rect 8067 15113 8079 15147
rect 9858 15144 9864 15156
rect 9819 15116 9864 15144
rect 8021 15107 8079 15113
rect 9858 15104 9864 15116
rect 9916 15144 9922 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 9916 15116 10149 15144
rect 9916 15104 9922 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 11940 15116 12173 15144
rect 11940 15104 11946 15116
rect 12161 15113 12173 15116
rect 12207 15144 12219 15147
rect 12437 15147 12495 15153
rect 12437 15144 12449 15147
rect 12207 15116 12449 15144
rect 12207 15113 12219 15116
rect 12161 15107 12219 15113
rect 12437 15113 12449 15116
rect 12483 15113 12495 15147
rect 12437 15107 12495 15113
rect 13078 15104 13084 15156
rect 13136 15144 13142 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13136 15116 13461 15144
rect 13136 15104 13142 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 17218 15144 17224 15156
rect 13872 15116 13917 15144
rect 17179 15116 17224 15144
rect 13872 15104 13878 15116
rect 17218 15104 17224 15116
rect 17276 15104 17282 15156
rect 20257 15147 20315 15153
rect 20257 15113 20269 15147
rect 20303 15144 20315 15147
rect 20622 15144 20628 15156
rect 20303 15116 20628 15144
rect 20303 15113 20315 15116
rect 20257 15107 20315 15113
rect 20622 15104 20628 15116
rect 20680 15144 20686 15156
rect 21082 15144 21088 15156
rect 20680 15116 21088 15144
rect 20680 15104 20686 15116
rect 21082 15104 21088 15116
rect 21140 15104 21146 15156
rect 22649 15147 22707 15153
rect 22649 15113 22661 15147
rect 22695 15144 22707 15147
rect 23017 15147 23075 15153
rect 23017 15144 23029 15147
rect 22695 15116 23029 15144
rect 22695 15113 22707 15116
rect 22649 15107 22707 15113
rect 23017 15113 23029 15116
rect 23063 15144 23075 15147
rect 23106 15144 23112 15156
rect 23063 15116 23112 15144
rect 23063 15113 23075 15116
rect 23017 15107 23075 15113
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 2038 15036 2044 15088
rect 2096 15076 2102 15088
rect 5442 15076 5448 15088
rect 2096 15048 5448 15076
rect 2096 15036 2102 15048
rect 5442 15036 5448 15048
rect 5500 15076 5506 15088
rect 5629 15079 5687 15085
rect 5629 15076 5641 15079
rect 5500 15048 5641 15076
rect 5500 15036 5506 15048
rect 5629 15045 5641 15048
rect 5675 15045 5687 15079
rect 5629 15039 5687 15045
rect 9766 15036 9772 15088
rect 9824 15076 9830 15088
rect 11333 15079 11391 15085
rect 11333 15076 11345 15079
rect 9824 15048 11345 15076
rect 9824 15036 9830 15048
rect 11333 15045 11345 15048
rect 11379 15045 11391 15079
rect 11333 15039 11391 15045
rect 15562 15036 15568 15088
rect 15620 15076 15626 15088
rect 21177 15079 21235 15085
rect 21177 15076 21189 15079
rect 15620 15048 21189 15076
rect 15620 15036 15626 15048
rect 21177 15045 21189 15048
rect 21223 15045 21235 15079
rect 21177 15039 21235 15045
rect 2682 15008 2688 15020
rect 2643 14980 2688 15008
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 3326 15008 3332 15020
rect 3287 14980 3332 15008
rect 3326 14968 3332 14980
rect 3384 14968 3390 15020
rect 3620 14980 4614 15008
rect 1448 14943 1506 14949
rect 1448 14909 1460 14943
rect 1494 14940 1506 14943
rect 1854 14940 1860 14952
rect 1494 14912 1860 14940
rect 1494 14909 1506 14912
rect 1448 14903 1506 14909
rect 1854 14900 1860 14912
rect 1912 14900 1918 14952
rect 1535 14875 1593 14881
rect 1535 14841 1547 14875
rect 1581 14872 1593 14875
rect 1946 14872 1952 14884
rect 1581 14844 1952 14872
rect 1581 14841 1593 14844
rect 1535 14835 1593 14841
rect 1946 14832 1952 14844
rect 2004 14832 2010 14884
rect 2777 14875 2835 14881
rect 2777 14841 2789 14875
rect 2823 14872 2835 14875
rect 2958 14872 2964 14884
rect 2823 14844 2964 14872
rect 2823 14841 2835 14844
rect 2777 14835 2835 14841
rect 2958 14832 2964 14844
rect 3016 14872 3022 14884
rect 3620 14872 3648 14980
rect 4157 14943 4215 14949
rect 4157 14909 4169 14943
rect 4203 14940 4215 14943
rect 4430 14940 4436 14952
rect 4203 14912 4436 14940
rect 4203 14909 4215 14912
rect 4157 14903 4215 14909
rect 4430 14900 4436 14912
rect 4488 14900 4494 14952
rect 4586 14940 4614 14980
rect 8846 14968 8852 15020
rect 8904 15008 8910 15020
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8904 14980 8953 15008
rect 8904 14968 8910 14980
rect 8941 14977 8953 14980
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 10781 15011 10839 15017
rect 10781 14977 10793 15011
rect 10827 15008 10839 15011
rect 10870 15008 10876 15020
rect 10827 14980 10876 15008
rect 10827 14977 10839 14980
rect 10781 14971 10839 14977
rect 10870 14968 10876 14980
rect 10928 14968 10934 15020
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11296 14980 11805 15008
rect 11296 14968 11302 14980
rect 11793 14977 11805 14980
rect 11839 15008 11851 15011
rect 12894 15008 12900 15020
rect 11839 14980 12900 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 14826 14968 14832 15020
rect 14884 15008 14890 15020
rect 15657 15011 15715 15017
rect 15657 15008 15669 15011
rect 14884 14980 15669 15008
rect 14884 14968 14890 14980
rect 15657 14977 15669 14980
rect 15703 15008 15715 15011
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 15703 14980 16865 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 17865 15011 17923 15017
rect 17865 14977 17877 15011
rect 17911 15008 17923 15011
rect 18230 15008 18236 15020
rect 17911 14980 18236 15008
rect 17911 14977 17923 14980
rect 17865 14971 17923 14977
rect 18230 14968 18236 14980
rect 18288 15008 18294 15020
rect 19337 15011 19395 15017
rect 18288 14980 19288 15008
rect 18288 14968 18294 14980
rect 5077 14943 5135 14949
rect 5077 14940 5089 14943
rect 4586 14912 5089 14940
rect 5077 14909 5089 14912
rect 5123 14909 5135 14943
rect 5077 14903 5135 14909
rect 6273 14943 6331 14949
rect 6273 14909 6285 14943
rect 6319 14940 6331 14943
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6319 14912 6837 14940
rect 6319 14909 6331 14912
rect 6273 14903 6331 14909
rect 6825 14909 6837 14912
rect 6871 14940 6883 14943
rect 6914 14940 6920 14952
rect 6871 14912 6920 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14940 12587 14943
rect 12710 14940 12716 14952
rect 12575 14912 12716 14940
rect 12575 14909 12587 14912
rect 12529 14903 12587 14909
rect 12710 14900 12716 14912
rect 12768 14940 12774 14952
rect 13630 14940 13636 14952
rect 12768 14912 13636 14940
rect 12768 14900 12774 14912
rect 13630 14900 13636 14912
rect 13688 14900 13694 14952
rect 19260 14949 19288 14980
rect 19337 14977 19349 15011
rect 19383 15008 19395 15011
rect 19426 15008 19432 15020
rect 19383 14980 19432 15008
rect 19383 14977 19395 14980
rect 19337 14971 19395 14977
rect 19426 14968 19432 14980
rect 19484 14968 19490 15020
rect 20254 14968 20260 15020
rect 20312 15008 20318 15020
rect 20533 15011 20591 15017
rect 20533 15008 20545 15011
rect 20312 14980 20545 15008
rect 20312 14968 20318 14980
rect 20533 14977 20545 14980
rect 20579 14977 20591 15011
rect 21192 15008 21220 15039
rect 23474 15036 23480 15088
rect 23532 15076 23538 15088
rect 23842 15076 23848 15088
rect 23532 15048 23848 15076
rect 23532 15036 23538 15048
rect 23842 15036 23848 15048
rect 23900 15076 23906 15088
rect 23900 15048 24072 15076
rect 23900 15036 23906 15048
rect 21729 15011 21787 15017
rect 21729 15008 21741 15011
rect 21192 14980 21741 15008
rect 20533 14971 20591 14977
rect 21729 14977 21741 14980
rect 21775 14977 21787 15011
rect 21729 14971 21787 14977
rect 23753 15011 23811 15017
rect 23753 14977 23765 15011
rect 23799 15008 23811 15011
rect 23934 15008 23940 15020
rect 23799 14980 23940 15008
rect 23799 14977 23811 14980
rect 23753 14971 23811 14977
rect 23934 14968 23940 14980
rect 23992 14968 23998 15020
rect 24044 15017 24072 15048
rect 24029 15011 24087 15017
rect 24029 14977 24041 15011
rect 24075 14977 24087 15011
rect 24762 15008 24768 15020
rect 24675 14980 24768 15008
rect 24029 14971 24087 14977
rect 24762 14968 24768 14980
rect 24820 15008 24826 15020
rect 27614 15008 27620 15020
rect 24820 14980 27620 15008
rect 24820 14968 24826 14980
rect 27614 14968 27620 14980
rect 27672 14968 27678 15020
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 13786 14912 14289 14940
rect 3016 14844 3648 14872
rect 3697 14875 3755 14881
rect 3016 14832 3022 14844
rect 3697 14841 3709 14875
rect 3743 14872 3755 14875
rect 4062 14872 4068 14884
rect 3743 14844 4068 14872
rect 3743 14841 3755 14844
rect 3697 14835 3755 14841
rect 2317 14807 2375 14813
rect 2317 14773 2329 14807
rect 2363 14804 2375 14807
rect 2406 14804 2412 14816
rect 2363 14776 2412 14804
rect 2363 14773 2375 14776
rect 2317 14767 2375 14773
rect 2406 14764 2412 14776
rect 2464 14764 2470 14816
rect 2498 14764 2504 14816
rect 2556 14804 2562 14816
rect 3712 14804 3740 14835
rect 4062 14832 4068 14844
rect 4120 14832 4126 14884
rect 4246 14832 4252 14884
rect 4304 14872 4310 14884
rect 4304 14844 4654 14872
rect 4304 14832 4310 14844
rect 4522 14804 4528 14816
rect 2556 14776 3740 14804
rect 4483 14776 4528 14804
rect 2556 14764 2562 14776
rect 4522 14764 4528 14776
rect 4580 14764 4586 14816
rect 4626 14804 4654 14844
rect 6454 14832 6460 14884
rect 6512 14872 6518 14884
rect 6641 14875 6699 14881
rect 6641 14872 6653 14875
rect 6512 14844 6653 14872
rect 6512 14832 6518 14844
rect 6641 14841 6653 14844
rect 6687 14872 6699 14875
rect 7187 14875 7245 14881
rect 7187 14872 7199 14875
rect 6687 14844 7199 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 7187 14841 7199 14844
rect 7233 14872 7245 14875
rect 8849 14875 8907 14881
rect 8849 14872 8861 14875
rect 7233 14844 8861 14872
rect 7233 14841 7245 14844
rect 7187 14835 7245 14841
rect 8849 14841 8861 14844
rect 8895 14872 8907 14875
rect 9303 14875 9361 14881
rect 9303 14872 9315 14875
rect 8895 14844 9315 14872
rect 8895 14841 8907 14844
rect 8849 14835 8907 14841
rect 9303 14841 9315 14844
rect 9349 14872 9361 14875
rect 9858 14872 9864 14884
rect 9349 14844 9864 14872
rect 9349 14841 9361 14844
rect 9303 14835 9361 14841
rect 9858 14832 9864 14844
rect 9916 14832 9922 14884
rect 10873 14875 10931 14881
rect 10873 14841 10885 14875
rect 10919 14841 10931 14875
rect 10873 14835 10931 14841
rect 12437 14875 12495 14881
rect 12437 14841 12449 14875
rect 12483 14872 12495 14875
rect 12850 14875 12908 14881
rect 12850 14872 12862 14875
rect 12483 14844 12862 14872
rect 12483 14841 12495 14844
rect 12437 14835 12495 14841
rect 12850 14841 12862 14844
rect 12896 14841 12908 14875
rect 12850 14835 12908 14841
rect 10505 14807 10563 14813
rect 10505 14804 10517 14807
rect 4626 14776 10517 14804
rect 10505 14773 10517 14776
rect 10551 14804 10563 14807
rect 10686 14804 10692 14816
rect 10551 14776 10692 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 10686 14764 10692 14776
rect 10744 14804 10750 14816
rect 10888 14804 10916 14835
rect 13446 14832 13452 14884
rect 13504 14872 13510 14884
rect 13786 14872 13814 14912
rect 14277 14909 14289 14912
rect 14323 14940 14335 14943
rect 14737 14943 14795 14949
rect 14737 14940 14749 14943
rect 14323 14912 14749 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 14737 14909 14749 14912
rect 14783 14909 14795 14943
rect 14737 14903 14795 14909
rect 18376 14943 18434 14949
rect 18376 14909 18388 14943
rect 18422 14909 18434 14943
rect 18376 14903 18434 14909
rect 19245 14943 19303 14949
rect 19245 14909 19257 14943
rect 19291 14940 19303 14943
rect 19291 14912 19564 14940
rect 19291 14909 19303 14912
rect 19245 14903 19303 14909
rect 13504 14844 13814 14872
rect 15197 14875 15255 14881
rect 13504 14832 13510 14844
rect 15197 14841 15209 14875
rect 15243 14872 15255 14875
rect 15565 14875 15623 14881
rect 15565 14872 15577 14875
rect 15243 14844 15577 14872
rect 15243 14841 15255 14844
rect 15197 14835 15255 14841
rect 15565 14841 15577 14844
rect 15611 14872 15623 14875
rect 16019 14875 16077 14881
rect 16019 14872 16031 14875
rect 15611 14844 16031 14872
rect 15611 14841 15623 14844
rect 15565 14835 15623 14841
rect 16019 14841 16031 14844
rect 16065 14872 16077 14875
rect 16114 14872 16120 14884
rect 16065 14844 16120 14872
rect 16065 14841 16077 14844
rect 16019 14835 16077 14841
rect 16114 14832 16120 14844
rect 16172 14832 16178 14884
rect 10744 14776 10916 14804
rect 14461 14807 14519 14813
rect 10744 14764 10750 14776
rect 14461 14773 14473 14807
rect 14507 14804 14519 14807
rect 14550 14804 14556 14816
rect 14507 14776 14556 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 16574 14804 16580 14816
rect 16487 14776 16580 14804
rect 16574 14764 16580 14776
rect 16632 14804 16638 14816
rect 17678 14804 17684 14816
rect 16632 14776 17684 14804
rect 16632 14764 16638 14776
rect 17678 14764 17684 14776
rect 17736 14764 17742 14816
rect 18391 14804 18419 14903
rect 18463 14875 18521 14881
rect 18463 14841 18475 14875
rect 18509 14872 18521 14875
rect 19426 14872 19432 14884
rect 18509 14844 19432 14872
rect 18509 14841 18521 14844
rect 18463 14835 18521 14841
rect 19426 14832 19432 14844
rect 19484 14832 19490 14884
rect 19536 14872 19564 14912
rect 22830 14900 22836 14952
rect 22888 14940 22894 14952
rect 23385 14943 23443 14949
rect 23385 14940 23397 14943
rect 22888 14912 23397 14940
rect 22888 14900 22894 14912
rect 23385 14909 23397 14912
rect 23431 14940 23443 14943
rect 25276 14943 25334 14949
rect 23431 14912 23520 14940
rect 23431 14909 23443 14912
rect 23385 14903 23443 14909
rect 19699 14875 19757 14881
rect 19699 14872 19711 14875
rect 19536 14844 19711 14872
rect 19699 14841 19711 14844
rect 19745 14872 19757 14875
rect 20070 14872 20076 14884
rect 19745 14844 20076 14872
rect 19745 14841 19757 14844
rect 19699 14835 19757 14841
rect 20070 14832 20076 14844
rect 20128 14872 20134 14884
rect 23492 14872 23520 14912
rect 25276 14909 25288 14943
rect 25322 14940 25334 14943
rect 25322 14912 25820 14940
rect 25322 14909 25334 14912
rect 25276 14903 25334 14909
rect 23845 14875 23903 14881
rect 23845 14872 23857 14875
rect 20128 14844 21680 14872
rect 23492 14844 23857 14872
rect 20128 14832 20134 14844
rect 18877 14807 18935 14813
rect 18877 14804 18889 14807
rect 18391 14776 18889 14804
rect 18877 14773 18889 14776
rect 18923 14804 18935 14807
rect 20714 14804 20720 14816
rect 18923 14776 20720 14804
rect 18923 14773 18935 14776
rect 18877 14767 18935 14773
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 21652 14813 21680 14844
rect 23845 14841 23857 14844
rect 23891 14841 23903 14875
rect 23845 14835 23903 14841
rect 24486 14832 24492 14884
rect 24544 14872 24550 14884
rect 25363 14875 25421 14881
rect 25363 14872 25375 14875
rect 24544 14844 25375 14872
rect 24544 14832 24550 14844
rect 25363 14841 25375 14844
rect 25409 14841 25421 14875
rect 25363 14835 25421 14841
rect 25792 14816 25820 14912
rect 21637 14807 21695 14813
rect 21637 14773 21649 14807
rect 21683 14804 21695 14807
rect 22097 14807 22155 14813
rect 22097 14804 22109 14807
rect 21683 14776 22109 14804
rect 21683 14773 21695 14776
rect 21637 14767 21695 14773
rect 22097 14773 22109 14776
rect 22143 14773 22155 14807
rect 25774 14804 25780 14816
rect 25735 14776 25780 14804
rect 22097 14767 22155 14773
rect 25774 14764 25780 14776
rect 25832 14764 25838 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2958 14600 2964 14612
rect 2919 14572 2964 14600
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 3510 14600 3516 14612
rect 3471 14572 3516 14600
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 4522 14600 4528 14612
rect 4483 14572 4528 14600
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 6454 14600 6460 14612
rect 6415 14572 6460 14600
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 7282 14560 7288 14612
rect 7340 14600 7346 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 7340 14572 7665 14600
rect 7340 14560 7346 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 7653 14563 7711 14569
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 7800 14572 8064 14600
rect 7800 14560 7806 14572
rect 1762 14492 1768 14544
rect 1820 14532 1826 14544
rect 2038 14532 2044 14544
rect 1820 14504 2044 14532
rect 1820 14492 1826 14504
rect 2038 14492 2044 14504
rect 2096 14492 2102 14544
rect 2593 14535 2651 14541
rect 2593 14501 2605 14535
rect 2639 14532 2651 14535
rect 2682 14532 2688 14544
rect 2639 14504 2688 14532
rect 2639 14501 2651 14504
rect 2593 14495 2651 14501
rect 2682 14492 2688 14504
rect 2740 14492 2746 14544
rect 7190 14492 7196 14544
rect 7248 14532 7254 14544
rect 7926 14532 7932 14544
rect 7248 14504 7932 14532
rect 7248 14492 7254 14504
rect 7926 14492 7932 14504
rect 7984 14492 7990 14544
rect 8036 14541 8064 14572
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 8904 14572 8953 14600
rect 8904 14560 8910 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 8941 14563 8999 14569
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 10686 14600 10692 14612
rect 10643 14572 10692 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 10870 14600 10876 14612
rect 10831 14572 10876 14600
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 13078 14600 13084 14612
rect 13039 14572 13084 14600
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 13630 14600 13636 14612
rect 13591 14572 13636 14600
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 18782 14560 18788 14612
rect 18840 14600 18846 14612
rect 18969 14603 19027 14609
rect 18969 14600 18981 14603
rect 18840 14572 18981 14600
rect 18840 14560 18846 14572
rect 18969 14569 18981 14572
rect 19015 14569 19027 14603
rect 19978 14600 19984 14612
rect 19939 14572 19984 14600
rect 18969 14563 19027 14569
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20622 14600 20628 14612
rect 20583 14572 20628 14600
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 22278 14600 22284 14612
rect 21008 14572 22284 14600
rect 8021 14535 8079 14541
rect 8021 14501 8033 14535
rect 8067 14501 8079 14535
rect 8021 14495 8079 14501
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 10039 14535 10097 14541
rect 10039 14532 10051 14535
rect 9916 14504 10051 14532
rect 9916 14492 9922 14504
rect 10039 14501 10051 14504
rect 10085 14532 10097 14535
rect 11882 14532 11888 14544
rect 10085 14504 11888 14532
rect 10085 14501 10097 14504
rect 10039 14495 10097 14501
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 12158 14532 12164 14544
rect 12119 14504 12164 14532
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 15927 14535 15985 14541
rect 15927 14501 15939 14535
rect 15973 14532 15985 14535
rect 16114 14532 16120 14544
rect 15973 14504 16120 14532
rect 15973 14501 15985 14504
rect 15927 14495 15985 14501
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 16666 14492 16672 14544
rect 16724 14532 16730 14544
rect 17402 14532 17408 14544
rect 16724 14504 17408 14532
rect 16724 14492 16730 14504
rect 17402 14492 17408 14504
rect 17460 14532 17466 14544
rect 17497 14535 17555 14541
rect 17497 14532 17509 14535
rect 17460 14504 17509 14532
rect 17460 14492 17466 14504
rect 17497 14501 17509 14504
rect 17543 14501 17555 14535
rect 17497 14495 17555 14501
rect 17678 14492 17684 14544
rect 17736 14532 17742 14544
rect 20162 14532 20168 14544
rect 17736 14504 20168 14532
rect 17736 14492 17742 14504
rect 20162 14492 20168 14504
rect 20220 14492 20226 14544
rect 21008 14541 21036 14572
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 20993 14535 21051 14541
rect 20993 14501 21005 14535
rect 21039 14501 21051 14535
rect 20993 14495 21051 14501
rect 21082 14492 21088 14544
rect 21140 14532 21146 14544
rect 21140 14504 21185 14532
rect 21140 14492 21146 14504
rect 22922 14492 22928 14544
rect 22980 14532 22986 14544
rect 23293 14535 23351 14541
rect 23293 14532 23305 14535
rect 22980 14504 23305 14532
rect 22980 14492 22986 14504
rect 23293 14501 23305 14504
rect 23339 14501 23351 14535
rect 23842 14532 23848 14544
rect 23803 14504 23848 14532
rect 23293 14495 23351 14501
rect 23842 14492 23848 14504
rect 23900 14492 23906 14544
rect 24854 14532 24860 14544
rect 24815 14504 24860 14532
rect 24854 14492 24860 14504
rect 24912 14492 24918 14544
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14464 4215 14467
rect 4338 14464 4344 14476
rect 4203 14436 4344 14464
rect 4203 14433 4215 14436
rect 4157 14427 4215 14433
rect 4338 14424 4344 14436
rect 4396 14424 4402 14476
rect 5442 14424 5448 14476
rect 5500 14464 5506 14476
rect 7009 14467 7067 14473
rect 7009 14464 7021 14467
rect 5500 14436 7021 14464
rect 5500 14424 5506 14436
rect 7009 14433 7021 14436
rect 7055 14464 7067 14467
rect 7742 14464 7748 14476
rect 7055 14436 7748 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 13998 14464 14004 14476
rect 13872 14436 13917 14464
rect 13959 14436 14004 14464
rect 13872 14424 13878 14436
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 15286 14424 15292 14476
rect 15344 14464 15350 14476
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 15344 14436 15577 14464
rect 15344 14424 15350 14436
rect 15565 14433 15577 14436
rect 15611 14433 15623 14467
rect 18874 14464 18880 14476
rect 18835 14436 18880 14464
rect 15565 14427 15623 14433
rect 18874 14424 18880 14436
rect 18932 14424 18938 14476
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 19337 14467 19395 14473
rect 19337 14464 19349 14467
rect 19300 14436 19349 14464
rect 19300 14424 19306 14436
rect 19337 14433 19349 14436
rect 19383 14433 19395 14467
rect 19337 14427 19395 14433
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 1949 14399 2007 14405
rect 1949 14396 1961 14399
rect 1811 14368 1961 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 1949 14365 1961 14368
rect 1995 14396 2007 14399
rect 2038 14396 2044 14408
rect 1995 14368 2044 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 6086 14396 6092 14408
rect 6047 14368 6092 14396
rect 6086 14356 6092 14368
rect 6144 14356 6150 14408
rect 8202 14396 8208 14408
rect 8163 14368 8208 14396
rect 8202 14356 8208 14368
rect 8260 14396 8266 14408
rect 9401 14399 9459 14405
rect 9401 14396 9413 14399
rect 8260 14368 9413 14396
rect 8260 14356 8266 14368
rect 9401 14365 9413 14368
rect 9447 14365 9459 14399
rect 9674 14396 9680 14408
rect 9635 14368 9680 14396
rect 9401 14359 9459 14365
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 12342 14396 12348 14408
rect 12115 14368 12348 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 12710 14396 12716 14408
rect 12671 14368 12716 14396
rect 12710 14356 12716 14368
rect 12768 14396 12774 14408
rect 13354 14396 13360 14408
rect 12768 14368 13360 14396
rect 12768 14356 12774 14368
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 17405 14399 17463 14405
rect 17405 14396 17417 14399
rect 17092 14368 17417 14396
rect 17092 14356 17098 14368
rect 17405 14365 17417 14368
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 17681 14399 17739 14405
rect 17681 14396 17693 14399
rect 17644 14368 17693 14396
rect 17644 14356 17650 14368
rect 17681 14365 17693 14368
rect 17727 14365 17739 14399
rect 21358 14396 21364 14408
rect 21319 14368 21364 14396
rect 17681 14359 17739 14365
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 23017 14399 23075 14405
rect 23017 14365 23029 14399
rect 23063 14396 23075 14399
rect 23201 14399 23259 14405
rect 23201 14396 23213 14399
rect 23063 14368 23213 14396
rect 23063 14365 23075 14368
rect 23017 14359 23075 14365
rect 23201 14365 23213 14368
rect 23247 14396 23259 14399
rect 24486 14396 24492 14408
rect 23247 14368 24492 14396
rect 23247 14365 23259 14368
rect 23201 14359 23259 14365
rect 24486 14356 24492 14368
rect 24544 14356 24550 14408
rect 24762 14396 24768 14408
rect 24723 14368 24768 14396
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 25038 14396 25044 14408
rect 24999 14368 25044 14396
rect 25038 14356 25044 14368
rect 25096 14356 25102 14408
rect 3881 14331 3939 14337
rect 3881 14297 3893 14331
rect 3927 14328 3939 14331
rect 3970 14328 3976 14340
rect 3927 14300 3976 14328
rect 3927 14297 3939 14300
rect 3881 14291 3939 14297
rect 3970 14288 3976 14300
rect 4028 14328 4034 14340
rect 5077 14331 5135 14337
rect 5077 14328 5089 14331
rect 4028 14300 5089 14328
rect 4028 14288 4034 14300
rect 5077 14297 5089 14300
rect 5123 14297 5135 14331
rect 5077 14291 5135 14297
rect 10962 14288 10968 14340
rect 11020 14328 11026 14340
rect 13262 14328 13268 14340
rect 11020 14300 13268 14328
rect 11020 14288 11026 14300
rect 13262 14288 13268 14300
rect 13320 14288 13326 14340
rect 20530 14328 20536 14340
rect 16500 14300 20536 14328
rect 16500 14272 16528 14300
rect 20530 14288 20536 14300
rect 20588 14328 20594 14340
rect 22922 14328 22928 14340
rect 20588 14300 22928 14328
rect 20588 14288 20594 14300
rect 22922 14288 22928 14300
rect 22980 14288 22986 14340
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 5534 14260 5540 14272
rect 4120 14232 5540 14260
rect 4120 14220 4126 14232
rect 5534 14220 5540 14232
rect 5592 14260 5598 14272
rect 5629 14263 5687 14269
rect 5629 14260 5641 14263
rect 5592 14232 5641 14260
rect 5592 14220 5598 14232
rect 5629 14229 5641 14232
rect 5675 14229 5687 14263
rect 7282 14260 7288 14272
rect 7243 14232 7288 14260
rect 5629 14223 5687 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 11054 14220 11060 14272
rect 11112 14260 11118 14272
rect 11241 14263 11299 14269
rect 11241 14260 11253 14263
rect 11112 14232 11253 14260
rect 11112 14220 11118 14232
rect 11241 14229 11253 14232
rect 11287 14229 11299 14263
rect 16482 14260 16488 14272
rect 16443 14232 16488 14260
rect 11241 14223 11299 14229
rect 16482 14220 16488 14232
rect 16540 14220 16546 14272
rect 16850 14220 16856 14272
rect 16908 14260 16914 14272
rect 17862 14260 17868 14272
rect 16908 14232 17868 14260
rect 16908 14220 16914 14232
rect 17862 14220 17868 14232
rect 17920 14260 17926 14272
rect 18325 14263 18383 14269
rect 18325 14260 18337 14263
rect 17920 14232 18337 14260
rect 17920 14220 17926 14232
rect 18325 14229 18337 14232
rect 18371 14229 18383 14263
rect 22646 14260 22652 14272
rect 22559 14232 22652 14260
rect 18325 14223 18383 14229
rect 22646 14220 22652 14232
rect 22704 14260 22710 14272
rect 23290 14260 23296 14272
rect 22704 14232 23296 14260
rect 22704 14220 22710 14232
rect 23290 14220 23296 14232
rect 23348 14220 23354 14272
rect 23842 14220 23848 14272
rect 23900 14260 23906 14272
rect 24213 14263 24271 14269
rect 24213 14260 24225 14263
rect 23900 14232 24225 14260
rect 23900 14220 23906 14232
rect 24213 14229 24225 14232
rect 24259 14260 24271 14263
rect 24946 14260 24952 14272
rect 24259 14232 24952 14260
rect 24259 14229 24271 14232
rect 24213 14223 24271 14229
rect 24946 14220 24952 14232
rect 25004 14220 25010 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1762 14056 1768 14068
rect 1723 14028 1768 14056
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 7800 14028 7849 14056
rect 7800 14016 7806 14028
rect 7837 14025 7849 14028
rect 7883 14025 7895 14059
rect 7837 14019 7895 14025
rect 8018 14016 8024 14068
rect 8076 14056 8082 14068
rect 8573 14059 8631 14065
rect 8573 14056 8585 14059
rect 8076 14028 8585 14056
rect 8076 14016 8082 14028
rect 8573 14025 8585 14028
rect 8619 14025 8631 14059
rect 9858 14056 9864 14068
rect 9819 14028 9864 14056
rect 8573 14019 8631 14025
rect 2869 13991 2927 13997
rect 2869 13988 2881 13991
rect 1780 13960 2881 13988
rect 1670 13744 1676 13796
rect 1728 13784 1734 13796
rect 1780 13784 1808 13960
rect 2869 13957 2881 13960
rect 2915 13957 2927 13991
rect 5994 13988 6000 14000
rect 2869 13951 2927 13957
rect 5787 13960 6000 13988
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 3510 13920 3516 13932
rect 2639 13892 3516 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 3510 13880 3516 13892
rect 3568 13920 3574 13932
rect 3789 13923 3847 13929
rect 3789 13920 3801 13923
rect 3568 13892 3801 13920
rect 3568 13880 3574 13892
rect 3789 13889 3801 13892
rect 3835 13889 3847 13923
rect 5787 13920 5815 13960
rect 5994 13948 6000 13960
rect 6052 13988 6058 14000
rect 6270 13988 6276 14000
rect 6052 13960 6276 13988
rect 6052 13948 6058 13960
rect 6270 13948 6276 13960
rect 6328 13948 6334 14000
rect 8588 13988 8616 14019
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 11885 14059 11943 14065
rect 11885 14025 11897 14059
rect 11931 14056 11943 14059
rect 12158 14056 12164 14068
rect 11931 14028 12164 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 15841 14059 15899 14065
rect 15841 14025 15853 14059
rect 15887 14056 15899 14059
rect 16114 14056 16120 14068
rect 15887 14028 16120 14056
rect 15887 14025 15899 14028
rect 15841 14019 15899 14025
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 17034 14016 17040 14068
rect 17092 14056 17098 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 17092 14028 17693 14056
rect 17092 14016 17098 14028
rect 17681 14025 17693 14028
rect 17727 14025 17739 14059
rect 18874 14056 18880 14068
rect 18835 14028 18880 14056
rect 17681 14019 17739 14025
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14056 20131 14059
rect 21082 14056 21088 14068
rect 20119 14028 21088 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 21082 14016 21088 14028
rect 21140 14056 21146 14068
rect 21821 14059 21879 14065
rect 21140 14028 21772 14056
rect 21140 14016 21146 14028
rect 13541 13991 13599 13997
rect 13541 13988 13553 13991
rect 8588 13960 8708 13988
rect 3789 13883 3847 13889
rect 5368 13892 5815 13920
rect 5905 13923 5963 13929
rect 5368 13861 5396 13892
rect 5905 13889 5917 13923
rect 5951 13920 5963 13923
rect 6086 13920 6092 13932
rect 5951 13892 6092 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 6086 13880 6092 13892
rect 6144 13880 6150 13932
rect 5077 13855 5135 13861
rect 2792 13824 2912 13852
rect 1949 13787 2007 13793
rect 1949 13784 1961 13787
rect 1728 13756 1961 13784
rect 1728 13744 1734 13756
rect 1949 13753 1961 13756
rect 1995 13753 2007 13787
rect 1949 13747 2007 13753
rect 2041 13787 2099 13793
rect 2041 13753 2053 13787
rect 2087 13784 2099 13787
rect 2130 13784 2136 13796
rect 2087 13756 2136 13784
rect 2087 13753 2099 13756
rect 2041 13747 2099 13753
rect 2130 13744 2136 13756
rect 2188 13784 2194 13796
rect 2590 13784 2596 13796
rect 2188 13756 2596 13784
rect 2188 13744 2194 13756
rect 2590 13744 2596 13756
rect 2648 13744 2654 13796
rect 1486 13676 1492 13728
rect 1544 13716 1550 13728
rect 2792 13716 2820 13824
rect 2884 13784 2912 13824
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5353 13855 5411 13861
rect 5353 13852 5365 13855
rect 5123 13824 5365 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5353 13821 5365 13824
rect 5399 13821 5411 13855
rect 5353 13815 5411 13821
rect 5629 13855 5687 13861
rect 5629 13821 5641 13855
rect 5675 13821 5687 13855
rect 5629 13815 5687 13821
rect 3510 13784 3516 13796
rect 2884 13756 3516 13784
rect 3510 13744 3516 13756
rect 3568 13744 3574 13796
rect 3605 13787 3663 13793
rect 3605 13753 3617 13787
rect 3651 13753 3663 13787
rect 3605 13747 3663 13753
rect 1544 13688 2820 13716
rect 3329 13719 3387 13725
rect 1544 13676 1550 13688
rect 3329 13685 3341 13719
rect 3375 13716 3387 13719
rect 3418 13716 3424 13728
rect 3375 13688 3424 13716
rect 3375 13685 3387 13688
rect 3329 13679 3387 13685
rect 3418 13676 3424 13688
rect 3476 13716 3482 13728
rect 3620 13716 3648 13747
rect 5166 13744 5172 13796
rect 5224 13784 5230 13796
rect 5644 13784 5672 13815
rect 6362 13812 6368 13864
rect 6420 13852 6426 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6420 13824 6837 13852
rect 6420 13812 6426 13824
rect 6825 13821 6837 13824
rect 6871 13852 6883 13855
rect 7098 13852 7104 13864
rect 6871 13824 7104 13852
rect 6871 13821 6883 13824
rect 6825 13815 6883 13821
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 8205 13855 8263 13861
rect 8205 13852 8217 13855
rect 7340 13824 8217 13852
rect 7340 13812 7346 13824
rect 8205 13821 8217 13824
rect 8251 13852 8263 13855
rect 8570 13852 8576 13864
rect 8251 13824 8576 13852
rect 8251 13821 8263 13824
rect 8205 13815 8263 13821
rect 8570 13812 8576 13824
rect 8628 13812 8634 13864
rect 8680 13852 8708 13960
rect 11256 13960 13553 13988
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13920 9551 13923
rect 9674 13920 9680 13932
rect 9539 13892 9680 13920
rect 9539 13889 9551 13892
rect 9493 13883 9551 13889
rect 9674 13880 9680 13892
rect 9732 13920 9738 13932
rect 10137 13923 10195 13929
rect 10137 13920 10149 13923
rect 9732 13892 10149 13920
rect 9732 13880 9738 13892
rect 10137 13889 10149 13892
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 8757 13855 8815 13861
rect 8757 13852 8769 13855
rect 8680 13824 8769 13852
rect 8757 13821 8769 13824
rect 8803 13821 8815 13855
rect 8757 13815 8815 13821
rect 7300 13784 7328 13812
rect 5224 13756 7328 13784
rect 8772 13784 8800 13815
rect 8846 13812 8852 13864
rect 8904 13852 8910 13864
rect 9217 13855 9275 13861
rect 9217 13852 9229 13855
rect 8904 13824 9229 13852
rect 8904 13812 8910 13824
rect 9217 13821 9229 13824
rect 9263 13821 9275 13855
rect 9217 13815 9275 13821
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13852 9643 13855
rect 10689 13855 10747 13861
rect 10689 13852 10701 13855
rect 9631 13824 10701 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 10689 13821 10701 13824
rect 10735 13852 10747 13855
rect 10962 13852 10968 13864
rect 10735 13824 10968 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11256 13861 11284 13960
rect 13541 13957 13553 13960
rect 13587 13988 13599 13991
rect 13998 13988 14004 14000
rect 13587 13960 14004 13988
rect 13587 13957 13599 13960
rect 13541 13951 13599 13957
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 14734 13948 14740 14000
rect 14792 13988 14798 14000
rect 17494 13988 17500 14000
rect 14792 13960 17500 13988
rect 14792 13948 14798 13960
rect 17494 13948 17500 13960
rect 17552 13988 17558 14000
rect 18233 13991 18291 13997
rect 18233 13988 18245 13991
rect 17552 13960 18245 13988
rect 17552 13948 17558 13960
rect 18233 13957 18245 13960
rect 18279 13957 18291 13991
rect 19978 13988 19984 14000
rect 18233 13951 18291 13957
rect 19260 13960 19984 13988
rect 12802 13920 12808 13932
rect 12763 13892 12808 13920
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 15473 13923 15531 13929
rect 15473 13889 15485 13923
rect 15519 13920 15531 13923
rect 16850 13920 16856 13932
rect 15519 13892 16856 13920
rect 15519 13889 15531 13892
rect 15473 13883 15531 13889
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17586 13920 17592 13932
rect 17083 13892 17592 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17586 13880 17592 13892
rect 17644 13880 17650 13932
rect 19260 13929 19288 13960
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 20162 13948 20168 14000
rect 20220 13988 20226 14000
rect 20625 13991 20683 13997
rect 20625 13988 20637 13991
rect 20220 13960 20637 13988
rect 20220 13948 20226 13960
rect 20625 13957 20637 13960
rect 20671 13988 20683 13991
rect 20898 13988 20904 14000
rect 20671 13960 20904 13988
rect 20671 13957 20683 13960
rect 20625 13951 20683 13957
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 21358 13988 21364 14000
rect 21319 13960 21364 13988
rect 21358 13948 21364 13960
rect 21416 13948 21422 14000
rect 21744 13988 21772 14028
rect 21821 14025 21833 14059
rect 21867 14056 21879 14059
rect 22278 14056 22284 14068
rect 21867 14028 22284 14056
rect 21867 14025 21879 14028
rect 21821 14019 21879 14025
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 22695 14059 22753 14065
rect 22695 14025 22707 14059
rect 22741 14056 22753 14059
rect 24118 14056 24124 14068
rect 22741 14028 24124 14056
rect 22741 14025 22753 14028
rect 22695 14019 22753 14025
rect 24118 14016 24124 14028
rect 24176 14016 24182 14068
rect 24765 14059 24823 14065
rect 24765 14025 24777 14059
rect 24811 14056 24823 14059
rect 24854 14056 24860 14068
rect 24811 14028 24860 14056
rect 24811 14025 24823 14028
rect 24765 14019 24823 14025
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 24946 14016 24952 14068
rect 25004 14056 25010 14068
rect 25363 14059 25421 14065
rect 25363 14056 25375 14059
rect 25004 14028 25375 14056
rect 25004 14016 25010 14028
rect 25363 14025 25375 14028
rect 25409 14025 25421 14059
rect 25363 14019 25421 14025
rect 22097 13991 22155 13997
rect 22097 13988 22109 13991
rect 21744 13960 22109 13988
rect 22097 13957 22109 13960
rect 22143 13988 22155 13991
rect 22830 13988 22836 14000
rect 22143 13960 22836 13988
rect 22143 13957 22155 13960
rect 22097 13951 22155 13957
rect 22830 13948 22836 13960
rect 22888 13948 22894 14000
rect 22922 13948 22928 14000
rect 22980 13988 22986 14000
rect 23017 13991 23075 13997
rect 23017 13988 23029 13991
rect 22980 13960 23029 13988
rect 22980 13948 22986 13960
rect 23017 13957 23029 13960
rect 23063 13957 23075 13991
rect 23017 13951 23075 13957
rect 19245 13923 19303 13929
rect 19245 13889 19257 13923
rect 19291 13889 19303 13923
rect 19245 13883 19303 13889
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 20438 13920 20444 13932
rect 19484 13892 20444 13920
rect 19484 13880 19490 13892
rect 20438 13880 20444 13892
rect 20496 13920 20502 13932
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 20496 13892 20821 13920
rect 20496 13880 20502 13892
rect 20809 13889 20821 13892
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 23753 13923 23811 13929
rect 23753 13889 23765 13923
rect 23799 13920 23811 13923
rect 23842 13920 23848 13932
rect 23799 13892 23848 13920
rect 23799 13889 23811 13892
rect 23753 13883 23811 13889
rect 23842 13880 23848 13892
rect 23900 13880 23906 13932
rect 23934 13880 23940 13932
rect 23992 13920 23998 13932
rect 24029 13923 24087 13929
rect 24029 13920 24041 13923
rect 23992 13892 24041 13920
rect 23992 13880 23998 13892
rect 24029 13889 24041 13892
rect 24075 13889 24087 13923
rect 24029 13883 24087 13889
rect 24762 13880 24768 13932
rect 24820 13920 24826 13932
rect 25041 13923 25099 13929
rect 25041 13920 25053 13923
rect 24820 13892 25053 13920
rect 24820 13880 24826 13892
rect 25041 13889 25053 13892
rect 25087 13889 25099 13923
rect 25041 13883 25099 13889
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 11112 13824 11253 13852
rect 11112 13812 11118 13824
rect 11241 13821 11253 13824
rect 11287 13821 11299 13855
rect 11241 13815 11299 13821
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 13872 13824 14013 13852
rect 13872 13812 13878 13824
rect 14001 13821 14013 13824
rect 14047 13852 14059 13855
rect 14458 13852 14464 13864
rect 14047 13824 14464 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 14734 13852 14740 13864
rect 14695 13824 14740 13852
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13852 18107 13855
rect 18506 13852 18512 13864
rect 18095 13824 18512 13852
rect 18095 13821 18107 13824
rect 18049 13815 18107 13821
rect 9858 13784 9864 13796
rect 8772 13756 9864 13784
rect 5224 13744 5230 13756
rect 9858 13744 9864 13756
rect 9916 13744 9922 13796
rect 11422 13744 11428 13796
rect 11480 13784 11486 13796
rect 11517 13787 11575 13793
rect 11517 13784 11529 13787
rect 11480 13756 11529 13784
rect 11480 13744 11486 13756
rect 11517 13753 11529 13756
rect 11563 13753 11575 13787
rect 12526 13784 12532 13796
rect 12487 13756 12532 13784
rect 11517 13747 11575 13753
rect 12526 13744 12532 13756
rect 12584 13744 12590 13796
rect 12621 13787 12679 13793
rect 12621 13753 12633 13787
rect 12667 13753 12679 13787
rect 14550 13784 14556 13796
rect 14511 13756 14556 13784
rect 12621 13747 12679 13753
rect 3476 13688 3648 13716
rect 4525 13719 4583 13725
rect 3476 13676 3482 13688
rect 4525 13685 4537 13719
rect 4571 13716 4583 13719
rect 5994 13716 6000 13728
rect 4571 13688 6000 13716
rect 4571 13685 4583 13688
rect 4525 13679 4583 13685
rect 5994 13676 6000 13688
rect 6052 13716 6058 13728
rect 6181 13719 6239 13725
rect 6181 13716 6193 13719
rect 6052 13688 6193 13716
rect 6052 13676 6058 13688
rect 6181 13685 6193 13688
rect 6227 13685 6239 13719
rect 6181 13679 6239 13685
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 6420 13688 6561 13716
rect 6420 13676 6426 13688
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 6914 13716 6920 13728
rect 6875 13688 6920 13716
rect 6549 13679 6607 13685
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 9585 13719 9643 13725
rect 9585 13716 9597 13719
rect 7156 13688 9597 13716
rect 7156 13676 7162 13688
rect 9585 13685 9597 13688
rect 9631 13685 9643 13719
rect 9585 13679 9643 13685
rect 12158 13676 12164 13728
rect 12216 13716 12222 13728
rect 12636 13716 12664 13747
rect 14550 13744 14556 13756
rect 14608 13784 14614 13796
rect 15212 13784 15240 13815
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 19889 13855 19947 13861
rect 19889 13821 19901 13855
rect 19935 13852 19947 13855
rect 20254 13852 20260 13864
rect 19935 13824 20260 13852
rect 19935 13821 19947 13824
rect 19889 13815 19947 13821
rect 20254 13812 20260 13824
rect 20312 13812 20318 13864
rect 22557 13855 22615 13861
rect 22557 13821 22569 13855
rect 22603 13852 22615 13855
rect 22646 13852 22652 13864
rect 22603 13824 22652 13852
rect 22603 13821 22615 13824
rect 22557 13815 22615 13821
rect 22646 13812 22652 13824
rect 22704 13812 22710 13864
rect 25276 13855 25334 13861
rect 25276 13821 25288 13855
rect 25322 13852 25334 13855
rect 25322 13824 25820 13852
rect 25322 13821 25334 13824
rect 25276 13815 25334 13821
rect 25792 13796 25820 13824
rect 16390 13784 16396 13796
rect 14608 13756 15240 13784
rect 16040 13756 16396 13784
rect 14608 13744 14614 13756
rect 12216 13688 12664 13716
rect 12216 13676 12222 13688
rect 14274 13676 14280 13728
rect 14332 13716 14338 13728
rect 16040 13716 16068 13756
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 16482 13744 16488 13796
rect 16540 13784 16546 13796
rect 19337 13787 19395 13793
rect 16540 13756 16585 13784
rect 16540 13744 16546 13756
rect 19337 13753 19349 13787
rect 19383 13784 19395 13787
rect 19702 13784 19708 13796
rect 19383 13756 19708 13784
rect 19383 13753 19395 13756
rect 19337 13747 19395 13753
rect 19702 13744 19708 13756
rect 19760 13744 19766 13796
rect 19978 13744 19984 13796
rect 20036 13784 20042 13796
rect 20165 13787 20223 13793
rect 20165 13784 20177 13787
rect 20036 13756 20177 13784
rect 20036 13744 20042 13756
rect 20165 13753 20177 13756
rect 20211 13753 20223 13787
rect 20898 13784 20904 13796
rect 20859 13756 20904 13784
rect 20165 13747 20223 13753
rect 20898 13744 20904 13756
rect 20956 13784 20962 13796
rect 23385 13787 23443 13793
rect 23385 13784 23397 13787
rect 20956 13756 23397 13784
rect 20956 13744 20962 13756
rect 23385 13753 23397 13756
rect 23431 13784 23443 13787
rect 23845 13787 23903 13793
rect 23845 13784 23857 13787
rect 23431 13756 23857 13784
rect 23431 13753 23443 13756
rect 23385 13747 23443 13753
rect 23845 13753 23857 13756
rect 23891 13753 23903 13787
rect 25774 13784 25780 13796
rect 25687 13756 25780 13784
rect 23845 13747 23903 13753
rect 25774 13744 25780 13756
rect 25832 13744 25838 13796
rect 14332 13688 16068 13716
rect 16209 13719 16267 13725
rect 14332 13676 14338 13688
rect 16209 13685 16221 13719
rect 16255 13716 16267 13719
rect 16500 13716 16528 13744
rect 17402 13716 17408 13728
rect 16255 13688 16528 13716
rect 17315 13688 17408 13716
rect 16255 13685 16267 13688
rect 16209 13679 16267 13685
rect 17402 13676 17408 13688
rect 17460 13716 17466 13728
rect 20073 13719 20131 13725
rect 20073 13716 20085 13719
rect 17460 13688 20085 13716
rect 17460 13676 17466 13688
rect 20073 13685 20085 13688
rect 20119 13685 20131 13719
rect 20073 13679 20131 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 2130 13512 2136 13524
rect 1995 13484 2136 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 2130 13472 2136 13484
rect 2188 13472 2194 13524
rect 3510 13512 3516 13524
rect 3471 13484 3516 13512
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 3881 13515 3939 13521
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 4338 13512 4344 13524
rect 3927 13484 4344 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 4338 13472 4344 13484
rect 4396 13472 4402 13524
rect 5074 13472 5080 13524
rect 5132 13512 5138 13524
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 5132 13484 5181 13512
rect 5132 13472 5138 13484
rect 5169 13481 5181 13484
rect 5215 13481 5227 13515
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 5169 13475 5227 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 7926 13512 7932 13524
rect 7887 13484 7932 13512
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 8018 13472 8024 13524
rect 8076 13512 8082 13524
rect 8076 13484 8248 13512
rect 8076 13472 8082 13484
rect 2409 13447 2467 13453
rect 2409 13413 2421 13447
rect 2455 13444 2467 13447
rect 2498 13444 2504 13456
rect 2455 13416 2504 13444
rect 2455 13413 2467 13416
rect 2409 13407 2467 13413
rect 2498 13404 2504 13416
rect 2556 13404 2562 13456
rect 4246 13444 4252 13456
rect 4207 13416 4252 13444
rect 4246 13404 4252 13416
rect 4304 13404 4310 13456
rect 6638 13444 6644 13456
rect 6599 13416 6644 13444
rect 6638 13404 6644 13416
rect 6696 13404 6702 13456
rect 8220 13453 8248 13484
rect 9398 13472 9404 13524
rect 9456 13512 9462 13524
rect 9769 13515 9827 13521
rect 9769 13512 9781 13515
rect 9456 13484 9781 13512
rect 9456 13472 9462 13484
rect 9769 13481 9781 13484
rect 9815 13481 9827 13515
rect 12158 13512 12164 13524
rect 12119 13484 12164 13512
rect 9769 13475 9827 13481
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 14734 13512 14740 13524
rect 14695 13484 14740 13512
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 15344 13484 16313 13512
rect 15344 13472 15350 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 16390 13472 16396 13524
rect 16448 13512 16454 13524
rect 16669 13515 16727 13521
rect 16669 13512 16681 13515
rect 16448 13484 16681 13512
rect 16448 13472 16454 13484
rect 16669 13481 16681 13484
rect 16715 13481 16727 13515
rect 16669 13475 16727 13481
rect 18969 13515 19027 13521
rect 18969 13481 18981 13515
rect 19015 13512 19027 13515
rect 19242 13512 19248 13524
rect 19015 13484 19248 13512
rect 19015 13481 19027 13484
rect 18969 13475 19027 13481
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 20438 13472 20444 13524
rect 20496 13512 20502 13524
rect 20625 13515 20683 13521
rect 20625 13512 20637 13515
rect 20496 13484 20637 13512
rect 20496 13472 20502 13484
rect 20625 13481 20637 13484
rect 20671 13481 20683 13515
rect 23750 13512 23756 13524
rect 23663 13484 23756 13512
rect 20625 13475 20683 13481
rect 23750 13472 23756 13484
rect 23808 13512 23814 13524
rect 25038 13512 25044 13524
rect 23808 13484 25044 13512
rect 23808 13472 23814 13484
rect 25038 13472 25044 13484
rect 25096 13472 25102 13524
rect 8205 13447 8263 13453
rect 8205 13413 8217 13447
rect 8251 13413 8263 13447
rect 8205 13407 8263 13413
rect 11603 13447 11661 13453
rect 11603 13413 11615 13447
rect 11649 13444 11661 13447
rect 11882 13444 11888 13456
rect 11649 13416 11888 13444
rect 11649 13413 11661 13416
rect 11603 13407 11661 13413
rect 11882 13404 11888 13416
rect 11940 13404 11946 13456
rect 14366 13444 14372 13456
rect 14327 13416 14372 13444
rect 14366 13404 14372 13416
rect 14424 13404 14430 13456
rect 19426 13444 19432 13456
rect 19387 13416 19432 13444
rect 19426 13404 19432 13416
rect 19484 13404 19490 13456
rect 19981 13447 20039 13453
rect 19981 13413 19993 13447
rect 20027 13444 20039 13447
rect 20254 13444 20260 13456
rect 20027 13416 20260 13444
rect 20027 13413 20039 13416
rect 19981 13407 20039 13413
rect 20254 13404 20260 13416
rect 20312 13404 20318 13456
rect 20990 13444 20996 13456
rect 20951 13416 20996 13444
rect 20990 13404 20996 13416
rect 21048 13404 21054 13456
rect 21082 13404 21088 13456
rect 21140 13444 21146 13456
rect 22741 13447 22799 13453
rect 21140 13416 21185 13444
rect 21140 13404 21146 13416
rect 22741 13413 22753 13447
rect 22787 13444 22799 13447
rect 22922 13444 22928 13456
rect 22787 13416 22928 13444
rect 22787 13413 22799 13416
rect 22741 13407 22799 13413
rect 22922 13404 22928 13416
rect 22980 13404 22986 13456
rect 23474 13404 23480 13456
rect 23532 13444 23538 13456
rect 24305 13447 24363 13453
rect 24305 13444 24317 13447
rect 23532 13416 24317 13444
rect 23532 13404 23538 13416
rect 24305 13413 24317 13416
rect 24351 13444 24363 13447
rect 24854 13444 24860 13456
rect 24351 13416 24860 13444
rect 24351 13413 24363 13416
rect 24305 13407 24363 13413
rect 24854 13404 24860 13416
rect 24912 13404 24918 13456
rect 9858 13376 9864 13388
rect 9819 13348 9864 13376
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 10134 13376 10140 13388
rect 10095 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 12342 13376 12348 13388
rect 10657 13348 12348 13376
rect 2130 13268 2136 13320
rect 2188 13308 2194 13320
rect 2317 13311 2375 13317
rect 2317 13308 2329 13311
rect 2188 13280 2329 13308
rect 2188 13268 2194 13280
rect 2317 13277 2329 13280
rect 2363 13277 2375 13311
rect 2958 13308 2964 13320
rect 2919 13280 2964 13308
rect 2317 13271 2375 13277
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 4522 13308 4528 13320
rect 4212 13280 4257 13308
rect 4483 13280 4528 13308
rect 4212 13268 4218 13280
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 5534 13268 5540 13320
rect 5592 13308 5598 13320
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 5592 13280 6561 13308
rect 5592 13268 5598 13280
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 8110 13308 8116 13320
rect 7984 13280 8116 13308
rect 7984 13268 7990 13280
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 8386 13308 8392 13320
rect 8347 13280 8392 13308
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 10657 13308 10685 13348
rect 12342 13336 12348 13348
rect 12400 13376 12406 13388
rect 12437 13379 12495 13385
rect 12437 13376 12449 13379
rect 12400 13348 12449 13376
rect 12400 13336 12406 13348
rect 12437 13345 12449 13348
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13345 13691 13379
rect 13633 13339 13691 13345
rect 9272 13280 10685 13308
rect 11241 13311 11299 13317
rect 9272 13268 9278 13280
rect 11241 13277 11253 13311
rect 11287 13308 11299 13311
rect 11422 13308 11428 13320
rect 11287 13280 11428 13308
rect 11287 13277 11299 13280
rect 11241 13271 11299 13277
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 13648 13308 13676 13339
rect 13722 13336 13728 13388
rect 13780 13376 13786 13388
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 13780 13348 14105 13376
rect 13780 13336 13786 13348
rect 14093 13345 14105 13348
rect 14139 13376 14151 13379
rect 14550 13376 14556 13388
rect 14139 13348 14556 13376
rect 14139 13345 14151 13348
rect 14093 13339 14151 13345
rect 14550 13336 14556 13348
rect 14608 13336 14614 13388
rect 15930 13376 15936 13388
rect 15891 13348 15936 13376
rect 15930 13336 15936 13348
rect 15988 13336 15994 13388
rect 17862 13376 17868 13388
rect 17823 13348 17868 13376
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18141 13379 18199 13385
rect 18141 13345 18153 13379
rect 18187 13345 18199 13379
rect 18141 13339 18199 13345
rect 13998 13308 14004 13320
rect 13648 13280 14004 13308
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 17218 13268 17224 13320
rect 17276 13308 17282 13320
rect 18156 13308 18184 13339
rect 18414 13308 18420 13320
rect 17276 13280 18184 13308
rect 18375 13280 18420 13308
rect 17276 13268 17282 13280
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 19337 13311 19395 13317
rect 19337 13277 19349 13311
rect 19383 13277 19395 13311
rect 20272 13308 20300 13404
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 20272 13280 21281 13308
rect 19337 13271 19395 13277
rect 21269 13277 21281 13280
rect 21315 13308 21327 13311
rect 21913 13311 21971 13317
rect 21913 13308 21925 13311
rect 21315 13280 21925 13308
rect 21315 13277 21327 13280
rect 21269 13271 21327 13277
rect 21913 13277 21925 13280
rect 21959 13308 21971 13311
rect 22002 13308 22008 13320
rect 21959 13280 22008 13308
rect 21959 13277 21971 13280
rect 21913 13271 21971 13277
rect 7101 13243 7159 13249
rect 7101 13209 7113 13243
rect 7147 13240 7159 13243
rect 8404 13240 8432 13268
rect 7147 13212 8432 13240
rect 7147 13209 7159 13212
rect 7101 13203 7159 13209
rect 11330 13200 11336 13252
rect 11388 13240 11394 13252
rect 12526 13240 12532 13252
rect 11388 13212 12532 13240
rect 11388 13200 11394 13212
rect 12526 13200 12532 13212
rect 12584 13240 12590 13252
rect 12805 13243 12863 13249
rect 12805 13240 12817 13243
rect 12584 13212 12817 13240
rect 12584 13200 12590 13212
rect 12805 13209 12817 13212
rect 12851 13209 12863 13243
rect 12805 13203 12863 13209
rect 12986 13200 12992 13252
rect 13044 13240 13050 13252
rect 19352 13240 19380 13271
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 22649 13311 22707 13317
rect 22649 13277 22661 13311
rect 22695 13277 22707 13311
rect 24210 13308 24216 13320
rect 24171 13280 24216 13308
rect 22649 13271 22707 13277
rect 19610 13240 19616 13252
rect 13044 13212 19616 13240
rect 13044 13200 13050 13212
rect 19610 13200 19616 13212
rect 19668 13200 19674 13252
rect 22664 13184 22692 13271
rect 24210 13268 24216 13280
rect 24268 13268 24274 13320
rect 24489 13311 24547 13317
rect 24489 13308 24501 13311
rect 24320 13280 24501 13308
rect 23198 13240 23204 13252
rect 23159 13212 23204 13240
rect 23198 13200 23204 13212
rect 23256 13200 23262 13252
rect 24320 13240 24348 13280
rect 24489 13277 24501 13280
rect 24535 13277 24547 13311
rect 24489 13271 24547 13277
rect 23446 13212 24348 13240
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 7469 13175 7527 13181
rect 7469 13172 7481 13175
rect 6880 13144 7481 13172
rect 6880 13132 6886 13144
rect 7469 13141 7481 13144
rect 7515 13141 7527 13175
rect 7469 13135 7527 13141
rect 10873 13175 10931 13181
rect 10873 13141 10885 13175
rect 10919 13172 10931 13175
rect 11054 13172 11060 13184
rect 10919 13144 11060 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 15562 13172 15568 13184
rect 15523 13144 15568 13172
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 22646 13132 22652 13184
rect 22704 13172 22710 13184
rect 23446 13172 23474 13212
rect 22704 13144 23474 13172
rect 22704 13132 22710 13144
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 4246 12928 4252 12980
rect 4304 12968 4310 12980
rect 4709 12971 4767 12977
rect 4709 12968 4721 12971
rect 4304 12940 4721 12968
rect 4304 12928 4310 12940
rect 4709 12937 4721 12940
rect 4755 12968 4767 12971
rect 5074 12968 5080 12980
rect 4755 12940 5080 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5258 12928 5264 12980
rect 5316 12968 5322 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5316 12940 5917 12968
rect 5316 12928 5322 12940
rect 5905 12937 5917 12940
rect 5951 12937 5963 12971
rect 5905 12931 5963 12937
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 10134 12968 10140 12980
rect 8628 12940 10140 12968
rect 8628 12928 8634 12940
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 11882 12968 11888 12980
rect 11843 12940 11888 12968
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 13722 12968 13728 12980
rect 13683 12940 13728 12968
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 13998 12968 14004 12980
rect 13911 12940 14004 12968
rect 13998 12928 14004 12940
rect 14056 12968 14062 12980
rect 17126 12968 17132 12980
rect 14056 12940 17132 12968
rect 14056 12928 14062 12940
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 17770 12968 17776 12980
rect 17731 12940 17776 12968
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 19610 12968 19616 12980
rect 19571 12940 19616 12968
rect 19610 12928 19616 12940
rect 19668 12928 19674 12980
rect 20070 12968 20076 12980
rect 20031 12940 20076 12968
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 21082 12928 21088 12980
rect 21140 12968 21146 12980
rect 21361 12971 21419 12977
rect 21361 12968 21373 12971
rect 21140 12940 21373 12968
rect 21140 12928 21146 12940
rect 21361 12937 21373 12940
rect 21407 12937 21419 12971
rect 23474 12968 23480 12980
rect 21361 12931 21419 12937
rect 23446 12928 23480 12968
rect 23532 12968 23538 12980
rect 23532 12940 23577 12968
rect 23532 12928 23538 12940
rect 24210 12928 24216 12980
rect 24268 12968 24274 12980
rect 24673 12971 24731 12977
rect 24673 12968 24685 12971
rect 24268 12940 24685 12968
rect 24268 12928 24274 12940
rect 24673 12937 24685 12940
rect 24719 12937 24731 12971
rect 24673 12931 24731 12937
rect 1765 12903 1823 12909
rect 1765 12869 1777 12903
rect 1811 12900 1823 12903
rect 2498 12900 2504 12912
rect 1811 12872 2504 12900
rect 1811 12869 1823 12872
rect 1765 12863 1823 12869
rect 1780 12696 1808 12863
rect 2498 12860 2504 12872
rect 2556 12900 2562 12912
rect 2869 12903 2927 12909
rect 2869 12900 2881 12903
rect 2556 12872 2881 12900
rect 2556 12860 2562 12872
rect 2869 12869 2881 12872
rect 2915 12900 2927 12903
rect 7006 12900 7012 12912
rect 2915 12872 7012 12900
rect 2915 12869 2927 12872
rect 2869 12863 2927 12869
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 9858 12900 9864 12912
rect 9771 12872 9864 12900
rect 9858 12860 9864 12872
rect 9916 12900 9922 12912
rect 10689 12903 10747 12909
rect 10689 12900 10701 12903
rect 9916 12872 10701 12900
rect 9916 12860 9922 12872
rect 10689 12869 10701 12872
rect 10735 12900 10747 12903
rect 14016 12900 14044 12928
rect 10735 12872 14044 12900
rect 10735 12869 10747 12872
rect 10689 12863 10747 12869
rect 1946 12832 1952 12844
rect 1907 12804 1952 12832
rect 1946 12792 1952 12804
rect 2004 12792 2010 12844
rect 2958 12792 2964 12844
rect 3016 12832 3022 12844
rect 3786 12832 3792 12844
rect 3016 12804 3792 12832
rect 3016 12792 3022 12804
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 4154 12792 4160 12844
rect 4212 12832 4218 12844
rect 5077 12835 5135 12841
rect 5077 12832 5089 12835
rect 4212 12804 5089 12832
rect 4212 12792 4218 12804
rect 5077 12801 5089 12804
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12764 5779 12767
rect 6181 12767 6239 12773
rect 6181 12764 6193 12767
rect 5767 12736 6193 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 6181 12733 6193 12736
rect 6227 12764 6239 12767
rect 6730 12764 6736 12776
rect 6227 12736 6736 12764
rect 6227 12733 6239 12736
rect 6181 12727 6239 12733
rect 6730 12724 6736 12736
rect 6788 12724 6794 12776
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12764 7619 12767
rect 8386 12764 8392 12776
rect 7607 12736 8392 12764
rect 7607 12733 7619 12736
rect 7561 12727 7619 12733
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12764 8631 12767
rect 8754 12764 8760 12776
rect 8619 12736 8760 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 10980 12773 11008 12872
rect 14090 12860 14096 12912
rect 14148 12900 14154 12912
rect 16022 12900 16028 12912
rect 14148 12872 16028 12900
rect 14148 12860 14154 12872
rect 16022 12860 16028 12872
rect 16080 12900 16086 12912
rect 16393 12903 16451 12909
rect 16393 12900 16405 12903
rect 16080 12872 16405 12900
rect 16080 12860 16086 12872
rect 16393 12869 16405 12872
rect 16439 12869 16451 12903
rect 16393 12863 16451 12869
rect 19337 12903 19395 12909
rect 19337 12869 19349 12903
rect 19383 12900 19395 12903
rect 19426 12900 19432 12912
rect 19383 12872 19432 12900
rect 19383 12869 19395 12872
rect 19337 12863 19395 12869
rect 19426 12860 19432 12872
rect 19484 12900 19490 12912
rect 23446 12900 23474 12928
rect 19484 12872 23474 12900
rect 19484 12860 19490 12872
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12768 12804 12817 12832
rect 12768 12792 12774 12804
rect 12805 12801 12817 12804
rect 12851 12801 12863 12835
rect 12805 12795 12863 12801
rect 13538 12792 13544 12844
rect 13596 12832 13602 12844
rect 14550 12832 14556 12844
rect 13596 12804 13814 12832
rect 14511 12804 14556 12832
rect 13596 12792 13602 12804
rect 10965 12767 11023 12773
rect 10965 12733 10977 12767
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 11112 12736 11253 12764
rect 11112 12724 11118 12736
rect 11241 12733 11253 12736
rect 11287 12733 11299 12767
rect 11241 12727 11299 12733
rect 2041 12699 2099 12705
rect 2041 12696 2053 12699
rect 1780 12668 2053 12696
rect 2041 12665 2053 12668
rect 2087 12665 2099 12699
rect 2590 12696 2596 12708
rect 2551 12668 2596 12696
rect 2041 12659 2099 12665
rect 2590 12656 2596 12668
rect 2648 12656 2654 12708
rect 3878 12705 3884 12708
rect 3605 12699 3663 12705
rect 3605 12665 3617 12699
rect 3651 12696 3663 12699
rect 3874 12696 3884 12705
rect 3651 12668 3884 12696
rect 3651 12665 3663 12668
rect 3605 12659 3663 12665
rect 3874 12659 3884 12668
rect 3878 12656 3884 12659
rect 3936 12656 3942 12708
rect 4433 12699 4491 12705
rect 4433 12665 4445 12699
rect 4479 12696 4491 12699
rect 4522 12696 4528 12708
rect 4479 12668 4528 12696
rect 4479 12665 4491 12668
rect 4433 12659 4491 12665
rect 4522 12656 4528 12668
rect 4580 12656 4586 12708
rect 6917 12699 6975 12705
rect 6917 12665 6929 12699
rect 6963 12665 6975 12699
rect 6917 12659 6975 12665
rect 5534 12628 5540 12640
rect 5495 12600 5540 12628
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 6638 12628 6644 12640
rect 6599 12600 6644 12628
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 6822 12588 6828 12640
rect 6880 12628 6886 12640
rect 6932 12628 6960 12659
rect 7006 12656 7012 12708
rect 7064 12696 7070 12708
rect 8481 12699 8539 12705
rect 7064 12668 7109 12696
rect 7064 12656 7070 12668
rect 8481 12665 8493 12699
rect 8527 12696 8539 12699
rect 8935 12699 8993 12705
rect 8935 12696 8947 12699
rect 8527 12668 8947 12696
rect 8527 12665 8539 12668
rect 8481 12659 8539 12665
rect 8935 12665 8947 12668
rect 8981 12696 8993 12699
rect 9766 12696 9772 12708
rect 8981 12668 9772 12696
rect 8981 12665 8993 12668
rect 8935 12659 8993 12665
rect 9766 12656 9772 12668
rect 9824 12656 9830 12708
rect 11517 12699 11575 12705
rect 11517 12665 11529 12699
rect 11563 12696 11575 12699
rect 11606 12696 11612 12708
rect 11563 12668 11612 12696
rect 11563 12665 11575 12668
rect 11517 12659 11575 12665
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 12526 12696 12532 12708
rect 12487 12668 12532 12696
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 12621 12699 12679 12705
rect 12621 12665 12633 12699
rect 12667 12665 12679 12699
rect 13786 12696 13814 12804
rect 14550 12792 14556 12804
rect 14608 12832 14614 12844
rect 15841 12835 15899 12841
rect 15841 12832 15853 12835
rect 14608 12804 15853 12832
rect 14608 12792 14614 12804
rect 15841 12801 15853 12804
rect 15887 12832 15899 12835
rect 16298 12832 16304 12844
rect 15887 12804 16304 12832
rect 15887 12801 15899 12804
rect 15841 12795 15899 12801
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 20346 12832 20352 12844
rect 16567 12804 20352 12832
rect 14274 12696 14280 12708
rect 13786 12668 14280 12696
rect 12621 12659 12679 12665
rect 8018 12628 8024 12640
rect 6880 12600 6960 12628
rect 7979 12600 8024 12628
rect 6880 12588 6886 12600
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 9490 12628 9496 12640
rect 9451 12600 9496 12628
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 12253 12631 12311 12637
rect 12253 12597 12265 12631
rect 12299 12628 12311 12631
rect 12434 12628 12440 12640
rect 12299 12600 12440 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 12434 12588 12440 12600
rect 12492 12628 12498 12640
rect 12636 12628 12664 12659
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 14369 12699 14427 12705
rect 14369 12665 14381 12699
rect 14415 12696 14427 12699
rect 14734 12696 14740 12708
rect 14415 12668 14740 12696
rect 14415 12665 14427 12668
rect 14369 12659 14427 12665
rect 14734 12656 14740 12668
rect 14792 12656 14798 12708
rect 15930 12696 15936 12708
rect 15843 12668 15936 12696
rect 15930 12656 15936 12668
rect 15988 12656 15994 12708
rect 16206 12656 16212 12708
rect 16264 12696 16270 12708
rect 16567 12696 16595 12804
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 22002 12832 22008 12844
rect 21963 12804 22008 12832
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 22649 12835 22707 12841
rect 22649 12801 22661 12835
rect 22695 12832 22707 12835
rect 23198 12832 23204 12844
rect 22695 12804 23204 12832
rect 22695 12801 22707 12804
rect 22649 12795 22707 12801
rect 23198 12792 23204 12804
rect 23256 12832 23262 12844
rect 24029 12835 24087 12841
rect 24029 12832 24041 12835
rect 23256 12804 24041 12832
rect 23256 12792 23262 12804
rect 24029 12801 24041 12804
rect 24075 12801 24087 12835
rect 24688 12832 24716 12931
rect 25225 12835 25283 12841
rect 25225 12832 25237 12835
rect 24688 12804 25237 12832
rect 24029 12795 24087 12801
rect 25225 12801 25237 12804
rect 25271 12801 25283 12835
rect 25225 12795 25283 12801
rect 17770 12724 17776 12776
rect 17828 12764 17834 12776
rect 18233 12767 18291 12773
rect 18233 12764 18245 12767
rect 17828 12736 18245 12764
rect 17828 12724 17834 12736
rect 18233 12733 18245 12736
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 18693 12767 18751 12773
rect 18693 12733 18705 12767
rect 18739 12733 18751 12767
rect 18693 12727 18751 12733
rect 20165 12767 20223 12773
rect 20165 12733 20177 12767
rect 20211 12764 20223 12767
rect 20254 12764 20260 12776
rect 20211 12736 20260 12764
rect 20211 12733 20223 12736
rect 20165 12727 20223 12733
rect 18708 12696 18736 12727
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 21085 12767 21143 12773
rect 21085 12733 21097 12767
rect 21131 12764 21143 12767
rect 21729 12767 21787 12773
rect 21729 12764 21741 12767
rect 21131 12736 21741 12764
rect 21131 12733 21143 12736
rect 21085 12727 21143 12733
rect 21729 12733 21741 12736
rect 21775 12733 21787 12767
rect 21729 12727 21787 12733
rect 16264 12668 16595 12696
rect 17788 12668 18736 12696
rect 18969 12699 19027 12705
rect 16264 12656 16270 12668
rect 12492 12600 12664 12628
rect 12492 12588 12498 12600
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 15197 12631 15255 12637
rect 15197 12628 15209 12631
rect 14884 12600 15209 12628
rect 14884 12588 14890 12600
rect 15197 12597 15209 12600
rect 15243 12628 15255 12631
rect 15565 12631 15623 12637
rect 15565 12628 15577 12631
rect 15243 12600 15577 12628
rect 15243 12597 15255 12600
rect 15197 12591 15255 12597
rect 15565 12597 15577 12600
rect 15611 12628 15623 12631
rect 15948 12628 15976 12656
rect 17788 12640 17816 12668
rect 18969 12665 18981 12699
rect 19015 12696 19027 12699
rect 20346 12696 20352 12708
rect 19015 12668 20352 12696
rect 19015 12665 19027 12668
rect 18969 12659 19027 12665
rect 20346 12656 20352 12668
rect 20404 12656 20410 12708
rect 20486 12699 20544 12705
rect 20486 12665 20498 12699
rect 20532 12665 20544 12699
rect 20486 12659 20544 12665
rect 15611 12600 15976 12628
rect 17129 12631 17187 12637
rect 15611 12597 15623 12600
rect 15565 12591 15623 12597
rect 17129 12597 17141 12631
rect 17175 12628 17187 12631
rect 17218 12628 17224 12640
rect 17175 12600 17224 12628
rect 17175 12597 17187 12600
rect 17129 12591 17187 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17497 12631 17555 12637
rect 17497 12597 17509 12631
rect 17543 12628 17555 12631
rect 17770 12628 17776 12640
rect 17543 12600 17776 12628
rect 17543 12597 17555 12600
rect 17497 12591 17555 12597
rect 17770 12588 17776 12600
rect 17828 12588 17834 12640
rect 20070 12588 20076 12640
rect 20128 12628 20134 12640
rect 20501 12628 20529 12659
rect 21542 12628 21548 12640
rect 20128 12600 21548 12628
rect 20128 12588 20134 12600
rect 21542 12588 21548 12600
rect 21600 12588 21606 12640
rect 21744 12628 21772 12727
rect 22097 12699 22155 12705
rect 22097 12665 22109 12699
rect 22143 12665 22155 12699
rect 23750 12696 23756 12708
rect 23711 12668 23756 12696
rect 22097 12659 22155 12665
rect 22112 12628 22140 12659
rect 23750 12656 23756 12668
rect 23808 12656 23814 12708
rect 23842 12656 23848 12708
rect 23900 12696 23906 12708
rect 23900 12668 23945 12696
rect 23900 12656 23906 12668
rect 22922 12628 22928 12640
rect 21744 12600 22140 12628
rect 22883 12600 22928 12628
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1673 12427 1731 12433
rect 1673 12393 1685 12427
rect 1719 12424 1731 12427
rect 1946 12424 1952 12436
rect 1719 12396 1952 12424
rect 1719 12393 1731 12396
rect 1673 12387 1731 12393
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 2130 12424 2136 12436
rect 2087 12396 2136 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2130 12384 2136 12396
rect 2188 12424 2194 12436
rect 3142 12424 3148 12436
rect 2188 12396 3148 12424
rect 2188 12384 2194 12396
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 3786 12424 3792 12436
rect 3747 12396 3792 12424
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 5074 12424 5080 12436
rect 5035 12396 5080 12424
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 6917 12427 6975 12433
rect 6917 12393 6929 12427
rect 6963 12424 6975 12427
rect 7006 12424 7012 12436
rect 6963 12396 7012 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7006 12384 7012 12396
rect 7064 12424 7070 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 7064 12396 7205 12424
rect 7064 12384 7070 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 7926 12424 7932 12436
rect 7887 12396 7932 12424
rect 7193 12387 7251 12393
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 11422 12424 11428 12436
rect 11383 12396 11428 12424
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 11977 12427 12035 12433
rect 11977 12424 11989 12427
rect 11940 12396 11989 12424
rect 11940 12384 11946 12396
rect 11977 12393 11989 12396
rect 12023 12393 12035 12427
rect 11977 12387 12035 12393
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12529 12427 12587 12433
rect 12529 12424 12541 12427
rect 12492 12396 12541 12424
rect 12492 12384 12498 12396
rect 12529 12393 12541 12396
rect 12575 12393 12587 12427
rect 12529 12387 12587 12393
rect 14274 12384 14280 12436
rect 14332 12424 14338 12436
rect 15013 12427 15071 12433
rect 15013 12424 15025 12427
rect 14332 12396 15025 12424
rect 14332 12384 14338 12396
rect 15013 12393 15025 12396
rect 15059 12393 15071 12427
rect 16298 12424 16304 12436
rect 16259 12396 16304 12424
rect 15013 12387 15071 12393
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19613 12427 19671 12433
rect 19613 12424 19625 12427
rect 19484 12396 19625 12424
rect 19484 12384 19490 12396
rect 19613 12393 19625 12396
rect 19659 12393 19671 12427
rect 19613 12387 19671 12393
rect 20717 12427 20775 12433
rect 20717 12393 20729 12427
rect 20763 12424 20775 12427
rect 20990 12424 20996 12436
rect 20763 12396 20996 12424
rect 20763 12393 20775 12396
rect 20717 12387 20775 12393
rect 20990 12384 20996 12396
rect 21048 12384 21054 12436
rect 21542 12424 21548 12436
rect 21503 12396 21548 12424
rect 21542 12384 21548 12396
rect 21600 12384 21606 12436
rect 22097 12427 22155 12433
rect 22097 12393 22109 12427
rect 22143 12424 22155 12427
rect 22922 12424 22928 12436
rect 22143 12396 22928 12424
rect 22143 12393 22155 12396
rect 22097 12387 22155 12393
rect 22922 12384 22928 12396
rect 22980 12384 22986 12436
rect 23753 12427 23811 12433
rect 23753 12393 23765 12427
rect 23799 12424 23811 12427
rect 23842 12424 23848 12436
rect 23799 12396 23848 12424
rect 23799 12393 23811 12396
rect 23753 12387 23811 12393
rect 23842 12384 23848 12396
rect 23900 12384 23906 12436
rect 2222 12316 2228 12368
rect 2280 12356 2286 12368
rect 2317 12359 2375 12365
rect 2317 12356 2329 12359
rect 2280 12328 2329 12356
rect 2280 12316 2286 12328
rect 2317 12325 2329 12328
rect 2363 12325 2375 12359
rect 2317 12319 2375 12325
rect 2590 12316 2596 12368
rect 2648 12356 2654 12368
rect 4154 12356 4160 12368
rect 2648 12328 4160 12356
rect 2648 12316 2654 12328
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 4338 12316 4344 12368
rect 4396 12356 4402 12368
rect 4478 12359 4536 12365
rect 4478 12356 4490 12359
rect 4396 12328 4490 12356
rect 4396 12316 4402 12328
rect 4478 12325 4490 12328
rect 4524 12325 4536 12359
rect 4478 12319 4536 12325
rect 5994 12316 6000 12368
rect 6052 12356 6058 12368
rect 6318 12359 6376 12365
rect 6318 12356 6330 12359
rect 6052 12328 6330 12356
rect 6052 12316 6058 12328
rect 6318 12325 6330 12328
rect 6364 12325 6376 12359
rect 6318 12319 6376 12325
rect 8205 12359 8263 12365
rect 8205 12325 8217 12359
rect 8251 12356 8263 12359
rect 9490 12356 9496 12368
rect 8251 12328 9496 12356
rect 8251 12325 8263 12328
rect 8205 12319 8263 12325
rect 9490 12316 9496 12328
rect 9548 12316 9554 12368
rect 13817 12359 13875 12365
rect 13817 12325 13829 12359
rect 13863 12356 13875 12359
rect 13906 12356 13912 12368
rect 13863 12328 13912 12356
rect 13863 12325 13875 12328
rect 13817 12319 13875 12325
rect 13906 12316 13912 12328
rect 13964 12316 13970 12368
rect 14369 12359 14427 12365
rect 14369 12325 14381 12359
rect 14415 12356 14427 12359
rect 14550 12356 14556 12368
rect 14415 12328 14556 12356
rect 14415 12325 14427 12328
rect 14369 12319 14427 12325
rect 14550 12316 14556 12328
rect 14608 12316 14614 12368
rect 15473 12359 15531 12365
rect 15473 12325 15485 12359
rect 15519 12356 15531 12359
rect 15562 12356 15568 12368
rect 15519 12328 15568 12356
rect 15519 12325 15531 12328
rect 15473 12319 15531 12325
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 16022 12356 16028 12368
rect 15983 12328 16028 12356
rect 16022 12316 16028 12328
rect 16080 12316 16086 12368
rect 18782 12316 18788 12368
rect 18840 12356 18846 12368
rect 19014 12359 19072 12365
rect 19014 12356 19026 12359
rect 18840 12328 19026 12356
rect 18840 12316 18846 12328
rect 19014 12325 19026 12328
rect 19060 12325 19072 12359
rect 19014 12319 19072 12325
rect 21082 12316 21088 12368
rect 21140 12356 21146 12368
rect 24305 12359 24363 12365
rect 24305 12356 24317 12359
rect 21140 12328 21404 12356
rect 21140 12316 21146 12328
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 16942 12288 16948 12300
rect 16903 12260 16948 12288
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 18414 12248 18420 12300
rect 18472 12288 18478 12300
rect 18693 12291 18751 12297
rect 18693 12288 18705 12291
rect 18472 12260 18705 12288
rect 18472 12248 18478 12260
rect 18693 12257 18705 12260
rect 18739 12257 18751 12291
rect 18693 12251 18751 12257
rect 20346 12248 20352 12300
rect 20404 12288 20410 12300
rect 21177 12291 21235 12297
rect 21177 12288 21189 12291
rect 20404 12260 21189 12288
rect 20404 12248 20410 12260
rect 21177 12257 21189 12260
rect 21223 12257 21235 12291
rect 21376 12288 21404 12328
rect 23446 12328 24317 12356
rect 23198 12288 23204 12300
rect 21376 12260 23204 12288
rect 21177 12251 21235 12257
rect 23198 12248 23204 12260
rect 23256 12288 23262 12300
rect 23446 12288 23474 12328
rect 24305 12325 24317 12328
rect 24351 12325 24363 12359
rect 24305 12319 24363 12325
rect 24857 12359 24915 12365
rect 24857 12325 24869 12359
rect 24903 12356 24915 12359
rect 25038 12356 25044 12368
rect 24903 12328 25044 12356
rect 24903 12325 24915 12328
rect 24857 12319 24915 12325
rect 25038 12316 25044 12328
rect 25096 12316 25102 12368
rect 23256 12260 23474 12288
rect 23256 12248 23262 12260
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12189 2283 12223
rect 2590 12220 2596 12232
rect 2551 12192 2596 12220
rect 2225 12183 2283 12189
rect 2240 12152 2268 12183
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 5442 12220 5448 12232
rect 4203 12192 5448 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 5997 12223 6055 12229
rect 5997 12189 6009 12223
rect 6043 12220 6055 12223
rect 6546 12220 6552 12232
rect 6043 12192 6552 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 8386 12220 8392 12232
rect 8159 12192 8392 12220
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 11606 12220 11612 12232
rect 11567 12192 11612 12220
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 13814 12220 13820 12232
rect 13771 12192 13820 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12220 15439 12223
rect 15746 12220 15752 12232
rect 15427 12192 15752 12220
rect 15427 12189 15439 12192
rect 15381 12183 15439 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 16850 12220 16856 12232
rect 16811 12192 16856 12220
rect 16850 12180 16856 12192
rect 16908 12180 16914 12232
rect 17034 12180 17040 12232
rect 17092 12220 17098 12232
rect 22925 12223 22983 12229
rect 22925 12220 22937 12223
rect 17092 12192 22937 12220
rect 17092 12180 17098 12192
rect 22925 12189 22937 12192
rect 22971 12189 22983 12223
rect 24210 12220 24216 12232
rect 24171 12192 24216 12220
rect 22925 12183 22983 12189
rect 24210 12180 24216 12192
rect 24268 12180 24274 12232
rect 3050 12152 3056 12164
rect 2240 12124 3056 12152
rect 3050 12112 3056 12124
rect 3108 12112 3114 12164
rect 3326 12112 3332 12164
rect 3384 12152 3390 12164
rect 4522 12152 4528 12164
rect 3384 12124 4528 12152
rect 3384 12112 3390 12124
rect 4522 12112 4528 12124
rect 4580 12152 4586 12164
rect 8665 12155 8723 12161
rect 8665 12152 8677 12155
rect 4580 12124 8677 12152
rect 4580 12112 4586 12124
rect 8665 12121 8677 12124
rect 8711 12121 8723 12155
rect 8665 12115 8723 12121
rect 17770 12112 17776 12164
rect 17828 12152 17834 12164
rect 18325 12155 18383 12161
rect 18325 12152 18337 12155
rect 17828 12124 18337 12152
rect 17828 12112 17834 12124
rect 18325 12121 18337 12124
rect 18371 12152 18383 12155
rect 18966 12152 18972 12164
rect 18371 12124 18972 12152
rect 18371 12121 18383 12124
rect 18325 12115 18383 12121
rect 18966 12112 18972 12124
rect 19024 12152 19030 12164
rect 20990 12152 20996 12164
rect 19024 12124 20996 12152
rect 19024 12112 19030 12124
rect 20990 12112 20996 12124
rect 21048 12112 21054 12164
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 2774 12084 2780 12096
rect 2096 12056 2780 12084
rect 2096 12044 2102 12056
rect 2774 12044 2780 12056
rect 2832 12044 2838 12096
rect 8754 12044 8760 12096
rect 8812 12084 8818 12096
rect 9033 12087 9091 12093
rect 9033 12084 9045 12087
rect 8812 12056 9045 12084
rect 8812 12044 8818 12056
rect 9033 12053 9045 12056
rect 9079 12053 9091 12087
rect 10502 12084 10508 12096
rect 10463 12056 10508 12084
rect 9033 12047 9091 12053
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 11054 12084 11060 12096
rect 11015 12056 11060 12084
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12894 12084 12900 12096
rect 12584 12056 12900 12084
rect 12584 12044 12590 12056
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 13541 12087 13599 12093
rect 13541 12053 13553 12087
rect 13587 12084 13599 12087
rect 13630 12084 13636 12096
rect 13587 12056 13636 12084
rect 13587 12053 13599 12056
rect 13541 12047 13599 12053
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 14734 12084 14740 12096
rect 14695 12056 14740 12084
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 19150 12084 19156 12096
rect 15436 12056 19156 12084
rect 15436 12044 15442 12056
rect 19150 12044 19156 12056
rect 19208 12044 19214 12096
rect 20254 12084 20260 12096
rect 20215 12056 20260 12084
rect 20254 12044 20260 12056
rect 20312 12044 20318 12096
rect 22646 12084 22652 12096
rect 22607 12056 22652 12084
rect 22646 12044 22652 12056
rect 22704 12044 22710 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2222 11840 2228 11892
rect 2280 11880 2286 11892
rect 3329 11883 3387 11889
rect 3329 11880 3341 11883
rect 2280 11852 3341 11880
rect 2280 11840 2286 11852
rect 3329 11849 3341 11852
rect 3375 11849 3387 11883
rect 3329 11843 3387 11849
rect 2590 11812 2596 11824
rect 2551 11784 2596 11812
rect 2590 11772 2596 11784
rect 2648 11772 2654 11824
rect 3344 11812 3372 11843
rect 3878 11840 3884 11892
rect 3936 11880 3942 11892
rect 5169 11883 5227 11889
rect 5169 11880 5181 11883
rect 3936 11852 5181 11880
rect 3936 11840 3942 11852
rect 5169 11849 5181 11852
rect 5215 11849 5227 11883
rect 5442 11880 5448 11892
rect 5403 11852 5448 11880
rect 5169 11843 5227 11849
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 7239 11883 7297 11889
rect 7239 11849 7251 11883
rect 7285 11880 7297 11883
rect 9214 11880 9220 11892
rect 7285 11852 9220 11880
rect 7285 11849 7297 11852
rect 7239 11843 7297 11849
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9398 11880 9404 11892
rect 9359 11852 9404 11880
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 9677 11883 9735 11889
rect 9677 11880 9689 11883
rect 9548 11852 9689 11880
rect 9548 11840 9554 11852
rect 9677 11849 9689 11852
rect 9723 11849 9735 11883
rect 9677 11843 9735 11849
rect 10502 11840 10508 11892
rect 10560 11880 10566 11892
rect 10597 11883 10655 11889
rect 10597 11880 10609 11883
rect 10560 11852 10609 11880
rect 10560 11840 10566 11852
rect 10597 11849 10609 11852
rect 10643 11880 10655 11883
rect 10962 11880 10968 11892
rect 10643 11852 10968 11880
rect 10643 11849 10655 11852
rect 10597 11843 10655 11849
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12805 11883 12863 11889
rect 12805 11849 12817 11883
rect 12851 11880 12863 11883
rect 13262 11880 13268 11892
rect 12851 11852 13268 11880
rect 12851 11849 12863 11852
rect 12805 11843 12863 11849
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 14553 11883 14611 11889
rect 14553 11849 14565 11883
rect 14599 11880 14611 11883
rect 14826 11880 14832 11892
rect 14599 11852 14832 11880
rect 14599 11849 14611 11852
rect 14553 11843 14611 11849
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 14921 11883 14979 11889
rect 14921 11849 14933 11883
rect 14967 11880 14979 11883
rect 15562 11880 15568 11892
rect 14967 11852 15568 11880
rect 14967 11849 14979 11852
rect 14921 11843 14979 11849
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 17865 11883 17923 11889
rect 17865 11849 17877 11883
rect 17911 11880 17923 11883
rect 18414 11880 18420 11892
rect 17911 11852 18420 11880
rect 17911 11849 17923 11852
rect 17865 11843 17923 11849
rect 18414 11840 18420 11852
rect 18472 11840 18478 11892
rect 19797 11883 19855 11889
rect 19797 11849 19809 11883
rect 19843 11880 19855 11883
rect 21082 11880 21088 11892
rect 19843 11852 21088 11880
rect 19843 11849 19855 11852
rect 19797 11843 19855 11849
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 21269 11883 21327 11889
rect 21269 11849 21281 11883
rect 21315 11880 21327 11883
rect 21542 11880 21548 11892
rect 21315 11852 21548 11880
rect 21315 11849 21327 11852
rect 21269 11843 21327 11849
rect 21542 11840 21548 11852
rect 21600 11880 21606 11892
rect 21637 11883 21695 11889
rect 21637 11880 21649 11883
rect 21600 11852 21649 11880
rect 21600 11840 21606 11852
rect 21637 11849 21649 11852
rect 21683 11849 21695 11883
rect 21637 11843 21695 11849
rect 22741 11883 22799 11889
rect 22741 11849 22753 11883
rect 22787 11880 22799 11883
rect 23842 11880 23848 11892
rect 22787 11852 23848 11880
rect 22787 11849 22799 11852
rect 22741 11843 22799 11849
rect 23842 11840 23848 11852
rect 23900 11840 23906 11892
rect 24210 11840 24216 11892
rect 24268 11880 24274 11892
rect 24854 11880 24860 11892
rect 24268 11852 24860 11880
rect 24268 11840 24274 11852
rect 24854 11840 24860 11852
rect 24912 11880 24918 11892
rect 25041 11883 25099 11889
rect 25041 11880 25053 11883
rect 24912 11852 25053 11880
rect 24912 11840 24918 11852
rect 25041 11849 25053 11852
rect 25087 11849 25099 11883
rect 25041 11843 25099 11849
rect 8018 11812 8024 11824
rect 3344 11784 8024 11812
rect 8018 11772 8024 11784
rect 8076 11812 8082 11824
rect 9033 11815 9091 11821
rect 9033 11812 9045 11815
rect 8076 11784 9045 11812
rect 8076 11772 8082 11784
rect 9033 11781 9045 11784
rect 9079 11781 9091 11815
rect 9033 11775 9091 11781
rect 6638 11744 6644 11756
rect 2700 11716 6644 11744
rect 1854 11568 1860 11620
rect 1912 11608 1918 11620
rect 2041 11611 2099 11617
rect 2041 11608 2053 11611
rect 1912 11580 2053 11608
rect 1912 11568 1918 11580
rect 2041 11577 2053 11580
rect 2087 11577 2099 11611
rect 2041 11571 2099 11577
rect 2133 11611 2191 11617
rect 2133 11577 2145 11611
rect 2179 11608 2191 11611
rect 2700 11608 2728 11716
rect 6638 11704 6644 11716
rect 6696 11744 6702 11756
rect 7006 11744 7012 11756
rect 6696 11716 7012 11744
rect 6696 11704 6702 11716
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11744 8171 11747
rect 9416 11744 9444 11840
rect 15378 11812 15384 11824
rect 12636 11784 15384 11812
rect 11146 11744 11152 11756
rect 8159 11716 9444 11744
rect 11107 11716 11152 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 3789 11679 3847 11685
rect 3789 11645 3801 11679
rect 3835 11676 3847 11679
rect 4246 11676 4252 11688
rect 3835 11648 4252 11676
rect 3835 11645 3847 11648
rect 3789 11639 3847 11645
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 4798 11636 4804 11688
rect 4856 11676 4862 11688
rect 7136 11679 7194 11685
rect 7136 11676 7148 11679
rect 4856 11648 7148 11676
rect 4856 11636 4862 11648
rect 7136 11645 7148 11648
rect 7182 11676 7194 11679
rect 7558 11676 7564 11688
rect 7182 11648 7564 11676
rect 7182 11645 7194 11648
rect 7136 11639 7194 11645
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 12636 11685 12664 11784
rect 15378 11772 15384 11784
rect 15436 11772 15442 11824
rect 16853 11815 16911 11821
rect 15488 11784 16528 11812
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11744 13231 11747
rect 13906 11744 13912 11756
rect 13219 11716 13912 11744
rect 13219 11713 13231 11716
rect 13173 11707 13231 11713
rect 13906 11704 13912 11716
rect 13964 11744 13970 11756
rect 15488 11753 15516 11784
rect 15473 11747 15531 11753
rect 13964 11716 15332 11744
rect 13964 11704 13970 11716
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11676 12311 11679
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12299 11648 12633 11676
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 13630 11676 13636 11688
rect 13591 11648 13636 11676
rect 12621 11639 12679 11645
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 2179 11580 2728 11608
rect 4157 11611 4215 11617
rect 2179 11577 2191 11580
rect 2133 11571 2191 11577
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4338 11608 4344 11620
rect 4203 11580 4344 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 1765 11543 1823 11549
rect 1765 11509 1777 11543
rect 1811 11540 1823 11543
rect 1946 11540 1952 11552
rect 1811 11512 1952 11540
rect 1811 11509 1823 11512
rect 1765 11503 1823 11509
rect 1946 11500 1952 11512
rect 2004 11540 2010 11552
rect 2148 11540 2176 11571
rect 4338 11568 4344 11580
rect 4396 11608 4402 11620
rect 4611 11611 4669 11617
rect 4611 11608 4623 11611
rect 4396 11580 4623 11608
rect 4396 11568 4402 11580
rect 4611 11577 4623 11580
rect 4657 11608 4669 11611
rect 5994 11608 6000 11620
rect 4657 11580 6000 11608
rect 4657 11577 4669 11580
rect 4611 11571 4669 11577
rect 5994 11568 6000 11580
rect 6052 11608 6058 11620
rect 6089 11611 6147 11617
rect 6089 11608 6101 11611
rect 6052 11580 6101 11608
rect 6052 11568 6058 11580
rect 6089 11577 6101 11580
rect 6135 11608 6147 11611
rect 8021 11611 8079 11617
rect 8021 11608 8033 11611
rect 6135 11580 8033 11608
rect 6135 11577 6147 11580
rect 6089 11571 6147 11577
rect 6196 11552 6224 11580
rect 8021 11577 8033 11580
rect 8067 11608 8079 11611
rect 8475 11611 8533 11617
rect 8475 11608 8487 11611
rect 8067 11580 8487 11608
rect 8067 11577 8079 11580
rect 8021 11571 8079 11577
rect 8475 11577 8487 11580
rect 8521 11608 8533 11611
rect 8662 11608 8668 11620
rect 8521 11580 8668 11608
rect 8521 11577 8533 11580
rect 8475 11571 8533 11577
rect 8662 11568 8668 11580
rect 8720 11568 8726 11620
rect 10873 11611 10931 11617
rect 10873 11577 10885 11611
rect 10919 11577 10931 11611
rect 10873 11571 10931 11577
rect 3050 11540 3056 11552
rect 2004 11512 2176 11540
rect 3011 11512 3056 11540
rect 2004 11500 2010 11512
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 6178 11500 6184 11552
rect 6236 11500 6242 11552
rect 6457 11543 6515 11549
rect 6457 11509 6469 11543
rect 6503 11540 6515 11543
rect 6546 11540 6552 11552
rect 6503 11512 6552 11540
rect 6503 11509 6515 11512
rect 6457 11503 6515 11509
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 10100 11512 10241 11540
rect 10100 11500 10106 11512
rect 10229 11509 10241 11512
rect 10275 11540 10287 11543
rect 10888 11540 10916 11571
rect 10962 11568 10968 11620
rect 11020 11608 11026 11620
rect 11020 11580 11065 11608
rect 11020 11568 11026 11580
rect 11238 11568 11244 11620
rect 11296 11608 11302 11620
rect 11882 11608 11888 11620
rect 11296 11580 11888 11608
rect 11296 11568 11302 11580
rect 11882 11568 11888 11580
rect 11940 11608 11946 11620
rect 13449 11611 13507 11617
rect 13449 11608 13461 11611
rect 11940 11580 13461 11608
rect 11940 11568 11946 11580
rect 13449 11577 13461 11580
rect 13495 11608 13507 11611
rect 13722 11608 13728 11620
rect 13495 11580 13728 11608
rect 13495 11577 13507 11580
rect 13449 11571 13507 11577
rect 13722 11568 13728 11580
rect 13780 11608 13786 11620
rect 13954 11611 14012 11617
rect 13954 11608 13966 11611
rect 13780 11580 13966 11608
rect 13780 11568 13786 11580
rect 13954 11577 13966 11580
rect 14000 11577 14012 11611
rect 13954 11571 14012 11577
rect 15304 11549 15332 11716
rect 15473 11713 15485 11747
rect 15519 11713 15531 11747
rect 15746 11744 15752 11756
rect 15707 11716 15752 11744
rect 15473 11707 15531 11713
rect 15746 11704 15752 11716
rect 15804 11704 15810 11756
rect 16500 11753 16528 11784
rect 16853 11781 16865 11815
rect 16899 11812 16911 11815
rect 16942 11812 16948 11824
rect 16899 11784 16948 11812
rect 16899 11781 16911 11784
rect 16853 11775 16911 11781
rect 16942 11772 16948 11784
rect 17000 11772 17006 11824
rect 17126 11812 17132 11824
rect 17087 11784 17132 11812
rect 17126 11772 17132 11784
rect 17184 11772 17190 11824
rect 19978 11772 19984 11824
rect 20036 11812 20042 11824
rect 20036 11784 22185 11812
rect 20036 11772 20042 11784
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 17034 11744 17040 11756
rect 16531 11716 17040 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 18417 11747 18475 11753
rect 18417 11713 18429 11747
rect 18463 11744 18475 11747
rect 18874 11744 18880 11756
rect 18463 11716 18880 11744
rect 18463 11713 18475 11716
rect 18417 11707 18475 11713
rect 18874 11704 18880 11716
rect 18932 11704 18938 11756
rect 20070 11744 20076 11756
rect 19213 11716 20076 11744
rect 16945 11679 17003 11685
rect 16945 11645 16957 11679
rect 16991 11676 17003 11679
rect 17218 11676 17224 11688
rect 16991 11648 17224 11676
rect 16991 11645 17003 11648
rect 16945 11639 17003 11645
rect 17218 11636 17224 11648
rect 17276 11676 17282 11688
rect 17276 11648 17540 11676
rect 17276 11636 17282 11648
rect 15565 11611 15623 11617
rect 15565 11577 15577 11611
rect 15611 11608 15623 11611
rect 16850 11608 16856 11620
rect 15611 11580 16856 11608
rect 15611 11577 15623 11580
rect 15565 11571 15623 11577
rect 10275 11512 10916 11540
rect 15289 11543 15347 11549
rect 10275 11509 10287 11512
rect 10229 11503 10287 11509
rect 15289 11509 15301 11543
rect 15335 11540 15347 11543
rect 15580 11540 15608 11571
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 17512 11552 17540 11648
rect 19213 11617 19241 11716
rect 20070 11704 20076 11716
rect 20128 11704 20134 11756
rect 20625 11679 20683 11685
rect 20625 11676 20637 11679
rect 20456 11648 20637 11676
rect 19198 11611 19256 11617
rect 19198 11608 19210 11611
rect 18800 11580 19210 11608
rect 18800 11552 18828 11580
rect 19198 11577 19210 11580
rect 19244 11577 19256 11611
rect 19198 11571 19256 11577
rect 20456 11552 20484 11648
rect 20625 11645 20637 11648
rect 20671 11645 20683 11679
rect 21818 11676 21824 11688
rect 21779 11648 21824 11676
rect 20625 11639 20683 11645
rect 21818 11636 21824 11648
rect 21876 11636 21882 11688
rect 22157 11676 22185 11784
rect 23934 11772 23940 11824
rect 23992 11812 23998 11824
rect 23992 11784 25176 11812
rect 23992 11772 23998 11784
rect 23477 11747 23535 11753
rect 23477 11713 23489 11747
rect 23523 11744 23535 11747
rect 24121 11747 24179 11753
rect 24121 11744 24133 11747
rect 23523 11716 24133 11744
rect 23523 11713 23535 11716
rect 23477 11707 23535 11713
rect 24121 11713 24133 11716
rect 24167 11744 24179 11747
rect 24210 11744 24216 11756
rect 24167 11716 24216 11744
rect 24167 11713 24179 11716
rect 24121 11707 24179 11713
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 24765 11747 24823 11753
rect 24765 11713 24777 11747
rect 24811 11744 24823 11747
rect 25038 11744 25044 11756
rect 24811 11716 25044 11744
rect 24811 11713 24823 11716
rect 24765 11707 24823 11713
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 23566 11676 23572 11688
rect 22157 11648 23572 11676
rect 23566 11636 23572 11648
rect 23624 11676 23630 11688
rect 23845 11679 23903 11685
rect 23845 11676 23857 11679
rect 23624 11648 23857 11676
rect 23624 11636 23630 11648
rect 23845 11645 23857 11648
rect 23891 11645 23903 11679
rect 25148 11676 25176 11784
rect 25628 11679 25686 11685
rect 25628 11676 25640 11679
rect 25148 11648 25640 11676
rect 23845 11639 23903 11645
rect 25628 11645 25640 11648
rect 25674 11676 25686 11679
rect 26053 11679 26111 11685
rect 26053 11676 26065 11679
rect 25674 11648 26065 11676
rect 25674 11645 25686 11648
rect 25628 11639 25686 11645
rect 26053 11645 26065 11648
rect 26099 11645 26111 11679
rect 26053 11639 26111 11645
rect 21542 11568 21548 11620
rect 21600 11608 21606 11620
rect 22142 11611 22200 11617
rect 22142 11608 22154 11611
rect 21600 11580 22154 11608
rect 21600 11568 21606 11580
rect 22142 11577 22154 11580
rect 22188 11577 22200 11611
rect 23860 11608 23888 11639
rect 24213 11611 24271 11617
rect 24213 11608 24225 11611
rect 23860 11580 24225 11608
rect 22142 11571 22200 11577
rect 24213 11577 24225 11580
rect 24259 11577 24271 11611
rect 24213 11571 24271 11577
rect 17494 11540 17500 11552
rect 15335 11512 15608 11540
rect 17455 11512 17500 11540
rect 15335 11509 15347 11512
rect 15289 11503 15347 11509
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 18782 11540 18788 11552
rect 18743 11512 18788 11540
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 20438 11540 20444 11552
rect 20399 11512 20444 11540
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 20809 11543 20867 11549
rect 20809 11509 20821 11543
rect 20855 11540 20867 11543
rect 20990 11540 20996 11552
rect 20855 11512 20996 11540
rect 20855 11509 20867 11512
rect 20809 11503 20867 11509
rect 20990 11500 20996 11512
rect 21048 11500 21054 11552
rect 25130 11500 25136 11552
rect 25188 11540 25194 11552
rect 25731 11543 25789 11549
rect 25731 11540 25743 11543
rect 25188 11512 25743 11540
rect 25188 11500 25194 11512
rect 25731 11509 25743 11512
rect 25777 11509 25789 11543
rect 25731 11503 25789 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 4246 11296 4252 11348
rect 4304 11336 4310 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4304 11308 4537 11336
rect 4304 11296 4310 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 7006 11336 7012 11348
rect 6967 11308 7012 11336
rect 4525 11299 4583 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7929 11339 7987 11345
rect 7929 11305 7941 11339
rect 7975 11336 7987 11339
rect 8386 11336 8392 11348
rect 7975 11308 8392 11336
rect 7975 11305 7987 11308
rect 7929 11299 7987 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11336 10198 11348
rect 11606 11336 11612 11348
rect 10192 11308 10548 11336
rect 11567 11308 11612 11336
rect 10192 11296 10198 11308
rect 1762 11228 1768 11280
rect 1820 11268 1826 11280
rect 2222 11268 2228 11280
rect 1820 11240 2228 11268
rect 1820 11228 1826 11240
rect 2222 11228 2228 11240
rect 2280 11228 2286 11280
rect 2777 11271 2835 11277
rect 2777 11237 2789 11271
rect 2823 11268 2835 11271
rect 2958 11268 2964 11280
rect 2823 11240 2964 11268
rect 2823 11237 2835 11240
rect 2777 11231 2835 11237
rect 2958 11228 2964 11240
rect 3016 11228 3022 11280
rect 4338 11268 4344 11280
rect 4299 11240 4344 11268
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 6178 11228 6184 11280
rect 6236 11268 6242 11280
rect 6410 11271 6468 11277
rect 6410 11268 6422 11271
rect 6236 11240 6422 11268
rect 6236 11228 6242 11240
rect 6410 11237 6422 11240
rect 6456 11237 6468 11271
rect 8754 11268 8760 11280
rect 8715 11240 8760 11268
rect 6410 11231 6468 11237
rect 8754 11228 8760 11240
rect 8812 11228 8818 11280
rect 10520 11277 10548 11308
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 12483 11339 12541 11345
rect 12483 11305 12495 11339
rect 12529 11336 12541 11339
rect 13814 11336 13820 11348
rect 12529 11308 13820 11336
rect 12529 11305 12541 11308
rect 12483 11299 12541 11305
rect 13814 11296 13820 11308
rect 13872 11336 13878 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 13872 11308 14933 11336
rect 13872 11296 13878 11308
rect 14921 11305 14933 11308
rect 14967 11305 14979 11339
rect 19978 11336 19984 11348
rect 19939 11308 19984 11336
rect 14921 11299 14979 11305
rect 19978 11296 19984 11308
rect 20036 11296 20042 11348
rect 20254 11296 20260 11348
rect 20312 11336 20318 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20312 11308 21005 11336
rect 20312 11296 20318 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 20993 11299 21051 11305
rect 24394 11296 24400 11348
rect 24452 11336 24458 11348
rect 24719 11339 24777 11345
rect 24719 11336 24731 11339
rect 24452 11308 24731 11336
rect 24452 11296 24458 11308
rect 24719 11305 24731 11308
rect 24765 11305 24777 11339
rect 24719 11299 24777 11305
rect 10505 11271 10563 11277
rect 10505 11237 10517 11271
rect 10551 11237 10563 11271
rect 10505 11231 10563 11237
rect 11057 11271 11115 11277
rect 11057 11237 11069 11271
rect 11103 11268 11115 11271
rect 11146 11268 11152 11280
rect 11103 11240 11152 11268
rect 11103 11237 11115 11240
rect 11057 11231 11115 11237
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 13722 11277 13728 11280
rect 13719 11268 13728 11277
rect 13683 11240 13728 11268
rect 13719 11231 13728 11240
rect 13722 11228 13728 11231
rect 13780 11228 13786 11280
rect 14734 11268 14740 11280
rect 14292 11240 14740 11268
rect 4246 11160 4252 11212
rect 4304 11200 4310 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4304 11172 4445 11200
rect 4304 11160 4310 11172
rect 4433 11169 4445 11172
rect 4479 11200 4491 11203
rect 4614 11200 4620 11212
rect 4479 11172 4620 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 4982 11200 4988 11212
rect 4943 11172 4988 11200
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 8294 11200 8300 11212
rect 8255 11172 8300 11200
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 8570 11200 8576 11212
rect 8531 11172 8576 11200
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 12380 11203 12438 11209
rect 12380 11200 12392 11203
rect 11618 11172 12392 11200
rect 2130 11132 2136 11144
rect 2091 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 6086 11132 6092 11144
rect 6047 11104 6092 11132
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 9416 11104 10425 11132
rect 1854 10996 1860 11008
rect 1815 10968 1860 10996
rect 1854 10956 1860 10968
rect 1912 10956 1918 11008
rect 8754 10956 8760 11008
rect 8812 10996 8818 11008
rect 9416 11005 9444 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 11330 11092 11336 11144
rect 11388 11132 11394 11144
rect 11618 11132 11646 11172
rect 12380 11169 12392 11172
rect 12426 11200 12438 11203
rect 12618 11200 12624 11212
rect 12426 11172 12624 11200
rect 12426 11169 12438 11172
rect 12380 11163 12438 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 14292 11209 14320 11240
rect 14734 11228 14740 11240
rect 14792 11268 14798 11280
rect 15473 11271 15531 11277
rect 15473 11268 15485 11271
rect 14792 11240 15485 11268
rect 14792 11228 14798 11240
rect 15473 11237 15485 11240
rect 15519 11268 15531 11271
rect 16942 11268 16948 11280
rect 15519 11240 16948 11268
rect 15519 11237 15531 11240
rect 15473 11231 15531 11237
rect 16942 11228 16948 11240
rect 17000 11228 17006 11280
rect 18782 11228 18788 11280
rect 18840 11268 18846 11280
rect 19382 11271 19440 11277
rect 19382 11268 19394 11271
rect 18840 11240 19394 11268
rect 18840 11228 18846 11240
rect 19382 11237 19394 11240
rect 19428 11237 19440 11271
rect 21818 11268 21824 11280
rect 19382 11231 19440 11237
rect 20501 11240 21824 11268
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11169 14335 11203
rect 17770 11200 17776 11212
rect 17731 11172 17776 11200
rect 14277 11163 14335 11169
rect 17770 11160 17776 11172
rect 17828 11160 17834 11212
rect 17954 11200 17960 11212
rect 17915 11172 17960 11200
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 18233 11203 18291 11209
rect 18233 11169 18245 11203
rect 18279 11200 18291 11203
rect 20501 11200 20529 11240
rect 21818 11228 21824 11240
rect 21876 11268 21882 11280
rect 21913 11271 21971 11277
rect 21913 11268 21925 11271
rect 21876 11240 21925 11268
rect 21876 11228 21882 11240
rect 21913 11237 21925 11240
rect 21959 11237 21971 11271
rect 23198 11268 23204 11280
rect 23159 11240 23204 11268
rect 21913 11231 21971 11237
rect 23198 11228 23204 11240
rect 23256 11268 23262 11280
rect 24121 11271 24179 11277
rect 24121 11268 24133 11271
rect 23256 11240 24133 11268
rect 23256 11228 23262 11240
rect 24121 11237 24133 11240
rect 24167 11237 24179 11271
rect 24121 11231 24179 11237
rect 20990 11200 20996 11212
rect 18279 11172 20529 11200
rect 20951 11172 20996 11200
rect 18279 11169 18291 11172
rect 18233 11163 18291 11169
rect 20990 11160 20996 11172
rect 21048 11160 21054 11212
rect 21266 11160 21272 11212
rect 21324 11200 21330 11212
rect 21361 11203 21419 11209
rect 21361 11200 21373 11203
rect 21324 11172 21373 11200
rect 21324 11160 21330 11172
rect 21361 11169 21373 11172
rect 21407 11169 21419 11203
rect 21361 11163 21419 11169
rect 24648 11203 24706 11209
rect 24648 11169 24660 11203
rect 24694 11200 24706 11203
rect 24762 11200 24768 11212
rect 24694 11172 24768 11200
rect 24694 11169 24706 11172
rect 24648 11163 24706 11169
rect 24762 11160 24768 11172
rect 24820 11160 24826 11212
rect 11388 11104 11646 11132
rect 13357 11135 13415 11141
rect 11388 11092 11394 11104
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 13814 11132 13820 11144
rect 13403 11104 13820 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 13814 11092 13820 11104
rect 13872 11132 13878 11144
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 13872 11104 14565 11132
rect 13872 11092 13878 11104
rect 14553 11101 14565 11104
rect 14599 11101 14611 11135
rect 14553 11095 14611 11101
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11101 15439 11135
rect 15746 11132 15752 11144
rect 15707 11104 15752 11132
rect 15381 11095 15439 11101
rect 11882 11024 11888 11076
rect 11940 11064 11946 11076
rect 15286 11064 15292 11076
rect 11940 11036 15292 11064
rect 11940 11024 11946 11036
rect 15286 11024 15292 11036
rect 15344 11024 15350 11076
rect 15396 11064 15424 11095
rect 15746 11092 15752 11104
rect 15804 11132 15810 11144
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 15804 11104 16681 11132
rect 15804 11092 15810 11104
rect 16669 11101 16681 11104
rect 16715 11101 16727 11135
rect 19058 11132 19064 11144
rect 19019 11104 19064 11132
rect 16669 11095 16727 11101
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 20346 11092 20352 11144
rect 20404 11132 20410 11144
rect 20625 11135 20683 11141
rect 20625 11132 20637 11135
rect 20404 11104 20637 11132
rect 20404 11092 20410 11104
rect 20625 11101 20637 11104
rect 20671 11101 20683 11135
rect 23106 11132 23112 11144
rect 23067 11104 23112 11132
rect 20625 11095 20683 11101
rect 23106 11092 23112 11104
rect 23164 11132 23170 11144
rect 25130 11132 25136 11144
rect 23164 11104 25136 11132
rect 23164 11092 23170 11104
rect 25130 11092 25136 11104
rect 25188 11092 25194 11144
rect 15396 11036 16436 11064
rect 16408 11008 16436 11036
rect 22646 11024 22652 11076
rect 22704 11064 22710 11076
rect 23661 11067 23719 11073
rect 23661 11064 23673 11067
rect 22704 11036 23673 11064
rect 22704 11024 22710 11036
rect 23661 11033 23673 11036
rect 23707 11064 23719 11067
rect 24026 11064 24032 11076
rect 23707 11036 24032 11064
rect 23707 11033 23719 11036
rect 23661 11027 23719 11033
rect 24026 11024 24032 11036
rect 24084 11024 24090 11076
rect 9401 10999 9459 11005
rect 9401 10996 9413 10999
rect 8812 10968 9413 10996
rect 8812 10956 8818 10968
rect 9401 10965 9413 10968
rect 9447 10965 9459 10999
rect 9401 10959 9459 10965
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 12897 10999 12955 11005
rect 12897 10996 12909 10999
rect 12768 10968 12909 10996
rect 12768 10956 12774 10968
rect 12897 10965 12909 10968
rect 12943 10965 12955 10999
rect 16390 10996 16396 11008
rect 16351 10968 16396 10996
rect 12897 10959 12955 10965
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 18782 10956 18788 11008
rect 18840 10996 18846 11008
rect 18877 10999 18935 11005
rect 18877 10996 18889 10999
rect 18840 10968 18889 10996
rect 18840 10956 18846 10968
rect 18877 10965 18889 10968
rect 18923 10965 18935 10999
rect 18877 10959 18935 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1762 10792 1768 10804
rect 1723 10764 1768 10792
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 1946 10752 1952 10804
rect 2004 10792 2010 10804
rect 2041 10795 2099 10801
rect 2041 10792 2053 10795
rect 2004 10764 2053 10792
rect 2004 10752 2010 10764
rect 2041 10761 2053 10764
rect 2087 10792 2099 10795
rect 2498 10792 2504 10804
rect 2087 10764 2504 10792
rect 2087 10761 2099 10764
rect 2041 10755 2099 10761
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 4246 10792 4252 10804
rect 4207 10764 4252 10792
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 5258 10752 5264 10804
rect 5316 10792 5322 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 5316 10764 5457 10792
rect 5316 10752 5322 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 6178 10792 6184 10804
rect 6139 10764 6184 10792
rect 5445 10755 5503 10761
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 7929 10795 7987 10801
rect 7929 10761 7941 10795
rect 7975 10792 7987 10795
rect 8294 10792 8300 10804
rect 7975 10764 8300 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 9861 10795 9919 10801
rect 9861 10761 9873 10795
rect 9907 10792 9919 10795
rect 10134 10792 10140 10804
rect 9907 10764 10140 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 10134 10752 10140 10764
rect 10192 10792 10198 10804
rect 11241 10795 11299 10801
rect 11241 10792 11253 10795
rect 10192 10764 11253 10792
rect 10192 10752 10198 10764
rect 11241 10761 11253 10764
rect 11287 10761 11299 10795
rect 12618 10792 12624 10804
rect 12579 10764 12624 10792
rect 11241 10755 11299 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 13722 10792 13728 10804
rect 13683 10764 13728 10792
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 15654 10752 15660 10804
rect 15712 10792 15718 10804
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 15712 10764 17141 10792
rect 15712 10752 15718 10764
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 17589 10795 17647 10801
rect 17589 10761 17601 10795
rect 17635 10792 17647 10795
rect 17770 10792 17776 10804
rect 17635 10764 17776 10792
rect 17635 10761 17647 10764
rect 17589 10755 17647 10761
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 22741 10795 22799 10801
rect 22741 10761 22753 10795
rect 22787 10792 22799 10795
rect 23106 10792 23112 10804
rect 22787 10764 23112 10792
rect 22787 10761 22799 10764
rect 22741 10755 22799 10761
rect 23106 10752 23112 10764
rect 23164 10752 23170 10804
rect 23477 10795 23535 10801
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 23566 10792 23572 10804
rect 23523 10764 23572 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 23566 10752 23572 10764
rect 23624 10752 23630 10804
rect 25406 10792 25412 10804
rect 25367 10764 25412 10792
rect 25406 10752 25412 10764
rect 25464 10752 25470 10804
rect 5276 10724 5304 10752
rect 4816 10696 5304 10724
rect 7193 10727 7251 10733
rect 2958 10656 2964 10668
rect 2919 10628 2964 10656
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 4709 10591 4767 10597
rect 4709 10588 4721 10591
rect 4672 10560 4721 10588
rect 4672 10548 4678 10560
rect 4709 10557 4721 10560
rect 4755 10588 4767 10591
rect 4816 10588 4844 10696
rect 7193 10693 7205 10727
rect 7239 10724 7251 10727
rect 11054 10724 11060 10736
rect 7239 10696 11060 10724
rect 7239 10693 7251 10696
rect 7193 10687 7251 10693
rect 11054 10684 11060 10696
rect 11112 10684 11118 10736
rect 15013 10727 15071 10733
rect 15013 10693 15025 10727
rect 15059 10724 15071 10727
rect 15197 10727 15255 10733
rect 15197 10724 15209 10727
rect 15059 10696 15209 10724
rect 15059 10693 15071 10696
rect 15013 10687 15071 10693
rect 15197 10693 15209 10696
rect 15243 10724 15255 10727
rect 15378 10724 15384 10736
rect 15243 10696 15384 10724
rect 15243 10693 15255 10696
rect 15197 10687 15255 10693
rect 15378 10684 15384 10696
rect 15436 10684 15442 10736
rect 16209 10727 16267 10733
rect 16209 10693 16221 10727
rect 16255 10724 16267 10727
rect 16942 10724 16948 10736
rect 16255 10696 16948 10724
rect 16255 10693 16267 10696
rect 16209 10687 16267 10693
rect 16942 10684 16948 10696
rect 17000 10684 17006 10736
rect 19058 10684 19064 10736
rect 19116 10724 19122 10736
rect 20073 10727 20131 10733
rect 20073 10724 20085 10727
rect 19116 10696 20085 10724
rect 19116 10684 19122 10696
rect 20073 10693 20085 10696
rect 20119 10724 20131 10727
rect 22186 10724 22192 10736
rect 20119 10696 22192 10724
rect 20119 10693 20131 10696
rect 20073 10687 20131 10693
rect 22186 10684 22192 10696
rect 22244 10684 22250 10736
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10656 5227 10659
rect 5442 10656 5448 10668
rect 5215 10628 5448 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 6454 10616 6460 10668
rect 6512 10656 6518 10668
rect 7561 10659 7619 10665
rect 7561 10656 7573 10659
rect 6512 10628 7573 10656
rect 6512 10616 6518 10628
rect 7561 10625 7573 10628
rect 7607 10656 7619 10659
rect 8570 10656 8576 10668
rect 7607 10628 8576 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 13449 10659 13507 10665
rect 13449 10625 13461 10659
rect 13495 10656 13507 10659
rect 20438 10656 20444 10668
rect 13495 10628 20444 10656
rect 13495 10625 13507 10628
rect 13449 10619 13507 10625
rect 20438 10616 20444 10628
rect 20496 10616 20502 10668
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10656 21327 10659
rect 21358 10656 21364 10668
rect 21315 10628 21364 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 23109 10659 23167 10665
rect 23109 10625 23121 10659
rect 23155 10656 23167 10659
rect 23198 10656 23204 10668
rect 23155 10628 23204 10656
rect 23155 10625 23167 10628
rect 23109 10619 23167 10625
rect 23198 10616 23204 10628
rect 23256 10616 23262 10668
rect 24026 10656 24032 10668
rect 23987 10628 24032 10656
rect 24026 10616 24032 10628
rect 24084 10616 24090 10668
rect 4982 10588 4988 10600
rect 4755 10560 4844 10588
rect 4895 10560 4988 10588
rect 4755 10557 4767 10560
rect 4709 10551 4767 10557
rect 4982 10548 4988 10560
rect 5040 10588 5046 10600
rect 6472 10588 6500 10616
rect 5040 10560 6500 10588
rect 7009 10591 7067 10597
rect 5040 10548 5046 10560
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 2317 10523 2375 10529
rect 2317 10489 2329 10523
rect 2363 10489 2375 10523
rect 2317 10483 2375 10489
rect 2409 10523 2467 10529
rect 2409 10489 2421 10523
rect 2455 10520 2467 10523
rect 2498 10520 2504 10532
rect 2455 10492 2504 10520
rect 2455 10489 2467 10492
rect 2409 10483 2467 10489
rect 2222 10412 2228 10464
rect 2280 10452 2286 10464
rect 2332 10452 2360 10483
rect 2498 10480 2504 10492
rect 2556 10480 2562 10532
rect 3605 10523 3663 10529
rect 3605 10489 3617 10523
rect 3651 10520 3663 10523
rect 3881 10523 3939 10529
rect 3881 10520 3893 10523
rect 3651 10492 3893 10520
rect 3651 10489 3663 10492
rect 3605 10483 3663 10489
rect 3881 10489 3893 10492
rect 3927 10520 3939 10523
rect 5000 10520 5028 10548
rect 3927 10492 5028 10520
rect 6641 10523 6699 10529
rect 3927 10489 3939 10492
rect 3881 10483 3939 10489
rect 6641 10489 6653 10523
rect 6687 10520 6699 10523
rect 7024 10520 7052 10551
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 8665 10591 8723 10597
rect 8665 10588 8677 10591
rect 8260 10560 8677 10588
rect 8260 10548 8266 10560
rect 8665 10557 8677 10560
rect 8711 10588 8723 10591
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 8711 10560 9045 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 9033 10557 9045 10560
rect 9079 10588 9091 10591
rect 9122 10588 9128 10600
rect 9079 10560 9128 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9493 10591 9551 10597
rect 9493 10557 9505 10591
rect 9539 10588 9551 10591
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 9539 10560 10333 10588
rect 9539 10557 9551 10560
rect 9493 10551 9551 10557
rect 10321 10557 10333 10560
rect 10367 10588 10379 10591
rect 10778 10588 10784 10600
rect 10367 10560 10784 10588
rect 10367 10557 10379 10560
rect 10321 10551 10379 10557
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 12768 10560 13093 10588
rect 12768 10548 12774 10560
rect 13081 10557 13093 10560
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 15105 10591 15163 10597
rect 15105 10588 15117 10591
rect 14875 10560 15117 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 15105 10557 15117 10560
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 15381 10591 15439 10597
rect 15381 10557 15393 10591
rect 15427 10588 15439 10591
rect 15470 10588 15476 10600
rect 15427 10560 15476 10588
rect 15427 10557 15439 10560
rect 15381 10551 15439 10557
rect 9858 10520 9864 10532
rect 6687 10492 9864 10520
rect 6687 10489 6699 10492
rect 6641 10483 6699 10489
rect 9858 10480 9864 10492
rect 9916 10480 9922 10532
rect 10229 10523 10287 10529
rect 10229 10489 10241 10523
rect 10275 10520 10287 10523
rect 10683 10523 10741 10529
rect 10683 10520 10695 10523
rect 10275 10492 10695 10520
rect 10275 10489 10287 10492
rect 10229 10483 10287 10489
rect 10683 10489 10695 10492
rect 10729 10520 10741 10523
rect 11238 10520 11244 10532
rect 10729 10492 11244 10520
rect 10729 10489 10741 10492
rect 10683 10483 10741 10489
rect 8294 10452 8300 10464
rect 2280 10424 2360 10452
rect 8255 10424 8300 10452
rect 2280 10412 2286 10424
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 10244 10452 10272 10483
rect 11238 10480 11244 10492
rect 11296 10480 11302 10532
rect 11330 10480 11336 10532
rect 11388 10520 11394 10532
rect 12161 10523 12219 10529
rect 12161 10520 12173 10523
rect 11388 10492 12173 10520
rect 11388 10480 11394 10492
rect 12161 10489 12173 10492
rect 12207 10520 12219 10523
rect 12894 10520 12900 10532
rect 12207 10492 12900 10520
rect 12207 10489 12219 10492
rect 12161 10483 12219 10489
rect 12894 10480 12900 10492
rect 12952 10480 12958 10532
rect 14277 10523 14335 10529
rect 14277 10489 14289 10523
rect 14323 10520 14335 10523
rect 15396 10520 15424 10551
rect 15470 10548 15476 10560
rect 15528 10548 15534 10600
rect 16945 10591 17003 10597
rect 16945 10557 16957 10591
rect 16991 10557 17003 10591
rect 16945 10551 17003 10557
rect 14323 10492 15424 10520
rect 14323 10489 14335 10492
rect 14277 10483 14335 10489
rect 8720 10424 10272 10452
rect 8720 10412 8726 10424
rect 10870 10412 10876 10464
rect 10928 10452 10934 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 10928 10424 11529 10452
rect 10928 10412 10934 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 11517 10415 11575 10421
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 14553 10455 14611 10461
rect 14553 10452 14565 10455
rect 14240 10424 14565 10452
rect 14240 10412 14246 10424
rect 14553 10421 14565 10424
rect 14599 10452 14611 10455
rect 14829 10455 14887 10461
rect 14829 10452 14841 10455
rect 14599 10424 14841 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 14829 10421 14841 10424
rect 14875 10421 14887 10455
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 14829 10415 14887 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 16853 10455 16911 10461
rect 16853 10421 16865 10455
rect 16899 10452 16911 10455
rect 16960 10452 16988 10551
rect 18874 10548 18880 10600
rect 18932 10588 18938 10600
rect 18969 10591 19027 10597
rect 18969 10588 18981 10591
rect 18932 10560 18981 10588
rect 18932 10548 18938 10560
rect 18969 10557 18981 10560
rect 19015 10557 19027 10591
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 18969 10551 19027 10557
rect 19352 10560 19441 10588
rect 19352 10532 19380 10560
rect 19429 10557 19441 10560
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 25225 10591 25283 10597
rect 25225 10557 25237 10591
rect 25271 10557 25283 10591
rect 25225 10551 25283 10557
rect 18509 10523 18567 10529
rect 18509 10489 18521 10523
rect 18555 10520 18567 10523
rect 19334 10520 19340 10532
rect 18555 10492 19340 10520
rect 18555 10489 18567 10492
rect 18509 10483 18567 10489
rect 19334 10480 19340 10492
rect 19392 10480 19398 10532
rect 19705 10523 19763 10529
rect 19705 10489 19717 10523
rect 19751 10520 19763 10523
rect 20162 10520 20168 10532
rect 19751 10492 20168 10520
rect 19751 10489 19763 10492
rect 19705 10483 19763 10489
rect 20162 10480 20168 10492
rect 20220 10480 20226 10532
rect 21266 10520 21272 10532
rect 20548 10492 21272 10520
rect 17218 10452 17224 10464
rect 16899 10424 17224 10452
rect 16899 10421 16911 10424
rect 16853 10415 16911 10421
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 18782 10452 18788 10464
rect 18743 10424 18788 10452
rect 18782 10412 18788 10424
rect 18840 10412 18846 10464
rect 19242 10412 19248 10464
rect 19300 10452 19306 10464
rect 20548 10461 20576 10492
rect 21266 10480 21272 10492
rect 21324 10480 21330 10532
rect 21361 10523 21419 10529
rect 21361 10489 21373 10523
rect 21407 10489 21419 10523
rect 21910 10520 21916 10532
rect 21871 10492 21916 10520
rect 21361 10483 21419 10489
rect 20533 10455 20591 10461
rect 20533 10452 20545 10455
rect 19300 10424 20545 10452
rect 19300 10412 19306 10424
rect 20533 10421 20545 10424
rect 20579 10421 20591 10455
rect 20990 10452 20996 10464
rect 20951 10424 20996 10452
rect 20533 10415 20591 10421
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 21082 10412 21088 10464
rect 21140 10452 21146 10464
rect 21376 10452 21404 10483
rect 21910 10480 21916 10492
rect 21968 10480 21974 10532
rect 23750 10520 23756 10532
rect 23711 10492 23756 10520
rect 23750 10480 23756 10492
rect 23808 10480 23814 10532
rect 23845 10523 23903 10529
rect 23845 10489 23857 10523
rect 23891 10489 23903 10523
rect 23845 10483 23903 10489
rect 22189 10455 22247 10461
rect 22189 10452 22201 10455
rect 21140 10424 22201 10452
rect 21140 10412 21146 10424
rect 22189 10421 22201 10424
rect 22235 10421 22247 10455
rect 22189 10415 22247 10421
rect 23566 10412 23572 10464
rect 23624 10452 23630 10464
rect 23860 10452 23888 10483
rect 24026 10480 24032 10532
rect 24084 10520 24090 10532
rect 25240 10520 25268 10551
rect 25685 10523 25743 10529
rect 25685 10520 25697 10523
rect 24084 10492 25697 10520
rect 24084 10480 24090 10492
rect 25685 10489 25697 10492
rect 25731 10489 25743 10523
rect 25685 10483 25743 10489
rect 24762 10452 24768 10464
rect 23624 10424 23888 10452
rect 24723 10424 24768 10452
rect 23624 10412 23630 10424
rect 24762 10412 24768 10424
rect 24820 10412 24826 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1535 10251 1593 10257
rect 1535 10217 1547 10251
rect 1581 10248 1593 10251
rect 1854 10248 1860 10260
rect 1581 10220 1860 10248
rect 1581 10217 1593 10220
rect 1535 10211 1593 10217
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 2314 10208 2320 10260
rect 2372 10248 2378 10260
rect 2547 10251 2605 10257
rect 2547 10248 2559 10251
rect 2372 10220 2559 10248
rect 2372 10208 2378 10220
rect 2547 10217 2559 10220
rect 2593 10217 2605 10251
rect 4430 10248 4436 10260
rect 4391 10220 4436 10248
rect 2547 10211 2605 10217
rect 4430 10208 4436 10220
rect 4488 10208 4494 10260
rect 6086 10208 6092 10260
rect 6144 10248 6150 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 6144 10220 6193 10248
rect 6144 10208 6150 10220
rect 6181 10217 6193 10220
rect 6227 10248 6239 10251
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 6227 10220 6929 10248
rect 6227 10217 6239 10220
rect 6181 10211 6239 10217
rect 6917 10217 6929 10220
rect 6963 10217 6975 10251
rect 10778 10248 10784 10260
rect 10739 10220 10784 10248
rect 6917 10211 6975 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13688 10220 13921 10248
rect 13688 10208 13694 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 13909 10211 13967 10217
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15344 10220 21541 10248
rect 15344 10208 15350 10220
rect 8202 10180 8208 10192
rect 8163 10152 8208 10180
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 10597 10183 10655 10189
rect 10597 10149 10609 10183
rect 10643 10180 10655 10183
rect 14182 10180 14188 10192
rect 10643 10152 14188 10180
rect 10643 10149 10655 10152
rect 10597 10143 10655 10149
rect 1302 10072 1308 10124
rect 1360 10112 1366 10124
rect 1432 10115 1490 10121
rect 1432 10112 1444 10115
rect 1360 10084 1444 10112
rect 1360 10072 1366 10084
rect 1432 10081 1444 10084
rect 1478 10081 1490 10115
rect 1432 10075 1490 10081
rect 2476 10115 2534 10121
rect 2476 10081 2488 10115
rect 2522 10112 2534 10115
rect 3326 10112 3332 10124
rect 2522 10084 3332 10112
rect 2522 10081 2534 10084
rect 2476 10075 2534 10081
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 3970 10072 3976 10124
rect 4028 10112 4034 10124
rect 4614 10112 4620 10124
rect 4028 10084 4620 10112
rect 4028 10072 4034 10084
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 4893 10115 4951 10121
rect 4893 10081 4905 10115
rect 4939 10112 4951 10115
rect 5166 10112 5172 10124
rect 4939 10084 5172 10112
rect 4939 10081 4951 10084
rect 4893 10075 4951 10081
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 6270 10112 6276 10124
rect 6227 10084 6276 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6454 10112 6460 10124
rect 6415 10084 6460 10112
rect 6454 10072 6460 10084
rect 6512 10072 6518 10124
rect 9728 10115 9786 10121
rect 9728 10081 9740 10115
rect 9774 10112 9786 10115
rect 10134 10112 10140 10124
rect 9774 10084 10140 10112
rect 9774 10081 9786 10084
rect 9728 10075 9786 10081
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10686 10112 10692 10124
rect 10647 10084 10692 10112
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 10870 10072 10876 10124
rect 10928 10112 10934 10124
rect 11149 10115 11207 10121
rect 11149 10112 11161 10115
rect 10928 10084 11161 10112
rect 10928 10072 10934 10084
rect 11149 10081 11161 10084
rect 11195 10081 11207 10115
rect 11606 10112 11612 10124
rect 11567 10084 11612 10112
rect 11149 10075 11207 10081
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 11900 10121 11928 10152
rect 11885 10115 11943 10121
rect 11885 10081 11897 10115
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 12710 10072 12716 10124
rect 12768 10112 12774 10124
rect 13786 10121 13814 10152
rect 14182 10140 14188 10152
rect 14240 10140 14246 10192
rect 16850 10140 16856 10192
rect 16908 10180 16914 10192
rect 17266 10183 17324 10189
rect 17266 10180 17278 10183
rect 16908 10152 17278 10180
rect 16908 10140 16914 10152
rect 17266 10149 17278 10152
rect 17312 10180 17324 10183
rect 18782 10180 18788 10192
rect 17312 10152 18788 10180
rect 17312 10149 17324 10152
rect 17266 10143 17324 10149
rect 18782 10140 18788 10152
rect 18840 10140 18846 10192
rect 21174 10180 21180 10192
rect 21135 10152 21180 10180
rect 21174 10140 21180 10152
rect 21232 10140 21238 10192
rect 21513 10180 21541 10220
rect 21910 10208 21916 10260
rect 21968 10248 21974 10260
rect 22097 10251 22155 10257
rect 22097 10248 22109 10251
rect 21968 10220 22109 10248
rect 21968 10208 21974 10220
rect 22097 10217 22109 10220
rect 22143 10217 22155 10251
rect 22097 10211 22155 10217
rect 22186 10208 22192 10260
rect 22244 10248 22250 10260
rect 22741 10251 22799 10257
rect 22741 10248 22753 10251
rect 22244 10220 22753 10248
rect 22244 10208 22250 10220
rect 22741 10217 22753 10220
rect 22787 10217 22799 10251
rect 23750 10248 23756 10260
rect 23711 10220 23756 10248
rect 22741 10211 22799 10217
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 24118 10208 24124 10260
rect 24176 10248 24182 10260
rect 24351 10251 24409 10257
rect 24351 10248 24363 10251
rect 24176 10220 24363 10248
rect 24176 10208 24182 10220
rect 24351 10217 24363 10220
rect 24397 10217 24409 10251
rect 24351 10211 24409 10217
rect 25222 10208 25228 10260
rect 25280 10248 25286 10260
rect 25363 10251 25421 10257
rect 25363 10248 25375 10251
rect 25280 10220 25375 10248
rect 25280 10208 25286 10220
rect 25363 10217 25375 10220
rect 25409 10217 25421 10251
rect 25363 10211 25421 10217
rect 22370 10180 22376 10192
rect 21513 10152 22376 10180
rect 22370 10140 22376 10152
rect 22428 10140 22434 10192
rect 12989 10115 13047 10121
rect 12989 10112 13001 10115
rect 12768 10084 13001 10112
rect 12768 10072 12774 10084
rect 12989 10081 13001 10084
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10081 13507 10115
rect 13449 10075 13507 10081
rect 13771 10115 13829 10121
rect 13771 10081 13783 10115
rect 13817 10081 13829 10115
rect 13771 10075 13829 10081
rect 14921 10115 14979 10121
rect 14921 10081 14933 10115
rect 14967 10112 14979 10115
rect 15197 10115 15255 10121
rect 15197 10112 15209 10115
rect 14967 10084 15209 10112
rect 14967 10081 14979 10084
rect 14921 10075 14979 10081
rect 15197 10081 15209 10084
rect 15243 10081 15255 10115
rect 15378 10112 15384 10124
rect 15339 10084 15384 10112
rect 15197 10075 15255 10081
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 7984 10016 8125 10044
rect 7984 10004 7990 10016
rect 8113 10013 8125 10016
rect 8159 10044 8171 10047
rect 9815 10047 9873 10053
rect 9815 10044 9827 10047
rect 8159 10016 9827 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 9815 10013 9827 10016
rect 9861 10013 9873 10047
rect 9815 10007 9873 10013
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10044 10287 10047
rect 10888 10044 10916 10072
rect 10275 10016 10916 10044
rect 11624 10044 11652 10072
rect 13464 10044 13492 10075
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 15470 10072 15476 10124
rect 15528 10112 15534 10124
rect 15565 10115 15623 10121
rect 15565 10112 15577 10115
rect 15528 10084 15577 10112
rect 15528 10072 15534 10084
rect 15565 10081 15577 10084
rect 15611 10081 15623 10115
rect 19242 10112 19248 10124
rect 19203 10084 19248 10112
rect 15565 10075 15623 10081
rect 19242 10072 19248 10084
rect 19300 10072 19306 10124
rect 19334 10072 19340 10124
rect 19392 10112 19398 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19392 10084 19717 10112
rect 19392 10072 19398 10084
rect 19705 10081 19717 10084
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 20990 10072 20996 10124
rect 21048 10112 21054 10124
rect 22922 10112 22928 10124
rect 21048 10084 22928 10112
rect 21048 10072 21054 10084
rect 22922 10072 22928 10084
rect 22980 10072 22986 10124
rect 23106 10112 23112 10124
rect 23067 10084 23112 10112
rect 23106 10072 23112 10084
rect 23164 10112 23170 10124
rect 24026 10112 24032 10124
rect 23164 10084 24032 10112
rect 23164 10072 23170 10084
rect 24026 10072 24032 10084
rect 24084 10072 24090 10124
rect 24248 10115 24306 10121
rect 24248 10081 24260 10115
rect 24294 10081 24306 10115
rect 24248 10075 24306 10081
rect 25225 10115 25283 10121
rect 25225 10081 25237 10115
rect 25271 10112 25283 10115
rect 25314 10112 25320 10124
rect 25271 10084 25320 10112
rect 25271 10081 25283 10084
rect 25225 10075 25283 10081
rect 11624 10016 13492 10044
rect 14737 10047 14795 10053
rect 10275 10013 10287 10016
rect 10229 10007 10287 10013
rect 14737 10013 14749 10047
rect 14783 10044 14795 10047
rect 15488 10044 15516 10072
rect 16022 10044 16028 10056
rect 14783 10016 15516 10044
rect 15983 10016 16028 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 16942 10044 16948 10056
rect 16903 10016 16948 10044
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 19978 10044 19984 10056
rect 19939 10016 19984 10044
rect 19978 10004 19984 10016
rect 20036 10004 20042 10056
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20772 10016 20913 10044
rect 20772 10004 20778 10016
rect 20901 10013 20913 10016
rect 20947 10013 20959 10047
rect 24118 10044 24124 10056
rect 20901 10007 20959 10013
rect 23446 10016 24124 10044
rect 8665 9979 8723 9985
rect 8665 9945 8677 9979
rect 8711 9976 8723 9979
rect 8754 9976 8760 9988
rect 8711 9948 8760 9976
rect 8711 9945 8723 9948
rect 8665 9939 8723 9945
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 17218 9936 17224 9988
rect 17276 9976 17282 9988
rect 17954 9976 17960 9988
rect 17276 9948 17960 9976
rect 17276 9936 17282 9948
rect 17954 9936 17960 9948
rect 18012 9976 18018 9988
rect 18141 9979 18199 9985
rect 18141 9976 18153 9979
rect 18012 9948 18153 9976
rect 18012 9936 18018 9948
rect 18141 9945 18153 9948
rect 18187 9945 18199 9979
rect 18141 9939 18199 9945
rect 22278 9936 22284 9988
rect 22336 9976 22342 9988
rect 23446 9976 23474 10016
rect 24118 10004 24124 10016
rect 24176 10044 24182 10056
rect 24263 10044 24291 10075
rect 25314 10072 25320 10084
rect 25372 10072 25378 10124
rect 24176 10016 24291 10044
rect 24176 10004 24182 10016
rect 22336 9948 23474 9976
rect 22336 9936 22342 9948
rect 2222 9908 2228 9920
rect 2183 9880 2228 9908
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 2866 9908 2872 9920
rect 2827 9880 2872 9908
rect 2866 9868 2872 9880
rect 2924 9868 2930 9920
rect 9125 9911 9183 9917
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9214 9908 9220 9920
rect 9171 9880 9220 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 9490 9908 9496 9920
rect 9451 9880 9496 9908
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 12710 9908 12716 9920
rect 12671 9880 12716 9908
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 14921 9911 14979 9917
rect 14921 9908 14933 9911
rect 14792 9880 14933 9908
rect 14792 9868 14798 9880
rect 14921 9877 14933 9880
rect 14967 9908 14979 9911
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14967 9880 15025 9908
rect 14967 9877 14979 9880
rect 14921 9871 14979 9877
rect 15013 9877 15025 9880
rect 15059 9877 15071 9911
rect 15013 9871 15071 9877
rect 15838 9868 15844 9920
rect 15896 9908 15902 9920
rect 16301 9911 16359 9917
rect 16301 9908 16313 9911
rect 15896 9880 16313 9908
rect 15896 9868 15902 9880
rect 16301 9877 16313 9880
rect 16347 9877 16359 9911
rect 17862 9908 17868 9920
rect 17823 9880 17868 9908
rect 16301 9871 16359 9877
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 18874 9868 18880 9920
rect 18932 9908 18938 9920
rect 18969 9911 19027 9917
rect 18969 9908 18981 9911
rect 18932 9880 18981 9908
rect 18932 9868 18938 9880
rect 18969 9877 18981 9880
rect 19015 9877 19027 9911
rect 18969 9871 19027 9877
rect 20717 9911 20775 9917
rect 20717 9877 20729 9911
rect 20763 9908 20775 9911
rect 21358 9908 21364 9920
rect 20763 9880 21364 9908
rect 20763 9877 20775 9880
rect 20717 9871 20775 9877
rect 21358 9868 21364 9880
rect 21416 9868 21422 9920
rect 21818 9908 21824 9920
rect 21779 9880 21824 9908
rect 21818 9868 21824 9880
rect 21876 9868 21882 9920
rect 23382 9868 23388 9920
rect 23440 9908 23446 9920
rect 23750 9908 23756 9920
rect 23440 9880 23756 9908
rect 23440 9868 23446 9880
rect 23750 9868 23756 9880
rect 23808 9868 23814 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1302 9664 1308 9716
rect 1360 9704 1366 9716
rect 1857 9707 1915 9713
rect 1857 9704 1869 9707
rect 1360 9676 1869 9704
rect 1360 9664 1366 9676
rect 1857 9673 1869 9676
rect 1903 9673 1915 9707
rect 3326 9704 3332 9716
rect 3287 9676 3332 9704
rect 1857 9667 1915 9673
rect 3326 9664 3332 9676
rect 3384 9664 3390 9716
rect 3970 9704 3976 9716
rect 3931 9676 3976 9704
rect 3970 9664 3976 9676
rect 4028 9664 4034 9716
rect 4341 9707 4399 9713
rect 4341 9673 4353 9707
rect 4387 9704 4399 9707
rect 5166 9704 5172 9716
rect 4387 9676 5172 9704
rect 4387 9673 4399 9676
rect 4341 9667 4399 9673
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 5859 9707 5917 9713
rect 5859 9704 5871 9707
rect 5592 9676 5871 9704
rect 5592 9664 5598 9676
rect 5859 9673 5871 9676
rect 5905 9673 5917 9707
rect 5859 9667 5917 9673
rect 6178 9664 6184 9716
rect 6236 9704 6242 9716
rect 6549 9707 6607 9713
rect 6549 9704 6561 9707
rect 6236 9676 6561 9704
rect 6236 9664 6242 9676
rect 6549 9673 6561 9676
rect 6595 9673 6607 9707
rect 6549 9667 6607 9673
rect 7745 9707 7803 9713
rect 7745 9673 7757 9707
rect 7791 9704 7803 9707
rect 8202 9704 8208 9716
rect 7791 9676 8208 9704
rect 7791 9673 7803 9676
rect 7745 9667 7803 9673
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 9122 9704 9128 9716
rect 9083 9676 9128 9704
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 9766 9704 9772 9716
rect 9679 9676 9772 9704
rect 9766 9664 9772 9676
rect 9824 9704 9830 9716
rect 10134 9704 10140 9716
rect 9824 9676 10140 9704
rect 9824 9664 9830 9676
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 15378 9704 15384 9716
rect 13872 9676 13917 9704
rect 15339 9676 15384 9704
rect 13872 9664 13878 9676
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 17497 9707 17555 9713
rect 17497 9673 17509 9707
rect 17543 9704 17555 9707
rect 17862 9704 17868 9716
rect 17543 9676 17868 9704
rect 17543 9673 17555 9676
rect 17497 9667 17555 9673
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 18506 9704 18512 9716
rect 18419 9676 18512 9704
rect 18506 9664 18512 9676
rect 18564 9704 18570 9716
rect 19242 9704 19248 9716
rect 18564 9676 19248 9704
rect 18564 9664 18570 9676
rect 19242 9664 19248 9676
rect 19300 9704 19306 9716
rect 19613 9707 19671 9713
rect 19613 9704 19625 9707
rect 19300 9676 19625 9704
rect 19300 9664 19306 9676
rect 19613 9673 19625 9676
rect 19659 9673 19671 9707
rect 21082 9704 21088 9716
rect 21043 9676 21088 9704
rect 19613 9667 19671 9673
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 21836 9676 22140 9704
rect 106 9596 112 9648
rect 164 9636 170 9648
rect 1535 9639 1593 9645
rect 164 9608 1507 9636
rect 164 9596 170 9608
rect 1479 9568 1507 9608
rect 1535 9605 1547 9639
rect 1581 9636 1593 9639
rect 2130 9636 2136 9648
rect 1581 9608 2136 9636
rect 1581 9605 1593 9608
rect 1535 9599 1593 9605
rect 2130 9596 2136 9608
rect 2188 9636 2194 9648
rect 2866 9636 2872 9648
rect 2188 9608 2872 9636
rect 2188 9596 2194 9608
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 3142 9596 3148 9648
rect 3200 9636 3206 9648
rect 4571 9639 4629 9645
rect 4571 9636 4583 9639
rect 3200 9608 4583 9636
rect 3200 9596 3206 9608
rect 4571 9605 4583 9608
rect 4617 9605 4629 9639
rect 4571 9599 4629 9605
rect 6273 9639 6331 9645
rect 6273 9605 6285 9639
rect 6319 9636 6331 9639
rect 7650 9636 7656 9648
rect 6319 9608 7656 9636
rect 6319 9605 6331 9608
rect 6273 9599 6331 9605
rect 2225 9571 2283 9577
rect 2225 9568 2237 9571
rect 1479 9540 2237 9568
rect 1479 9509 1507 9540
rect 2225 9537 2237 9540
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 3108 9540 3433 9568
rect 3108 9528 3114 9540
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 1464 9503 1522 9509
rect 1464 9469 1476 9503
rect 1510 9469 1522 9503
rect 1464 9463 1522 9469
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2444 9503 2502 9509
rect 2444 9500 2456 9503
rect 2096 9472 2456 9500
rect 2096 9460 2102 9472
rect 2444 9469 2456 9472
rect 2490 9500 2502 9503
rect 2869 9503 2927 9509
rect 2869 9500 2881 9503
rect 2490 9472 2881 9500
rect 2490 9469 2502 9472
rect 2444 9463 2502 9469
rect 2869 9469 2881 9472
rect 2915 9469 2927 9503
rect 2869 9463 2927 9469
rect 4500 9503 4558 9509
rect 4500 9469 4512 9503
rect 4546 9500 4558 9503
rect 5788 9503 5846 9509
rect 4546 9472 5028 9500
rect 4546 9469 4558 9472
rect 4500 9463 4558 9469
rect 1578 9392 1584 9444
rect 1636 9432 1642 9444
rect 2547 9435 2605 9441
rect 2547 9432 2559 9435
rect 1636 9404 2559 9432
rect 1636 9392 1642 9404
rect 2547 9401 2559 9404
rect 2593 9401 2605 9435
rect 2547 9395 2605 9401
rect 5000 9373 5028 9472
rect 5788 9469 5800 9503
rect 5834 9500 5846 9503
rect 6288 9500 6316 9599
rect 7650 9596 7656 9608
rect 7708 9596 7714 9648
rect 14458 9636 14464 9648
rect 13832 9608 14464 9636
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9568 7251 9571
rect 10042 9568 10048 9580
rect 7239 9540 10048 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 11330 9568 11336 9580
rect 10796 9540 11336 9568
rect 5834 9472 6316 9500
rect 8205 9503 8263 9509
rect 5834 9469 5846 9472
rect 5788 9463 5846 9469
rect 8205 9469 8217 9503
rect 8251 9500 8263 9503
rect 9214 9500 9220 9512
rect 8251 9472 9220 9500
rect 8251 9469 8263 9472
rect 8205 9463 8263 9469
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 9490 9460 9496 9512
rect 9548 9500 9554 9512
rect 10796 9509 10824 9540
rect 11330 9528 11336 9540
rect 11388 9528 11394 9580
rect 11514 9568 11520 9580
rect 11475 9540 11520 9568
rect 11514 9528 11520 9540
rect 11572 9528 11578 9580
rect 11698 9528 11704 9580
rect 11756 9568 11762 9580
rect 13832 9568 13860 9608
rect 14458 9596 14464 9608
rect 14516 9636 14522 9648
rect 15838 9636 15844 9648
rect 14516 9608 15844 9636
rect 14516 9596 14522 9608
rect 15838 9596 15844 9608
rect 15896 9596 15902 9648
rect 18524 9636 18552 9664
rect 21836 9636 21864 9676
rect 17696 9608 18552 9636
rect 18616 9608 21864 9636
rect 14182 9568 14188 9580
rect 11756 9540 13860 9568
rect 14095 9540 14188 9568
rect 11756 9528 11762 9540
rect 14182 9528 14188 9540
rect 14240 9568 14246 9580
rect 16206 9568 16212 9580
rect 14240 9540 16212 9568
rect 14240 9528 14246 9540
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 16577 9571 16635 9577
rect 16577 9537 16589 9571
rect 16623 9568 16635 9571
rect 16942 9568 16948 9580
rect 16623 9540 16948 9568
rect 16623 9537 16635 9540
rect 16577 9531 16635 9537
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 10781 9503 10839 9509
rect 10781 9500 10793 9503
rect 9548 9472 10793 9500
rect 9548 9460 9554 9472
rect 10781 9469 10793 9472
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 11057 9503 11115 9509
rect 10928 9472 10973 9500
rect 10928 9460 10934 9472
rect 11057 9469 11069 9503
rect 11103 9469 11115 9503
rect 12710 9500 12716 9512
rect 12671 9472 12716 9500
rect 11057 9463 11115 9469
rect 5629 9435 5687 9441
rect 5629 9401 5641 9435
rect 5675 9432 5687 9435
rect 6454 9432 6460 9444
rect 5675 9404 6460 9432
rect 5675 9401 5687 9404
rect 5629 9395 5687 9401
rect 6454 9392 6460 9404
rect 6512 9392 6518 9444
rect 8113 9435 8171 9441
rect 8113 9401 8125 9435
rect 8159 9432 8171 9435
rect 8567 9435 8625 9441
rect 8567 9432 8579 9435
rect 8159 9404 8579 9432
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 8567 9401 8579 9404
rect 8613 9432 8625 9435
rect 8662 9432 8668 9444
rect 8613 9404 8668 9432
rect 8613 9401 8625 9404
rect 8567 9395 8625 9401
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 4985 9367 5043 9373
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 9122 9364 9128 9376
rect 5031 9336 9128 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 10321 9367 10379 9373
rect 10321 9333 10333 9367
rect 10367 9364 10379 9367
rect 10686 9364 10692 9376
rect 10367 9336 10692 9364
rect 10367 9333 10379 9336
rect 10321 9327 10379 9333
rect 10686 9324 10692 9336
rect 10744 9364 10750 9376
rect 11072 9364 11100 9463
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 13541 9503 13599 9509
rect 13541 9469 13553 9503
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 14274 9500 14280 9512
rect 13771 9472 14280 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 10744 9336 11100 9364
rect 10744 9324 10750 9336
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 11885 9367 11943 9373
rect 11885 9364 11897 9367
rect 11664 9336 11897 9364
rect 11664 9324 11670 9336
rect 11885 9333 11897 9336
rect 11931 9364 11943 9367
rect 12250 9364 12256 9376
rect 11931 9336 12256 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 13556 9364 13584 9463
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14516 9472 14841 9500
rect 14516 9460 14522 9472
rect 14829 9469 14841 9472
rect 14875 9500 14887 9503
rect 15562 9500 15568 9512
rect 14875 9472 15568 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 15838 9500 15844 9512
rect 15799 9472 15844 9500
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 15930 9460 15936 9512
rect 15988 9500 15994 9512
rect 16301 9503 16359 9509
rect 16301 9500 16313 9503
rect 15988 9472 16313 9500
rect 15988 9460 15994 9472
rect 16301 9469 16313 9472
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 17696 9432 17724 9608
rect 18616 9580 18644 9608
rect 21910 9596 21916 9648
rect 21968 9636 21974 9648
rect 21968 9608 22048 9636
rect 21968 9596 21974 9608
rect 18598 9568 18604 9580
rect 18559 9540 18604 9568
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 18782 9528 18788 9580
rect 18840 9568 18846 9580
rect 19889 9571 19947 9577
rect 19889 9568 19901 9571
rect 18840 9540 19901 9568
rect 18840 9528 18846 9540
rect 19889 9537 19901 9540
rect 19935 9568 19947 9571
rect 19981 9571 20039 9577
rect 19981 9568 19993 9571
rect 19935 9540 19993 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 19981 9537 19993 9540
rect 20027 9537 20039 9571
rect 20162 9568 20168 9580
rect 20123 9540 20168 9568
rect 19981 9531 20039 9537
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 22020 9577 22048 9608
rect 22005 9571 22063 9577
rect 22005 9537 22017 9571
rect 22051 9537 22063 9571
rect 22112 9568 22140 9676
rect 22922 9664 22928 9716
rect 22980 9704 22986 9716
rect 23293 9707 23351 9713
rect 23293 9704 23305 9707
rect 22980 9676 23305 9704
rect 22980 9664 22986 9676
rect 23293 9673 23305 9676
rect 23339 9673 23351 9707
rect 24118 9704 24124 9716
rect 24079 9676 24124 9704
rect 23293 9667 23351 9673
rect 24118 9664 24124 9676
rect 24176 9664 24182 9716
rect 24581 9707 24639 9713
rect 24581 9673 24593 9707
rect 24627 9704 24639 9707
rect 24670 9704 24676 9716
rect 24627 9676 24676 9704
rect 24627 9673 24639 9676
rect 24581 9667 24639 9673
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 24854 9704 24860 9716
rect 24815 9676 24860 9704
rect 24854 9664 24860 9676
rect 24912 9664 24918 9716
rect 22370 9596 22376 9648
rect 22428 9636 22434 9648
rect 23842 9636 23848 9648
rect 22428 9608 23848 9636
rect 22428 9596 22434 9608
rect 23308 9580 23336 9608
rect 23842 9596 23848 9608
rect 23900 9596 23906 9648
rect 25314 9636 25320 9648
rect 25227 9608 25320 9636
rect 25314 9596 25320 9608
rect 25372 9636 25378 9648
rect 27614 9636 27620 9648
rect 25372 9608 27620 9636
rect 25372 9596 25378 9608
rect 27614 9596 27620 9608
rect 27672 9596 27678 9648
rect 22278 9568 22284 9580
rect 22112 9540 22284 9568
rect 22005 9531 22063 9537
rect 22278 9528 22284 9540
rect 22336 9528 22342 9580
rect 23290 9528 23296 9580
rect 23348 9528 23354 9580
rect 18874 9460 18880 9512
rect 18932 9500 18938 9512
rect 18932 9472 21864 9500
rect 18932 9460 18938 9472
rect 15580 9404 17724 9432
rect 17773 9435 17831 9441
rect 14366 9364 14372 9376
rect 13556 9336 14372 9364
rect 14366 9324 14372 9336
rect 14424 9364 14430 9376
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 14424 9336 14473 9364
rect 14424 9324 14430 9336
rect 14461 9333 14473 9336
rect 14507 9364 14519 9367
rect 14734 9364 14740 9376
rect 14507 9336 14740 9364
rect 14507 9333 14519 9336
rect 14461 9327 14519 9333
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 15013 9367 15071 9373
rect 15013 9333 15025 9367
rect 15059 9364 15071 9367
rect 15580 9364 15608 9404
rect 17773 9401 17785 9435
rect 17819 9432 17831 9435
rect 18138 9432 18144 9444
rect 17819 9404 18144 9432
rect 17819 9401 17831 9404
rect 17773 9395 17831 9401
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9401 18291 9435
rect 18233 9395 18291 9401
rect 19889 9435 19947 9441
rect 19889 9401 19901 9435
rect 19935 9432 19947 9435
rect 20486 9435 20544 9441
rect 20486 9432 20498 9435
rect 19935 9404 20498 9432
rect 19935 9401 19947 9404
rect 19889 9395 19947 9401
rect 20486 9401 20498 9404
rect 20532 9401 20544 9435
rect 20486 9395 20544 9401
rect 15059 9336 15608 9364
rect 15749 9367 15807 9373
rect 15059 9333 15071 9336
rect 15013 9327 15071 9333
rect 15749 9333 15761 9367
rect 15795 9364 15807 9367
rect 15838 9364 15844 9376
rect 15795 9336 15844 9364
rect 15795 9333 15807 9336
rect 15749 9327 15807 9333
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 16945 9367 17003 9373
rect 16945 9364 16957 9367
rect 16908 9336 16957 9364
rect 16908 9324 16914 9336
rect 16945 9333 16957 9336
rect 16991 9333 17003 9367
rect 16945 9327 17003 9333
rect 17862 9324 17868 9376
rect 17920 9364 17926 9376
rect 18248 9364 18276 9395
rect 19242 9364 19248 9376
rect 17920 9336 18276 9364
rect 19203 9336 19248 9364
rect 17920 9324 17926 9336
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 20501 9364 20529 9395
rect 20714 9392 20720 9444
rect 20772 9432 20778 9444
rect 21729 9435 21787 9441
rect 21729 9432 21741 9435
rect 20772 9404 21741 9432
rect 20772 9392 20778 9404
rect 21729 9401 21741 9404
rect 21775 9401 21787 9435
rect 21729 9395 21787 9401
rect 20990 9364 20996 9376
rect 20501 9336 20996 9364
rect 20990 9324 20996 9336
rect 21048 9364 21054 9376
rect 21174 9364 21180 9376
rect 21048 9336 21180 9364
rect 21048 9324 21054 9336
rect 21174 9324 21180 9336
rect 21232 9364 21238 9376
rect 21361 9367 21419 9373
rect 21361 9364 21373 9367
rect 21232 9336 21373 9364
rect 21232 9324 21238 9336
rect 21361 9333 21373 9336
rect 21407 9333 21419 9367
rect 21836 9364 21864 9472
rect 22094 9392 22100 9444
rect 22152 9432 22158 9444
rect 22152 9404 22197 9432
rect 22152 9392 22158 9404
rect 22925 9367 22983 9373
rect 22925 9364 22937 9367
rect 21836 9336 22937 9364
rect 21361 9327 21419 9333
rect 22925 9333 22937 9336
rect 22971 9364 22983 9367
rect 23106 9364 23112 9376
rect 22971 9336 23112 9364
rect 22971 9333 22983 9336
rect 22925 9327 22983 9333
rect 23106 9324 23112 9336
rect 23164 9324 23170 9376
rect 23658 9364 23664 9376
rect 23619 9336 23664 9364
rect 23658 9324 23664 9336
rect 23716 9324 23722 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 7926 9160 7932 9172
rect 7887 9132 7932 9160
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 10781 9163 10839 9169
rect 10781 9160 10793 9163
rect 9272 9132 10793 9160
rect 9272 9120 9278 9132
rect 10781 9129 10793 9132
rect 10827 9129 10839 9163
rect 14458 9160 14464 9172
rect 14419 9132 14464 9160
rect 10781 9123 10839 9129
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 15470 9120 15476 9172
rect 15528 9160 15534 9172
rect 15565 9163 15623 9169
rect 15565 9160 15577 9163
rect 15528 9132 15577 9160
rect 15528 9120 15534 9132
rect 15565 9129 15577 9132
rect 15611 9129 15623 9163
rect 16942 9160 16948 9172
rect 16903 9132 16948 9160
rect 15565 9123 15623 9129
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 20162 9160 20168 9172
rect 20123 9132 20168 9160
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 21821 9163 21879 9169
rect 21821 9129 21833 9163
rect 21867 9160 21879 9163
rect 22094 9160 22100 9172
rect 21867 9132 22100 9160
rect 21867 9129 21879 9132
rect 21821 9123 21879 9129
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 23382 9120 23388 9172
rect 23440 9160 23446 9172
rect 23799 9163 23857 9169
rect 23799 9160 23811 9163
rect 23440 9132 23811 9160
rect 23440 9120 23446 9132
rect 23799 9129 23811 9132
rect 23845 9129 23857 9163
rect 23799 9123 23857 9129
rect 6362 9092 6368 9104
rect 6012 9064 6368 9092
rect 6012 9036 6040 9064
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 6546 9092 6552 9104
rect 6507 9064 6552 9092
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 8205 9095 8263 9101
rect 8205 9061 8217 9095
rect 8251 9092 8263 9095
rect 8294 9092 8300 9104
rect 8251 9064 8300 9092
rect 8251 9061 8263 9064
rect 8205 9055 8263 9061
rect 8294 9052 8300 9064
rect 8352 9052 8358 9104
rect 8754 9092 8760 9104
rect 8715 9064 8760 9092
rect 8754 9052 8760 9064
rect 8812 9052 8818 9104
rect 8938 9052 8944 9104
rect 8996 9092 9002 9104
rect 9125 9095 9183 9101
rect 9125 9092 9137 9095
rect 8996 9064 9137 9092
rect 8996 9052 9002 9064
rect 9125 9061 9137 9064
rect 9171 9092 9183 9095
rect 10870 9092 10876 9104
rect 9171 9064 10876 9092
rect 9171 9061 9183 9064
rect 9125 9055 9183 9061
rect 10870 9052 10876 9064
rect 10928 9092 10934 9104
rect 12434 9092 12440 9104
rect 10928 9064 12440 9092
rect 10928 9052 10934 9064
rect 106 8984 112 9036
rect 164 9024 170 9036
rect 1432 9027 1490 9033
rect 1432 9024 1444 9027
rect 164 8996 1444 9024
rect 164 8984 170 8996
rect 1432 8993 1444 8996
rect 1478 9024 1490 9027
rect 1578 9024 1584 9036
rect 1478 8996 1584 9024
rect 1478 8993 1490 8996
rect 1432 8987 1490 8993
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 5994 9024 6000 9036
rect 5955 8996 6000 9024
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 6273 9027 6331 9033
rect 6273 8993 6285 9027
rect 6319 9024 6331 9027
rect 6454 9024 6460 9036
rect 6319 8996 6460 9024
rect 6319 8993 6331 8996
rect 6273 8987 6331 8993
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 9024 9551 9027
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9539 8996 9689 9024
rect 9539 8993 9551 8996
rect 9493 8987 9551 8993
rect 9677 8993 9689 8996
rect 9723 9024 9735 9027
rect 10502 9024 10508 9036
rect 9723 8996 10508 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 11440 9033 11468 9064
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 12710 9052 12716 9104
rect 12768 9092 12774 9104
rect 13817 9095 13875 9101
rect 13817 9092 13829 9095
rect 12768 9064 13829 9092
rect 12768 9052 12774 9064
rect 13817 9061 13829 9064
rect 13863 9061 13875 9095
rect 13817 9055 13875 9061
rect 19613 9095 19671 9101
rect 19613 9061 19625 9095
rect 19659 9092 19671 9095
rect 20714 9092 20720 9104
rect 19659 9064 20720 9092
rect 19659 9061 19671 9064
rect 19613 9055 19671 9061
rect 20714 9052 20720 9064
rect 20772 9052 20778 9104
rect 20990 9052 20996 9104
rect 21048 9092 21054 9104
rect 21222 9095 21280 9101
rect 21222 9092 21234 9095
rect 21048 9064 21234 9092
rect 21048 9052 21054 9064
rect 21222 9061 21234 9064
rect 21268 9061 21280 9095
rect 21222 9055 21280 9061
rect 21358 9052 21364 9104
rect 21416 9092 21422 9104
rect 22787 9095 22845 9101
rect 22787 9092 22799 9095
rect 21416 9064 22799 9092
rect 21416 9052 21422 9064
rect 22787 9061 22799 9064
rect 22833 9061 22845 9095
rect 22787 9055 22845 9061
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 10652 8996 10701 9024
rect 10652 8984 10658 8996
rect 10689 8993 10701 8996
rect 10735 8993 10747 9027
rect 10689 8987 10747 8993
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 8993 11483 9027
rect 11425 8987 11483 8993
rect 11609 9027 11667 9033
rect 11609 8993 11621 9027
rect 11655 9024 11667 9027
rect 12069 9027 12127 9033
rect 11655 8996 11836 9024
rect 11655 8993 11667 8996
rect 11609 8987 11667 8993
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8925 8171 8959
rect 11698 8956 11704 8968
rect 8113 8919 8171 8925
rect 9876 8928 11704 8956
rect 1535 8891 1593 8897
rect 1535 8857 1547 8891
rect 1581 8888 1593 8891
rect 8018 8888 8024 8900
rect 1581 8860 8024 8888
rect 1581 8857 1593 8860
rect 1535 8851 1593 8857
rect 8018 8848 8024 8860
rect 8076 8888 8082 8900
rect 8128 8888 8156 8919
rect 8076 8860 8156 8888
rect 8076 8848 8082 8860
rect 6730 8780 6736 8832
rect 6788 8820 6794 8832
rect 9876 8829 9904 8928
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 11808 8888 11836 8996
rect 12069 8993 12081 9027
rect 12115 9024 12127 9027
rect 12802 9024 12808 9036
rect 12115 8996 12808 9024
rect 12115 8993 12127 8996
rect 12069 8987 12127 8993
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 12986 9024 12992 9036
rect 12947 8996 12992 9024
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 13170 9024 13176 9036
rect 13131 8996 13176 9024
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 15654 9024 15660 9036
rect 15615 8996 15660 9024
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 17218 8984 17224 9036
rect 17276 9024 17282 9036
rect 17313 9027 17371 9033
rect 17313 9024 17325 9027
rect 17276 8996 17325 9024
rect 17276 8984 17282 8996
rect 17313 8993 17325 8996
rect 17359 8993 17371 9027
rect 17770 9024 17776 9036
rect 17731 8996 17776 9024
rect 17313 8987 17371 8993
rect 17770 8984 17776 8996
rect 17828 8984 17834 9036
rect 19150 9024 19156 9036
rect 19111 8996 19156 9024
rect 19150 8984 19156 8996
rect 19208 8984 19214 9036
rect 19242 8984 19248 9036
rect 19300 9024 19306 9036
rect 19337 9027 19395 9033
rect 19337 9024 19349 9027
rect 19300 8996 19349 9024
rect 19300 8984 19306 8996
rect 19337 8993 19349 8996
rect 19383 8993 19395 9027
rect 19337 8987 19395 8993
rect 19978 8984 19984 9036
rect 20036 9024 20042 9036
rect 20901 9027 20959 9033
rect 20901 9024 20913 9027
rect 20036 8996 20913 9024
rect 20036 8984 20042 8996
rect 20901 8993 20913 8996
rect 20947 8993 20959 9027
rect 22646 9024 22652 9036
rect 22607 8996 22652 9024
rect 20901 8987 20959 8993
rect 22646 8984 22652 8996
rect 22704 8984 22710 9036
rect 23728 9027 23786 9033
rect 23728 8993 23740 9027
rect 23774 9024 23786 9027
rect 23842 9024 23848 9036
rect 23774 8996 23848 9024
rect 23774 8993 23786 8996
rect 23728 8987 23786 8993
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 18046 8956 18052 8968
rect 17959 8928 18052 8956
rect 18046 8916 18052 8928
rect 18104 8956 18110 8968
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 18104 8928 18337 8956
rect 18104 8916 18110 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 12250 8888 12256 8900
rect 11808 8860 12256 8888
rect 12250 8848 12256 8860
rect 12308 8888 12314 8900
rect 12805 8891 12863 8897
rect 12805 8888 12817 8891
rect 12308 8860 12817 8888
rect 12308 8848 12314 8860
rect 12805 8857 12817 8860
rect 12851 8888 12863 8891
rect 14274 8888 14280 8900
rect 12851 8860 14280 8888
rect 12851 8857 12863 8860
rect 12805 8851 12863 8857
rect 14274 8848 14280 8860
rect 14332 8848 14338 8900
rect 9861 8823 9919 8829
rect 9861 8820 9873 8823
rect 6788 8792 9873 8820
rect 6788 8780 6794 8792
rect 9861 8789 9873 8792
rect 9907 8789 9919 8823
rect 9861 8783 9919 8789
rect 10321 8823 10379 8829
rect 10321 8789 10333 8823
rect 10367 8820 10379 8823
rect 10686 8820 10692 8832
rect 10367 8792 10692 8820
rect 10367 8789 10379 8792
rect 10321 8783 10379 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 13262 8820 13268 8832
rect 13223 8792 13268 8820
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 14366 8780 14372 8832
rect 14424 8820 14430 8832
rect 14737 8823 14795 8829
rect 14737 8820 14749 8823
rect 14424 8792 14749 8820
rect 14424 8780 14430 8792
rect 14737 8789 14749 8792
rect 14783 8789 14795 8823
rect 14737 8783 14795 8789
rect 16206 8780 16212 8832
rect 16264 8820 16270 8832
rect 16301 8823 16359 8829
rect 16301 8820 16313 8823
rect 16264 8792 16313 8820
rect 16264 8780 16270 8792
rect 16301 8789 16313 8792
rect 16347 8789 16359 8823
rect 16301 8783 16359 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 1995 8619 2053 8625
rect 1995 8585 2007 8619
rect 2041 8616 2053 8619
rect 2222 8616 2228 8628
rect 2041 8588 2228 8616
rect 2041 8585 2053 8588
rect 1995 8579 2053 8585
rect 2222 8576 2228 8588
rect 2280 8576 2286 8628
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 3007 8619 3065 8625
rect 3007 8616 3019 8619
rect 2832 8588 3019 8616
rect 2832 8576 2838 8588
rect 3007 8585 3019 8588
rect 3053 8585 3065 8619
rect 3007 8579 3065 8585
rect 5905 8619 5963 8625
rect 5905 8585 5917 8619
rect 5951 8616 5963 8619
rect 5994 8616 6000 8628
rect 5951 8588 6000 8616
rect 5951 8585 5963 8588
rect 5905 8579 5963 8585
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6454 8616 6460 8628
rect 6319 8588 6460 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 6822 8576 6828 8628
rect 6880 8616 6886 8628
rect 6963 8619 7021 8625
rect 6963 8616 6975 8619
rect 6880 8588 6975 8616
rect 6880 8576 6886 8588
rect 6963 8585 6975 8588
rect 7009 8585 7021 8619
rect 6963 8579 7021 8585
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 8294 8616 8300 8628
rect 7883 8588 8300 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 8938 8616 8944 8628
rect 8899 8588 8944 8616
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9306 8616 9312 8628
rect 9267 8588 9312 8616
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10689 8619 10747 8625
rect 10689 8616 10701 8619
rect 10008 8588 10701 8616
rect 10008 8576 10014 8588
rect 10689 8585 10701 8588
rect 10735 8585 10747 8619
rect 11698 8616 11704 8628
rect 11611 8588 11704 8616
rect 10689 8579 10747 8585
rect 11698 8576 11704 8588
rect 11756 8616 11762 8628
rect 12250 8616 12256 8628
rect 11756 8588 12256 8616
rect 11756 8576 11762 8588
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 12710 8616 12716 8628
rect 12671 8588 12716 8616
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 12802 8576 12808 8628
rect 12860 8616 12866 8628
rect 14001 8619 14059 8625
rect 14001 8616 14013 8619
rect 12860 8588 14013 8616
rect 12860 8576 12866 8588
rect 14001 8585 14013 8588
rect 14047 8616 14059 8619
rect 14366 8616 14372 8628
rect 14047 8588 14372 8616
rect 14047 8585 14059 8588
rect 14001 8579 14059 8585
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 15838 8576 15844 8628
rect 15896 8616 15902 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 15896 8588 17325 8616
rect 15896 8576 15902 8588
rect 17313 8585 17325 8588
rect 17359 8616 17371 8619
rect 17770 8616 17776 8628
rect 17359 8588 17776 8616
rect 17359 8585 17371 8588
rect 17313 8579 17371 8585
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 19150 8576 19156 8628
rect 19208 8616 19214 8628
rect 19613 8619 19671 8625
rect 19613 8616 19625 8619
rect 19208 8588 19625 8616
rect 19208 8576 19214 8588
rect 19613 8585 19625 8588
rect 19659 8585 19671 8619
rect 19978 8616 19984 8628
rect 19939 8588 19984 8616
rect 19613 8579 19671 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 20717 8619 20775 8625
rect 20717 8585 20729 8619
rect 20763 8616 20775 8619
rect 20806 8616 20812 8628
rect 20763 8588 20812 8616
rect 20763 8585 20775 8588
rect 20717 8579 20775 8585
rect 10042 8508 10048 8560
rect 10100 8548 10106 8560
rect 10505 8551 10563 8557
rect 10505 8548 10517 8551
rect 10100 8520 10517 8548
rect 10100 8508 10106 8520
rect 10505 8517 10517 8520
rect 10551 8517 10563 8551
rect 14826 8548 14832 8560
rect 14739 8520 14832 8548
rect 10505 8511 10563 8517
rect 14826 8508 14832 8520
rect 14884 8548 14890 8560
rect 15378 8548 15384 8560
rect 14884 8520 15384 8548
rect 14884 8508 14890 8520
rect 15378 8508 15384 8520
rect 15436 8508 15442 8560
rect 17788 8548 17816 8576
rect 19242 8548 19248 8560
rect 17788 8520 19248 8548
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 6907 8452 7389 8480
rect 1394 8372 1400 8424
rect 1452 8412 1458 8424
rect 1892 8415 1950 8421
rect 1892 8412 1904 8415
rect 1452 8384 1904 8412
rect 1452 8372 1458 8384
rect 1892 8381 1904 8384
rect 1938 8412 1950 8415
rect 2314 8412 2320 8424
rect 1938 8384 2320 8412
rect 1938 8381 1950 8384
rect 1892 8375 1950 8381
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 2682 8372 2688 8424
rect 2740 8412 2746 8424
rect 6907 8421 6935 8452
rect 7377 8449 7389 8452
rect 7423 8480 7435 8483
rect 7834 8480 7840 8492
rect 7423 8452 7840 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 8619 8452 9045 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 9033 8449 9045 8452
rect 9079 8480 9091 8483
rect 9582 8480 9588 8492
rect 9079 8452 9588 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8480 10011 8483
rect 10594 8480 10600 8492
rect 9999 8452 10600 8480
rect 9999 8449 10011 8452
rect 9953 8443 10011 8449
rect 10594 8440 10600 8452
rect 10652 8480 10658 8492
rect 11241 8483 11299 8489
rect 11241 8480 11253 8483
rect 10652 8452 11253 8480
rect 10652 8440 10658 8452
rect 11241 8449 11253 8452
rect 11287 8480 11299 8483
rect 13170 8480 13176 8492
rect 11287 8452 13176 8480
rect 11287 8449 11299 8452
rect 11241 8443 11299 8449
rect 13170 8440 13176 8452
rect 13228 8480 13234 8492
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13228 8452 13645 8480
rect 13228 8440 13234 8452
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 16393 8483 16451 8489
rect 16393 8480 16405 8483
rect 16172 8452 16405 8480
rect 16172 8440 16178 8452
rect 16393 8449 16405 8452
rect 16439 8449 16451 8483
rect 16393 8443 16451 8449
rect 16850 8440 16856 8492
rect 16908 8480 16914 8492
rect 17773 8483 17831 8489
rect 17773 8480 17785 8483
rect 16908 8452 17785 8480
rect 16908 8440 16914 8452
rect 17773 8449 17785 8452
rect 17819 8449 17831 8483
rect 18046 8480 18052 8492
rect 18007 8452 18052 8480
rect 17773 8443 17831 8449
rect 2904 8415 2962 8421
rect 2904 8412 2916 8415
rect 2740 8384 2916 8412
rect 2740 8372 2746 8384
rect 2904 8381 2916 8384
rect 2950 8412 2962 8415
rect 3329 8415 3387 8421
rect 3329 8412 3341 8415
rect 2950 8384 3341 8412
rect 2950 8381 2962 8384
rect 2904 8375 2962 8381
rect 3329 8381 3341 8384
rect 3375 8381 3387 8415
rect 3329 8375 3387 8381
rect 6892 8415 6950 8421
rect 6892 8381 6904 8415
rect 6938 8381 6950 8415
rect 6892 8375 6950 8381
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8812 8415 8870 8421
rect 8812 8412 8824 8415
rect 8251 8384 8824 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8812 8381 8824 8384
rect 8858 8412 8870 8415
rect 10376 8415 10434 8421
rect 10376 8412 10388 8415
rect 8858 8384 10388 8412
rect 8858 8381 8870 8384
rect 8812 8375 8870 8381
rect 10376 8381 10388 8384
rect 10422 8412 10434 8415
rect 10686 8412 10692 8424
rect 10422 8384 10692 8412
rect 10422 8381 10434 8384
rect 10376 8375 10434 8381
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 10796 8384 12572 8412
rect 8665 8347 8723 8353
rect 8665 8313 8677 8347
rect 8711 8344 8723 8347
rect 9030 8344 9036 8356
rect 8711 8316 9036 8344
rect 8711 8313 8723 8316
rect 8665 8307 8723 8313
rect 9030 8304 9036 8316
rect 9088 8344 9094 8356
rect 10229 8347 10287 8353
rect 10229 8344 10241 8347
rect 9088 8316 10241 8344
rect 9088 8304 9094 8316
rect 10229 8313 10241 8316
rect 10275 8313 10287 8347
rect 10229 8307 10287 8313
rect 10502 8304 10508 8356
rect 10560 8344 10566 8356
rect 10796 8344 10824 8384
rect 12434 8344 12440 8356
rect 10560 8316 10824 8344
rect 12395 8316 12440 8344
rect 10560 8304 10566 8316
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 12544 8344 12572 8384
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 12676 8384 12721 8412
rect 12676 8372 12682 8384
rect 14366 8372 14372 8424
rect 14424 8412 14430 8424
rect 14737 8415 14795 8421
rect 14737 8412 14749 8415
rect 14424 8384 14749 8412
rect 14424 8372 14430 8384
rect 14737 8381 14749 8384
rect 14783 8412 14795 8415
rect 14918 8412 14924 8424
rect 14783 8384 14924 8412
rect 14783 8381 14795 8384
rect 14737 8375 14795 8381
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 15013 8415 15071 8421
rect 15013 8381 15025 8415
rect 15059 8412 15071 8415
rect 15654 8412 15660 8424
rect 15059 8384 15660 8412
rect 15059 8381 15071 8384
rect 15013 8375 15071 8381
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 16206 8372 16212 8424
rect 16264 8412 16270 8424
rect 16301 8415 16359 8421
rect 16301 8412 16313 8415
rect 16264 8384 16313 8412
rect 16264 8372 16270 8384
rect 16301 8381 16313 8384
rect 16347 8381 16359 8415
rect 16301 8375 16359 8381
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 16577 8415 16635 8421
rect 16577 8412 16589 8415
rect 16540 8384 16589 8412
rect 16540 8372 16546 8384
rect 16577 8381 16589 8384
rect 16623 8381 16635 8415
rect 16577 8375 16635 8381
rect 17788 8344 17816 8443
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 20232 8415 20290 8421
rect 20232 8412 20244 8415
rect 19392 8384 20244 8412
rect 19392 8372 19398 8384
rect 20232 8381 20244 8384
rect 20278 8412 20290 8415
rect 20732 8412 20760 8579
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 20990 8616 20996 8628
rect 20951 8588 20996 8616
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 21818 8576 21824 8628
rect 21876 8616 21882 8628
rect 22189 8619 22247 8625
rect 22189 8616 22201 8619
rect 21876 8588 22201 8616
rect 21876 8576 21882 8588
rect 22189 8585 22201 8588
rect 22235 8585 22247 8619
rect 23842 8616 23848 8628
rect 23803 8588 23848 8616
rect 22189 8579 22247 8585
rect 23842 8576 23848 8588
rect 23900 8576 23906 8628
rect 21910 8480 21916 8492
rect 21871 8452 21916 8480
rect 21910 8440 21916 8452
rect 21968 8440 21974 8492
rect 20278 8384 20760 8412
rect 20278 8381 20290 8384
rect 20232 8375 20290 8381
rect 18370 8347 18428 8353
rect 18370 8344 18382 8347
rect 12544 8316 16436 8344
rect 17788 8316 18382 8344
rect 9674 8276 9680 8288
rect 9635 8248 9680 8276
rect 9674 8236 9680 8248
rect 9732 8276 9738 8288
rect 9953 8279 10011 8285
rect 9953 8276 9965 8279
rect 9732 8248 9965 8276
rect 9732 8236 9738 8248
rect 9953 8245 9965 8248
rect 9999 8245 10011 8279
rect 9953 8239 10011 8245
rect 10042 8236 10048 8288
rect 10100 8276 10106 8288
rect 12158 8276 12164 8288
rect 10100 8248 10145 8276
rect 12119 8248 12164 8276
rect 10100 8236 10106 8248
rect 12158 8236 12164 8248
rect 12216 8276 12222 8288
rect 12618 8276 12624 8288
rect 12216 8248 12624 8276
rect 12216 8236 12222 8248
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 13357 8279 13415 8285
rect 13357 8276 13369 8279
rect 13044 8248 13369 8276
rect 13044 8236 13050 8248
rect 13357 8245 13369 8248
rect 13403 8276 13415 8279
rect 13630 8276 13636 8288
rect 13403 8248 13636 8276
rect 13403 8245 13415 8248
rect 13357 8239 13415 8245
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 14550 8276 14556 8288
rect 14511 8248 14556 8276
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 15197 8279 15255 8285
rect 15197 8245 15209 8279
rect 15243 8276 15255 8279
rect 15286 8276 15292 8288
rect 15243 8248 15292 8276
rect 15243 8245 15255 8248
rect 15197 8239 15255 8245
rect 15286 8236 15292 8248
rect 15344 8236 15350 8288
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 15749 8279 15807 8285
rect 15749 8276 15761 8279
rect 15712 8248 15761 8276
rect 15712 8236 15718 8248
rect 15749 8245 15761 8248
rect 15795 8276 15807 8279
rect 16117 8279 16175 8285
rect 16117 8276 16129 8279
rect 15795 8248 16129 8276
rect 15795 8245 15807 8248
rect 15749 8239 15807 8245
rect 16117 8245 16129 8248
rect 16163 8276 16175 8279
rect 16298 8276 16304 8288
rect 16163 8248 16304 8276
rect 16163 8245 16175 8248
rect 16117 8239 16175 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 16408 8276 16436 8316
rect 18370 8313 18382 8316
rect 18416 8313 18428 8347
rect 21269 8347 21327 8353
rect 21269 8344 21281 8347
rect 18370 8307 18428 8313
rect 20548 8316 21281 8344
rect 20548 8288 20576 8316
rect 21269 8313 21281 8316
rect 21315 8313 21327 8347
rect 21269 8307 21327 8313
rect 21361 8347 21419 8353
rect 21361 8313 21373 8347
rect 21407 8344 21419 8347
rect 21726 8344 21732 8356
rect 21407 8316 21732 8344
rect 21407 8313 21419 8316
rect 21361 8307 21419 8313
rect 21726 8304 21732 8316
rect 21784 8304 21790 8356
rect 16761 8279 16819 8285
rect 16761 8276 16773 8279
rect 16408 8248 16773 8276
rect 16761 8245 16773 8248
rect 16807 8245 16819 8279
rect 18966 8276 18972 8288
rect 18927 8248 18972 8276
rect 16761 8239 16819 8245
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 20303 8279 20361 8285
rect 20303 8245 20315 8279
rect 20349 8276 20361 8279
rect 20530 8276 20536 8288
rect 20349 8248 20536 8276
rect 20349 8245 20361 8248
rect 20303 8239 20361 8245
rect 20530 8236 20536 8248
rect 20588 8236 20594 8288
rect 22646 8276 22652 8288
rect 22607 8248 22652 8276
rect 22646 8236 22652 8248
rect 22704 8276 22710 8288
rect 27706 8276 27712 8288
rect 22704 8248 27712 8276
rect 22704 8236 22710 8248
rect 27706 8236 27712 8248
rect 27764 8236 27770 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1535 8075 1593 8081
rect 1535 8041 1547 8075
rect 1581 8072 1593 8075
rect 8938 8072 8944 8084
rect 1581 8044 8944 8072
rect 1581 8041 1593 8044
rect 1535 8035 1593 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 9030 8032 9036 8084
rect 9088 8072 9094 8084
rect 9398 8072 9404 8084
rect 9088 8044 9404 8072
rect 9088 8032 9094 8044
rect 9398 8032 9404 8044
rect 9456 8072 9462 8084
rect 9456 8044 9812 8072
rect 9456 8032 9462 8044
rect 2547 8007 2605 8013
rect 2547 7973 2559 8007
rect 2593 8004 2605 8007
rect 4154 8004 4160 8016
rect 2593 7976 4160 8004
rect 2593 7973 2605 7976
rect 2547 7967 2605 7973
rect 4154 7964 4160 7976
rect 4212 7964 4218 8016
rect 8018 8004 8024 8016
rect 7979 7976 8024 8004
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 9784 8013 9812 8044
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 11793 8075 11851 8081
rect 11793 8072 11805 8075
rect 9916 8044 11805 8072
rect 9916 8032 9922 8044
rect 11793 8041 11805 8044
rect 11839 8041 11851 8075
rect 12434 8072 12440 8084
rect 12347 8044 12440 8072
rect 11793 8035 11851 8041
rect 12434 8032 12440 8044
rect 12492 8072 12498 8084
rect 12713 8075 12771 8081
rect 12713 8072 12725 8075
rect 12492 8044 12725 8072
rect 12492 8032 12498 8044
rect 12713 8041 12725 8044
rect 12759 8041 12771 8075
rect 12713 8035 12771 8041
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 13081 8075 13139 8081
rect 13081 8072 13093 8075
rect 12952 8044 13093 8072
rect 12952 8032 12958 8044
rect 13081 8041 13093 8044
rect 13127 8041 13139 8075
rect 14826 8072 14832 8084
rect 14787 8044 14832 8072
rect 13081 8035 13139 8041
rect 14826 8032 14832 8044
rect 14884 8032 14890 8084
rect 17037 8075 17095 8081
rect 17037 8041 17049 8075
rect 17083 8072 17095 8075
rect 17494 8072 17500 8084
rect 17083 8044 17500 8072
rect 17083 8041 17095 8044
rect 17037 8035 17095 8041
rect 17494 8032 17500 8044
rect 17552 8072 17558 8084
rect 19150 8072 19156 8084
rect 17552 8044 19156 8072
rect 17552 8032 17558 8044
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 19751 8075 19809 8081
rect 19751 8072 19763 8075
rect 19576 8044 19763 8072
rect 19576 8032 19582 8044
rect 19751 8041 19763 8044
rect 19797 8041 19809 8075
rect 19751 8035 19809 8041
rect 20530 8032 20536 8084
rect 20588 8072 20594 8084
rect 20625 8075 20683 8081
rect 20625 8072 20637 8075
rect 20588 8044 20637 8072
rect 20588 8032 20594 8044
rect 20625 8041 20637 8044
rect 20671 8041 20683 8075
rect 20625 8035 20683 8041
rect 9769 8007 9827 8013
rect 9769 7973 9781 8007
rect 9815 8004 9827 8007
rect 10781 8007 10839 8013
rect 10781 8004 10793 8007
rect 9815 7976 10793 8004
rect 9815 7973 9827 7976
rect 9769 7967 9827 7973
rect 10781 7973 10793 7976
rect 10827 7973 10839 8007
rect 10781 7967 10839 7973
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 18233 8007 18291 8013
rect 18233 8004 18245 8007
rect 17920 7976 18245 8004
rect 17920 7964 17926 7976
rect 18233 7973 18245 7976
rect 18279 8004 18291 8007
rect 18966 8004 18972 8016
rect 18279 7976 18972 8004
rect 18279 7973 18291 7976
rect 18233 7967 18291 7973
rect 18966 7964 18972 7976
rect 19024 7964 19030 8016
rect 20990 7964 20996 8016
rect 21048 8004 21054 8016
rect 21222 8007 21280 8013
rect 21222 8004 21234 8007
rect 21048 7976 21234 8004
rect 21048 7964 21054 7976
rect 21222 7973 21234 7976
rect 21268 7973 21280 8007
rect 21222 7967 21280 7973
rect 1464 7939 1522 7945
rect 1464 7905 1476 7939
rect 1510 7905 1522 7939
rect 2406 7936 2412 7948
rect 2367 7908 2412 7936
rect 1464 7899 1522 7905
rect 106 7760 112 7812
rect 164 7800 170 7812
rect 1479 7800 1507 7899
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 9916 7939 9974 7945
rect 8619 7908 8800 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 1854 7800 1860 7812
rect 164 7772 1860 7800
rect 164 7760 170 7772
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 8662 7760 8668 7812
rect 8720 7800 8726 7812
rect 8772 7800 8800 7908
rect 9916 7905 9928 7939
rect 9962 7936 9974 7939
rect 10686 7936 10692 7948
rect 9962 7908 10692 7936
rect 9962 7905 9974 7908
rect 9916 7899 9974 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 11296 7908 11345 7936
rect 11296 7896 11302 7908
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 11609 7939 11667 7945
rect 11609 7905 11621 7939
rect 11655 7936 11667 7939
rect 12158 7936 12164 7948
rect 11655 7908 12164 7936
rect 11655 7905 11667 7908
rect 11609 7899 11667 7905
rect 9582 7828 9588 7880
rect 9640 7868 9646 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 9640 7840 10149 7868
rect 9640 7828 9646 7840
rect 10137 7837 10149 7840
rect 10183 7868 10195 7871
rect 11624 7868 11652 7899
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 14277 7939 14335 7945
rect 14277 7905 14289 7939
rect 14323 7936 14335 7939
rect 14826 7936 14832 7948
rect 14323 7908 14832 7936
rect 14323 7905 14335 7908
rect 14277 7899 14335 7905
rect 14826 7896 14832 7908
rect 14884 7896 14890 7948
rect 14918 7896 14924 7948
rect 14976 7936 14982 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 14976 7908 15301 7936
rect 14976 7896 14982 7908
rect 15289 7905 15301 7908
rect 15335 7936 15347 7939
rect 15470 7936 15476 7948
rect 15335 7908 15476 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 15470 7896 15476 7908
rect 15528 7896 15534 7948
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7936 15623 7939
rect 15654 7936 15660 7948
rect 15611 7908 15660 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 16022 7896 16028 7948
rect 16080 7936 16086 7948
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 16080 7908 16865 7936
rect 16080 7896 16086 7908
rect 16853 7905 16865 7908
rect 16899 7936 16911 7939
rect 17310 7936 17316 7948
rect 16899 7908 17316 7936
rect 16899 7905 16911 7908
rect 16853 7899 16911 7905
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 18782 7896 18788 7948
rect 18840 7936 18846 7948
rect 19680 7939 19738 7945
rect 19680 7936 19692 7939
rect 18840 7908 19692 7936
rect 18840 7896 18846 7908
rect 19680 7905 19692 7908
rect 19726 7936 19738 7939
rect 20073 7939 20131 7945
rect 20073 7936 20085 7939
rect 19726 7908 20085 7936
rect 19726 7905 19738 7908
rect 19680 7899 19738 7905
rect 20073 7905 20085 7908
rect 20119 7905 20131 7939
rect 20073 7899 20131 7905
rect 10183 7840 11652 7868
rect 14369 7871 14427 7877
rect 10183 7837 10195 7840
rect 10137 7831 10195 7837
rect 14369 7837 14381 7871
rect 14415 7868 14427 7871
rect 15381 7871 15439 7877
rect 15381 7868 15393 7871
rect 14415 7840 15393 7868
rect 14415 7837 14427 7840
rect 14369 7831 14427 7837
rect 15381 7837 15393 7840
rect 15427 7837 15439 7871
rect 15746 7868 15752 7880
rect 15707 7840 15752 7868
rect 15381 7831 15439 7837
rect 10229 7803 10287 7809
rect 10229 7800 10241 7803
rect 8720 7772 10241 7800
rect 8720 7760 8726 7772
rect 10229 7769 10241 7772
rect 10275 7769 10287 7803
rect 10229 7763 10287 7769
rect 11425 7803 11483 7809
rect 11425 7769 11437 7803
rect 11471 7800 11483 7803
rect 11514 7800 11520 7812
rect 11471 7772 11520 7800
rect 11471 7769 11483 7772
rect 11425 7763 11483 7769
rect 11514 7760 11520 7772
rect 11572 7760 11578 7812
rect 15396 7800 15424 7831
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18598 7868 18604 7880
rect 18559 7840 18604 7868
rect 18141 7831 18199 7837
rect 16114 7800 16120 7812
rect 15396 7772 16120 7800
rect 16114 7760 16120 7772
rect 16172 7800 16178 7812
rect 16301 7803 16359 7809
rect 16301 7800 16313 7803
rect 16172 7772 16313 7800
rect 16172 7760 16178 7772
rect 16301 7769 16313 7772
rect 16347 7769 16359 7803
rect 16301 7763 16359 7769
rect 8570 7692 8576 7744
rect 8628 7732 8634 7744
rect 8757 7735 8815 7741
rect 8757 7732 8769 7735
rect 8628 7704 8769 7732
rect 8628 7692 8634 7704
rect 8757 7701 8769 7704
rect 8803 7701 8815 7735
rect 9490 7732 9496 7744
rect 9451 7704 9496 7732
rect 8757 7695 8815 7701
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 10042 7732 10048 7744
rect 10003 7704 10048 7732
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 11238 7732 11244 7744
rect 11199 7704 11244 7732
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 16666 7732 16672 7744
rect 16627 7704 16672 7732
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 17218 7692 17224 7744
rect 17276 7732 17282 7744
rect 17313 7735 17371 7741
rect 17313 7732 17325 7735
rect 17276 7704 17325 7732
rect 17276 7692 17282 7704
rect 17313 7701 17325 7704
rect 17359 7701 17371 7735
rect 17313 7695 17371 7701
rect 17402 7692 17408 7744
rect 17460 7732 17466 7744
rect 17865 7735 17923 7741
rect 17865 7732 17877 7735
rect 17460 7704 17877 7732
rect 17460 7692 17466 7704
rect 17865 7701 17877 7704
rect 17911 7732 17923 7735
rect 18156 7732 18184 7831
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 20346 7828 20352 7880
rect 20404 7868 20410 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20404 7840 20913 7868
rect 20404 7828 20410 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 17911 7704 18184 7732
rect 17911 7701 17923 7704
rect 17865 7695 17923 7701
rect 18230 7692 18236 7744
rect 18288 7732 18294 7744
rect 19061 7735 19119 7741
rect 19061 7732 19073 7735
rect 18288 7704 19073 7732
rect 18288 7692 18294 7704
rect 19061 7701 19073 7704
rect 19107 7701 19119 7735
rect 21818 7732 21824 7744
rect 21779 7704 21824 7732
rect 19061 7695 19119 7701
rect 21818 7692 21824 7704
rect 21876 7692 21882 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1535 7531 1593 7537
rect 1535 7497 1547 7531
rect 1581 7528 1593 7531
rect 1670 7528 1676 7540
rect 1581 7500 1676 7528
rect 1581 7497 1593 7500
rect 1535 7491 1593 7497
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 1854 7528 1860 7540
rect 1815 7500 1860 7528
rect 1854 7488 1860 7500
rect 1912 7488 1918 7540
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 9401 7531 9459 7537
rect 9401 7497 9413 7531
rect 9447 7528 9459 7531
rect 9582 7528 9588 7540
rect 9447 7500 9588 7528
rect 9447 7497 9459 7500
rect 9401 7491 9459 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 9677 7531 9735 7537
rect 9677 7497 9689 7531
rect 9723 7528 9735 7531
rect 11698 7528 11704 7540
rect 9723 7500 11704 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 16114 7528 16120 7540
rect 16075 7500 16120 7528
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 17310 7488 17316 7540
rect 17368 7528 17374 7540
rect 17405 7531 17463 7537
rect 17405 7528 17417 7531
rect 17368 7500 17417 7528
rect 17368 7488 17374 7500
rect 17405 7497 17417 7500
rect 17451 7497 17463 7531
rect 17862 7528 17868 7540
rect 17823 7500 17868 7528
rect 17405 7491 17463 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 19058 7528 19064 7540
rect 19019 7500 19064 7528
rect 19058 7488 19064 7500
rect 19116 7488 19122 7540
rect 19242 7488 19248 7540
rect 19300 7528 19306 7540
rect 19429 7531 19487 7537
rect 19429 7528 19441 7531
rect 19300 7500 19441 7528
rect 19300 7488 19306 7500
rect 19429 7497 19441 7500
rect 19475 7497 19487 7531
rect 20990 7528 20996 7540
rect 20951 7500 20996 7528
rect 19429 7491 19487 7497
rect 9490 7420 9496 7472
rect 9548 7460 9554 7472
rect 9548 7432 9674 7460
rect 9548 7420 9554 7432
rect 1210 7352 1216 7404
rect 1268 7392 1274 7404
rect 9646 7392 9674 7432
rect 11054 7420 11060 7472
rect 11112 7460 11118 7472
rect 14185 7463 14243 7469
rect 14185 7460 14197 7463
rect 11112 7432 14197 7460
rect 11112 7420 11118 7432
rect 14185 7429 14197 7432
rect 14231 7460 14243 7463
rect 14826 7460 14832 7472
rect 14231 7432 14832 7460
rect 14231 7429 14243 7432
rect 14185 7423 14243 7429
rect 14826 7420 14832 7432
rect 14884 7420 14890 7472
rect 11238 7392 11244 7404
rect 1268 7364 1507 7392
rect 1268 7352 1274 7364
rect 1479 7333 1507 7364
rect 9646 7364 11244 7392
rect 1464 7327 1522 7333
rect 1464 7293 1476 7327
rect 1510 7293 1522 7327
rect 1464 7287 1522 7293
rect 9519 7327 9577 7333
rect 9519 7293 9531 7327
rect 9565 7324 9577 7327
rect 9646 7324 9674 7364
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 11514 7352 11520 7404
rect 11572 7392 11578 7404
rect 11609 7395 11667 7401
rect 11609 7392 11621 7395
rect 11572 7364 11621 7392
rect 11572 7352 11578 7364
rect 11609 7361 11621 7364
rect 11655 7392 11667 7395
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 11655 7364 13001 7392
rect 11655 7361 11667 7364
rect 11609 7355 11667 7361
rect 12989 7361 13001 7364
rect 13035 7392 13047 7395
rect 13173 7395 13231 7401
rect 13173 7392 13185 7395
rect 13035 7364 13185 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13173 7361 13185 7364
rect 13219 7392 13231 7395
rect 13630 7392 13636 7404
rect 13219 7364 13636 7392
rect 13219 7361 13231 7364
rect 13173 7355 13231 7361
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17494 7392 17500 7404
rect 17175 7364 17500 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17494 7352 17500 7364
rect 17552 7392 17558 7404
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 17552 7364 18153 7392
rect 17552 7352 17558 7364
rect 18141 7361 18153 7364
rect 18187 7392 18199 7395
rect 18230 7392 18236 7404
rect 18187 7364 18236 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 18230 7352 18236 7364
rect 18288 7352 18294 7404
rect 18782 7392 18788 7404
rect 18743 7364 18788 7392
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 19444 7392 19472 7491
rect 20990 7488 20996 7500
rect 21048 7528 21054 7540
rect 25958 7528 25964 7540
rect 21048 7500 25964 7528
rect 21048 7488 21054 7500
rect 25958 7488 25964 7500
rect 26016 7488 26022 7540
rect 21910 7392 21916 7404
rect 19444 7364 20116 7392
rect 21871 7364 21916 7392
rect 10042 7324 10048 7336
rect 9565 7296 9674 7324
rect 9955 7296 10048 7324
rect 9565 7293 9577 7296
rect 9519 7287 9577 7293
rect 10042 7284 10048 7296
rect 10100 7324 10106 7336
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 10100 7296 10425 7324
rect 10100 7284 10106 7296
rect 10413 7293 10425 7296
rect 10459 7324 10471 7327
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 10459 7296 11161 7324
rect 10459 7293 10471 7296
rect 10413 7287 10471 7293
rect 11149 7293 11161 7296
rect 11195 7324 11207 7327
rect 11532 7324 11560 7352
rect 11195 7296 11560 7324
rect 11195 7293 11207 7296
rect 11149 7287 11207 7293
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 13081 7327 13139 7333
rect 13081 7324 13093 7327
rect 12952 7296 13093 7324
rect 12952 7284 12958 7296
rect 13081 7293 13093 7296
rect 13127 7293 13139 7327
rect 13081 7287 13139 7293
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7293 13415 7327
rect 14734 7324 14740 7336
rect 14695 7296 14740 7324
rect 13357 7287 13415 7293
rect 9033 7259 9091 7265
rect 9033 7225 9045 7259
rect 9079 7256 9091 7259
rect 10686 7256 10692 7268
rect 9079 7228 10692 7256
rect 9079 7225 9091 7228
rect 9033 7219 9091 7225
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 11241 7259 11299 7265
rect 11241 7225 11253 7259
rect 11287 7256 11299 7259
rect 12434 7256 12440 7268
rect 11287 7228 12440 7256
rect 11287 7225 11299 7228
rect 11241 7219 11299 7225
rect 12434 7216 12440 7228
rect 12492 7216 12498 7268
rect 13170 7216 13176 7268
rect 13228 7256 13234 7268
rect 13372 7256 13400 7287
rect 14734 7284 14740 7296
rect 14792 7284 14798 7336
rect 15013 7327 15071 7333
rect 15013 7293 15025 7327
rect 15059 7324 15071 7327
rect 15654 7324 15660 7336
rect 15059 7296 15660 7324
rect 15059 7293 15071 7296
rect 15013 7287 15071 7293
rect 13228 7228 13400 7256
rect 13228 7216 13234 7228
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 13872 7228 13917 7256
rect 13872 7216 13878 7228
rect 2406 7148 2412 7200
rect 2464 7188 2470 7200
rect 2501 7191 2559 7197
rect 2501 7188 2513 7191
rect 2464 7160 2513 7188
rect 2464 7148 2470 7160
rect 2501 7157 2513 7160
rect 2547 7188 2559 7191
rect 5534 7188 5540 7200
rect 2547 7160 5540 7188
rect 2547 7157 2559 7160
rect 2501 7151 2559 7157
rect 5534 7148 5540 7160
rect 5592 7188 5598 7200
rect 7558 7188 7564 7200
rect 5592 7160 7564 7188
rect 5592 7148 5598 7160
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 10042 7148 10048 7200
rect 10100 7188 10106 7200
rect 11882 7188 11888 7200
rect 10100 7160 11888 7188
rect 10100 7148 10106 7160
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 11977 7191 12035 7197
rect 11977 7157 11989 7191
rect 12023 7188 12035 7191
rect 12158 7188 12164 7200
rect 12023 7160 12164 7188
rect 12023 7157 12035 7160
rect 11977 7151 12035 7157
rect 12158 7148 12164 7160
rect 12216 7188 12222 7200
rect 13188 7188 13216 7216
rect 14550 7188 14556 7200
rect 12216 7160 13216 7188
rect 14511 7160 14556 7188
rect 12216 7148 12222 7160
rect 14550 7148 14556 7160
rect 14608 7188 14614 7200
rect 15028 7188 15056 7287
rect 15654 7284 15660 7296
rect 15712 7324 15718 7336
rect 15749 7327 15807 7333
rect 15749 7324 15761 7327
rect 15712 7296 15761 7324
rect 15712 7284 15718 7296
rect 15749 7293 15761 7296
rect 15795 7293 15807 7327
rect 15749 7287 15807 7293
rect 19058 7284 19064 7336
rect 19116 7324 19122 7336
rect 20088 7333 20116 7364
rect 21910 7352 21916 7364
rect 21968 7352 21974 7404
rect 19613 7327 19671 7333
rect 19613 7324 19625 7327
rect 19116 7296 19625 7324
rect 19116 7284 19122 7296
rect 19613 7293 19625 7296
rect 19659 7293 19671 7327
rect 19613 7287 19671 7293
rect 20073 7327 20131 7333
rect 20073 7293 20085 7327
rect 20119 7293 20131 7327
rect 20073 7287 20131 7293
rect 15470 7256 15476 7268
rect 15431 7228 15476 7256
rect 15470 7216 15476 7228
rect 15528 7216 15534 7268
rect 16482 7256 16488 7268
rect 16443 7228 16488 7256
rect 16482 7216 16488 7228
rect 16540 7216 16546 7268
rect 16577 7259 16635 7265
rect 16577 7225 16589 7259
rect 16623 7256 16635 7259
rect 16666 7256 16672 7268
rect 16623 7228 16672 7256
rect 16623 7225 16635 7228
rect 16577 7219 16635 7225
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 18230 7216 18236 7268
rect 18288 7256 18294 7268
rect 18288 7228 18333 7256
rect 18288 7216 18294 7228
rect 14608 7160 15056 7188
rect 14608 7148 14614 7160
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 19076 7188 19104 7284
rect 20346 7256 20352 7268
rect 20307 7228 20352 7256
rect 20346 7216 20352 7228
rect 20404 7216 20410 7268
rect 21453 7259 21511 7265
rect 21453 7225 21465 7259
rect 21499 7225 21511 7259
rect 21453 7219 21511 7225
rect 21545 7259 21603 7265
rect 21545 7225 21557 7259
rect 21591 7256 21603 7259
rect 21818 7256 21824 7268
rect 21591 7228 21824 7256
rect 21591 7225 21603 7228
rect 21545 7219 21603 7225
rect 15436 7160 19104 7188
rect 21468 7188 21496 7219
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 22370 7188 22376 7200
rect 21468 7160 22376 7188
rect 15436 7148 15442 7160
rect 22370 7148 22376 7160
rect 22428 7148 22434 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1210 6944 1216 6996
rect 1268 6984 1274 6996
rect 1581 6987 1639 6993
rect 1581 6984 1593 6987
rect 1268 6956 1593 6984
rect 1268 6944 1274 6956
rect 1581 6953 1593 6956
rect 1627 6953 1639 6987
rect 9398 6984 9404 6996
rect 9359 6956 9404 6984
rect 1581 6947 1639 6953
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 14826 6984 14832 6996
rect 14787 6956 14832 6984
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 15378 6944 15384 6996
rect 15436 6984 15442 6996
rect 15473 6987 15531 6993
rect 15473 6984 15485 6987
rect 15436 6956 15485 6984
rect 15436 6944 15442 6956
rect 15473 6953 15485 6956
rect 15519 6953 15531 6987
rect 15473 6947 15531 6953
rect 15562 6944 15568 6996
rect 15620 6984 15626 6996
rect 16117 6987 16175 6993
rect 16117 6984 16129 6987
rect 15620 6956 16129 6984
rect 15620 6944 15626 6956
rect 16117 6953 16129 6956
rect 16163 6953 16175 6987
rect 16117 6947 16175 6953
rect 16482 6944 16488 6996
rect 16540 6984 16546 6996
rect 17681 6987 17739 6993
rect 17681 6984 17693 6987
rect 16540 6956 17693 6984
rect 16540 6944 16546 6956
rect 17681 6953 17693 6956
rect 17727 6984 17739 6987
rect 19843 6987 19901 6993
rect 19843 6984 19855 6987
rect 17727 6956 19855 6984
rect 17727 6953 17739 6956
rect 17681 6947 17739 6953
rect 19843 6953 19855 6956
rect 19889 6953 19901 6987
rect 19843 6947 19901 6953
rect 21453 6987 21511 6993
rect 21453 6953 21465 6987
rect 21499 6984 21511 6987
rect 21818 6984 21824 6996
rect 21499 6956 21824 6984
rect 21499 6953 21511 6956
rect 21453 6947 21511 6953
rect 21818 6944 21824 6956
rect 21876 6944 21882 6996
rect 9674 6916 9680 6928
rect 9635 6888 9680 6916
rect 9674 6876 9680 6888
rect 9732 6876 9738 6928
rect 14734 6916 14740 6928
rect 14108 6888 14740 6916
rect 10318 6848 10324 6860
rect 10279 6820 10324 6848
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 11330 6848 11336 6860
rect 11291 6820 11336 6848
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 13262 6848 13268 6860
rect 13223 6820 13268 6848
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 14108 6857 14136 6888
rect 14734 6876 14740 6888
rect 14792 6916 14798 6928
rect 15749 6919 15807 6925
rect 15749 6916 15761 6919
rect 14792 6888 15761 6916
rect 14792 6876 14798 6888
rect 15749 6885 15761 6888
rect 15795 6916 15807 6919
rect 16206 6916 16212 6928
rect 15795 6888 16212 6916
rect 15795 6885 15807 6888
rect 15749 6879 15807 6885
rect 16206 6876 16212 6888
rect 16264 6876 16270 6928
rect 16755 6919 16813 6925
rect 16755 6885 16767 6919
rect 16801 6916 16813 6919
rect 16850 6916 16856 6928
rect 16801 6888 16856 6916
rect 16801 6885 16813 6888
rect 16755 6879 16813 6885
rect 16850 6876 16856 6888
rect 16908 6876 16914 6928
rect 18322 6916 18328 6928
rect 18283 6888 18328 6916
rect 18322 6876 18328 6888
rect 18380 6876 18386 6928
rect 20346 6876 20352 6928
rect 20404 6916 20410 6928
rect 21729 6919 21787 6925
rect 21729 6916 21741 6919
rect 20404 6888 21741 6916
rect 20404 6876 20410 6888
rect 21729 6885 21741 6888
rect 21775 6885 21787 6919
rect 21729 6879 21787 6885
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13786 6820 14105 6848
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12986 6780 12992 6792
rect 12023 6752 12992 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12986 6740 12992 6752
rect 13044 6780 13050 6792
rect 13786 6780 13814 6820
rect 14093 6817 14105 6820
rect 14139 6817 14151 6851
rect 14274 6848 14280 6860
rect 14235 6820 14280 6848
rect 14093 6811 14151 6817
rect 14274 6808 14280 6820
rect 14332 6808 14338 6860
rect 15289 6851 15347 6857
rect 15289 6817 15301 6851
rect 15335 6848 15347 6851
rect 15470 6848 15476 6860
rect 15335 6820 15476 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 19518 6808 19524 6860
rect 19576 6848 19582 6860
rect 19740 6851 19798 6857
rect 19740 6848 19752 6851
rect 19576 6820 19752 6848
rect 19576 6808 19582 6820
rect 19740 6817 19752 6820
rect 19786 6817 19798 6851
rect 19740 6811 19798 6817
rect 13044 6752 13814 6780
rect 14369 6783 14427 6789
rect 13044 6740 13050 6752
rect 14369 6749 14381 6783
rect 14415 6780 14427 6783
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 14415 6752 16405 6780
rect 14415 6749 14427 6752
rect 14369 6743 14427 6749
rect 16393 6749 16405 6752
rect 16439 6780 16451 6783
rect 16574 6780 16580 6792
rect 16439 6752 16580 6780
rect 16439 6749 16451 6752
rect 16393 6743 16451 6749
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 18230 6780 18236 6792
rect 18191 6752 18236 6780
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 17313 6715 17371 6721
rect 17313 6681 17325 6715
rect 17359 6712 17371 6715
rect 18782 6712 18788 6724
rect 17359 6684 18092 6712
rect 18743 6684 18788 6712
rect 17359 6681 17371 6684
rect 17313 6675 17371 6681
rect 10870 6644 10876 6656
rect 10831 6616 10876 6644
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 13170 6644 13176 6656
rect 13131 6616 13176 6644
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 18064 6653 18092 6684
rect 18782 6672 18788 6684
rect 18840 6672 18846 6724
rect 18049 6647 18107 6653
rect 18049 6613 18061 6647
rect 18095 6644 18107 6647
rect 18138 6644 18144 6656
rect 18095 6616 18144 6644
rect 18095 6613 18107 6616
rect 18049 6607 18107 6613
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 9398 6400 9404 6452
rect 9456 6440 9462 6452
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 9456 6412 9689 6440
rect 9456 6400 9462 6412
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 10318 6440 10324 6452
rect 10231 6412 10324 6440
rect 9677 6403 9735 6409
rect 10318 6400 10324 6412
rect 10376 6440 10382 6452
rect 12158 6440 12164 6452
rect 10376 6412 12164 6440
rect 10376 6400 10382 6412
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 12621 6443 12679 6449
rect 12621 6409 12633 6443
rect 12667 6440 12679 6443
rect 12802 6440 12808 6452
rect 12667 6412 12808 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 13262 6400 13268 6452
rect 13320 6440 13326 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 13320 6412 13461 6440
rect 13320 6400 13326 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13449 6403 13507 6409
rect 16485 6443 16543 6449
rect 16485 6409 16497 6443
rect 16531 6440 16543 6443
rect 16666 6440 16672 6452
rect 16531 6412 16672 6440
rect 16531 6409 16543 6412
rect 16485 6403 16543 6409
rect 10870 6372 10876 6384
rect 10831 6344 10876 6372
rect 10870 6332 10876 6344
rect 10928 6332 10934 6384
rect 11330 6372 11336 6384
rect 10980 6344 11336 6372
rect 4798 6264 4804 6316
rect 4856 6304 4862 6316
rect 10980 6304 11008 6344
rect 11330 6332 11336 6344
rect 11388 6372 11394 6384
rect 11793 6375 11851 6381
rect 11793 6372 11805 6375
rect 11388 6344 11805 6372
rect 11388 6332 11394 6344
rect 11793 6341 11805 6344
rect 11839 6341 11851 6375
rect 11793 6335 11851 6341
rect 11238 6304 11244 6316
rect 4856 6276 11008 6304
rect 11199 6276 11244 6304
rect 4856 6264 4862 6276
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 11808 6304 11836 6335
rect 11808 6276 12480 6304
rect 9309 6239 9367 6245
rect 9309 6205 9321 6239
rect 9355 6236 9367 6239
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 9355 6208 9597 6236
rect 9355 6205 9367 6208
rect 9309 6199 9367 6205
rect 9585 6205 9597 6208
rect 9631 6205 9643 6239
rect 9585 6199 9643 6205
rect 9398 6168 9404 6180
rect 9359 6140 9404 6168
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 9600 6168 9628 6199
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10744 6208 10793 6236
rect 10744 6196 10750 6208
rect 10781 6205 10793 6208
rect 10827 6205 10839 6239
rect 10781 6199 10839 6205
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 11146 6236 11152 6248
rect 11103 6208 11152 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 11072 6168 11100 6199
rect 11146 6196 11152 6208
rect 11204 6236 11210 6248
rect 12452 6245 12480 6276
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11204 6208 12173 6236
rect 11204 6196 11210 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12897 6239 12955 6245
rect 12897 6236 12909 6239
rect 12483 6208 12909 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12897 6205 12909 6208
rect 12943 6205 12955 6239
rect 13464 6236 13492 6403
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 16850 6440 16856 6452
rect 16811 6412 16856 6440
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 19518 6400 19524 6452
rect 19576 6440 19582 6452
rect 19705 6443 19763 6449
rect 19705 6440 19717 6443
rect 19576 6412 19717 6440
rect 19576 6400 19582 6412
rect 19705 6409 19717 6412
rect 19751 6409 19763 6443
rect 19705 6403 19763 6409
rect 15473 6375 15531 6381
rect 15473 6341 15485 6375
rect 15519 6372 15531 6375
rect 16868 6372 16896 6400
rect 15519 6344 16896 6372
rect 15519 6341 15531 6344
rect 15473 6335 15531 6341
rect 14366 6264 14372 6316
rect 14424 6304 14430 6316
rect 14553 6307 14611 6313
rect 14553 6304 14565 6307
rect 14424 6276 14565 6304
rect 14424 6264 14430 6276
rect 14553 6273 14565 6276
rect 14599 6304 14611 6307
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 14599 6276 15025 6304
rect 14599 6273 14611 6276
rect 14553 6267 14611 6273
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 13464 6208 13645 6236
rect 12897 6199 12955 6205
rect 13633 6205 13645 6208
rect 13679 6205 13691 6239
rect 13633 6199 13691 6205
rect 14461 6239 14519 6245
rect 14461 6205 14473 6239
rect 14507 6205 14519 6239
rect 14461 6199 14519 6205
rect 14737 6239 14795 6245
rect 14737 6205 14749 6239
rect 14783 6236 14795 6239
rect 15562 6236 15568 6248
rect 14783 6208 15568 6236
rect 14783 6205 14795 6208
rect 14737 6199 14795 6205
rect 9600 6140 11100 6168
rect 12802 6128 12808 6180
rect 12860 6168 12866 6180
rect 13998 6168 14004 6180
rect 12860 6140 14004 6168
rect 12860 6128 12866 6140
rect 13998 6128 14004 6140
rect 14056 6168 14062 6180
rect 14476 6168 14504 6199
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 15901 6177 15929 6344
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 17911 6276 18061 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 18049 6273 18061 6276
rect 18095 6304 18107 6307
rect 18322 6304 18328 6316
rect 18095 6276 18328 6304
rect 18095 6273 18107 6276
rect 18049 6267 18107 6273
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 17497 6239 17555 6245
rect 17497 6205 17509 6239
rect 17543 6236 17555 6239
rect 18138 6236 18144 6248
rect 17543 6208 18144 6236
rect 17543 6205 17555 6208
rect 17497 6199 17555 6205
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 14056 6140 14504 6168
rect 15886 6171 15944 6177
rect 14056 6128 14062 6140
rect 15886 6137 15898 6171
rect 15932 6137 15944 6171
rect 15886 6131 15944 6137
rect 10686 6100 10692 6112
rect 10647 6072 10692 6100
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 9398 5896 9404 5908
rect 9359 5868 9404 5896
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 12986 5896 12992 5908
rect 12947 5868 12992 5896
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13446 5896 13452 5908
rect 13407 5868 13452 5896
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 14366 5896 14372 5908
rect 14327 5868 14372 5896
rect 14366 5856 14372 5868
rect 14424 5856 14430 5908
rect 15470 5896 15476 5908
rect 15431 5868 15476 5896
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 16209 5899 16267 5905
rect 16209 5896 16221 5899
rect 15620 5868 16221 5896
rect 15620 5856 15626 5868
rect 16209 5865 16221 5868
rect 16255 5865 16267 5899
rect 16574 5896 16580 5908
rect 16535 5868 16580 5896
rect 16209 5859 16267 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 18230 5896 18236 5908
rect 18191 5868 18236 5896
rect 18230 5856 18236 5868
rect 18288 5896 18294 5908
rect 18325 5899 18383 5905
rect 18325 5896 18337 5899
rect 18288 5868 18337 5896
rect 18288 5856 18294 5868
rect 18325 5865 18337 5868
rect 18371 5865 18383 5899
rect 18325 5859 18383 5865
rect 9416 5828 9444 5856
rect 10962 5828 10968 5840
rect 9416 5800 10968 5828
rect 10962 5788 10968 5800
rect 11020 5828 11026 5840
rect 11885 5831 11943 5837
rect 11020 5800 11100 5828
rect 11020 5788 11026 5800
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 11072 5769 11100 5800
rect 11885 5797 11897 5831
rect 11931 5828 11943 5831
rect 12894 5828 12900 5840
rect 11931 5800 12900 5828
rect 11931 5797 11943 5800
rect 11885 5791 11943 5797
rect 12894 5788 12900 5800
rect 12952 5788 12958 5840
rect 13173 5831 13231 5837
rect 13173 5797 13185 5831
rect 13219 5828 13231 5831
rect 13262 5828 13268 5840
rect 13219 5800 13268 5828
rect 13219 5797 13231 5800
rect 13173 5791 13231 5797
rect 13262 5788 13268 5800
rect 13320 5828 13326 5840
rect 14001 5831 14059 5837
rect 14001 5828 14013 5831
rect 13320 5800 14013 5828
rect 13320 5788 13326 5800
rect 14001 5797 14013 5800
rect 14047 5797 14059 5831
rect 16942 5828 16948 5840
rect 16903 5800 16948 5828
rect 14001 5791 14059 5797
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 17494 5828 17500 5840
rect 17455 5800 17500 5828
rect 17494 5788 17500 5800
rect 17552 5788 17558 5840
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 10744 5732 10885 5760
rect 10744 5720 10750 5732
rect 10873 5729 10885 5732
rect 10919 5729 10931 5763
rect 10873 5723 10931 5729
rect 11057 5763 11115 5769
rect 11057 5729 11069 5763
rect 11103 5729 11115 5763
rect 11422 5760 11428 5772
rect 11383 5732 11428 5760
rect 11057 5723 11115 5729
rect 10888 5692 10916 5723
rect 11422 5720 11428 5732
rect 11480 5720 11486 5772
rect 12912 5760 12940 5788
rect 13357 5763 13415 5769
rect 13357 5760 13369 5763
rect 12912 5732 13369 5760
rect 13357 5729 13369 5732
rect 13403 5760 13415 5763
rect 13538 5760 13544 5772
rect 13403 5732 13544 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 15746 5760 15752 5772
rect 15707 5732 15752 5760
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 11514 5692 11520 5704
rect 10888 5664 11520 5692
rect 11514 5652 11520 5664
rect 11572 5652 11578 5704
rect 16850 5692 16856 5704
rect 16811 5664 16856 5692
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 13170 5584 13176 5636
rect 13228 5624 13234 5636
rect 16758 5624 16764 5636
rect 13228 5596 16764 5624
rect 13228 5584 13234 5596
rect 16758 5584 16764 5596
rect 16816 5584 16822 5636
rect 15933 5559 15991 5565
rect 15933 5525 15945 5559
rect 15979 5556 15991 5559
rect 17218 5556 17224 5568
rect 15979 5528 17224 5556
rect 15979 5525 15991 5528
rect 15933 5519 15991 5525
rect 17218 5516 17224 5528
rect 17276 5516 17282 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 10962 5312 10968 5364
rect 11020 5352 11026 5364
rect 11793 5355 11851 5361
rect 11793 5352 11805 5355
rect 11020 5324 11805 5352
rect 11020 5312 11026 5324
rect 11793 5321 11805 5324
rect 11839 5321 11851 5355
rect 13262 5352 13268 5364
rect 13223 5324 13268 5352
rect 11793 5315 11851 5321
rect 13262 5312 13268 5324
rect 13320 5312 13326 5364
rect 13538 5352 13544 5364
rect 13499 5324 13544 5352
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 13998 5352 14004 5364
rect 13959 5324 14004 5352
rect 13998 5312 14004 5324
rect 14056 5312 14062 5364
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 16117 5355 16175 5361
rect 16117 5352 16129 5355
rect 15804 5324 16129 5352
rect 15804 5312 15810 5324
rect 16117 5321 16129 5324
rect 16163 5321 16175 5355
rect 16117 5315 16175 5321
rect 14461 5287 14519 5293
rect 14461 5253 14473 5287
rect 14507 5284 14519 5287
rect 15838 5284 15844 5296
rect 14507 5256 15844 5284
rect 14507 5253 14519 5256
rect 14461 5247 14519 5253
rect 15838 5244 15844 5256
rect 15896 5244 15902 5296
rect 11146 5216 11152 5228
rect 11107 5188 11152 5216
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 17000 5188 17049 5216
rect 17000 5176 17006 5188
rect 17037 5185 17049 5188
rect 17083 5216 17095 5219
rect 17313 5219 17371 5225
rect 17313 5216 17325 5219
rect 17083 5188 17325 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 17313 5185 17325 5188
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 9858 5148 9864 5160
rect 9819 5120 9864 5148
rect 9858 5108 9864 5120
rect 9916 5148 9922 5160
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 9916 5120 10241 5148
rect 9916 5108 9922 5120
rect 10229 5117 10241 5120
rect 10275 5148 10287 5151
rect 10505 5151 10563 5157
rect 10505 5148 10517 5151
rect 10275 5120 10517 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 10505 5117 10517 5120
rect 10551 5148 10563 5151
rect 11422 5148 11428 5160
rect 10551 5120 11428 5148
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 13872 5120 14289 5148
rect 13872 5108 13878 5120
rect 14277 5117 14289 5120
rect 14323 5148 14335 5151
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 14323 5120 14749 5148
rect 14323 5117 14335 5120
rect 14277 5111 14335 5117
rect 14737 5117 14749 5120
rect 14783 5117 14795 5151
rect 15286 5148 15292 5160
rect 15247 5120 15292 5148
rect 14737 5111 14795 5117
rect 15286 5108 15292 5120
rect 15344 5148 15350 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15344 5120 15761 5148
rect 15344 5108 15350 5120
rect 15749 5117 15761 5120
rect 15795 5117 15807 5151
rect 16666 5148 16672 5160
rect 16627 5120 16672 5148
rect 15749 5111 15807 5117
rect 16666 5108 16672 5120
rect 16724 5108 16730 5160
rect 11514 5012 11520 5024
rect 11475 4984 11520 5012
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 15473 5015 15531 5021
rect 15473 4981 15485 5015
rect 15519 5012 15531 5015
rect 18874 5012 18880 5024
rect 15519 4984 18880 5012
rect 15519 4981 15531 4984
rect 15473 4975 15531 4981
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 10962 4808 10968 4820
rect 10923 4780 10968 4808
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 16623 4811 16681 4817
rect 16623 4777 16635 4811
rect 16669 4808 16681 4811
rect 16850 4808 16856 4820
rect 16669 4780 16856 4808
rect 16669 4777 16681 4780
rect 16623 4771 16681 4777
rect 16850 4768 16856 4780
rect 16908 4808 16914 4820
rect 16945 4811 17003 4817
rect 16945 4808 16957 4811
rect 16908 4780 16957 4808
rect 16908 4768 16914 4780
rect 16945 4777 16957 4780
rect 16991 4777 17003 4811
rect 16945 4771 17003 4777
rect 21959 4811 22017 4817
rect 21959 4777 21971 4811
rect 22005 4808 22017 4811
rect 22370 4808 22376 4820
rect 22005 4780 22376 4808
rect 22005 4777 22017 4780
rect 21959 4771 22017 4777
rect 22370 4768 22376 4780
rect 22428 4768 22434 4820
rect 10870 4672 10876 4684
rect 10831 4644 10876 4672
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 16574 4681 16580 4684
rect 16552 4675 16580 4681
rect 16552 4672 16564 4675
rect 16487 4644 16564 4672
rect 16552 4641 16564 4644
rect 16632 4672 16638 4684
rect 17678 4672 17684 4684
rect 16632 4644 17684 4672
rect 16552 4635 16580 4641
rect 16574 4632 16580 4635
rect 16632 4632 16638 4644
rect 17678 4632 17684 4644
rect 17736 4632 17742 4684
rect 21726 4672 21732 4684
rect 21687 4644 21732 4672
rect 21726 4632 21732 4644
rect 21784 4632 21790 4684
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 16666 4604 16672 4616
rect 16439 4576 16672 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 16574 4264 16580 4276
rect 16535 4236 16580 4264
rect 16574 4224 16580 4236
rect 16632 4224 16638 4276
rect 21726 4224 21732 4276
rect 21784 4264 21790 4276
rect 21913 4267 21971 4273
rect 21913 4264 21925 4267
rect 21784 4236 21925 4264
rect 21784 4224 21790 4236
rect 21913 4233 21925 4236
rect 21959 4264 21971 4267
rect 27614 4264 27620 4276
rect 21959 4236 27620 4264
rect 21959 4233 21971 4236
rect 21913 4227 21971 4233
rect 27614 4224 27620 4236
rect 27672 4224 27678 4276
rect 10778 3924 10784 3936
rect 10739 3896 10784 3924
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 106 3544 112 3596
rect 164 3584 170 3596
rect 1394 3584 1400 3596
rect 1452 3593 1458 3596
rect 1452 3587 1490 3593
rect 164 3556 1400 3584
rect 164 3544 170 3556
rect 1394 3544 1400 3556
rect 1478 3553 1490 3587
rect 1452 3547 1490 3553
rect 1452 3544 1458 3547
rect 1535 3519 1593 3525
rect 1535 3485 1547 3519
rect 1581 3516 1593 3519
rect 11330 3516 11336 3528
rect 1581 3488 11336 3516
rect 1581 3485 1593 3488
rect 1535 3479 1593 3485
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1452 3148 1593 3176
rect 1452 3136 1458 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 1581 3139 1639 3145
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 24118 2592 24124 2644
rect 24176 2632 24182 2644
rect 24719 2635 24777 2641
rect 24719 2632 24731 2635
rect 24176 2604 24731 2632
rect 24176 2592 24182 2604
rect 24719 2601 24731 2604
rect 24765 2601 24777 2635
rect 24719 2595 24777 2601
rect 24648 2499 24706 2505
rect 24648 2465 24660 2499
rect 24694 2496 24706 2499
rect 25130 2496 25136 2508
rect 24694 2468 25136 2496
rect 24694 2465 24706 2468
rect 24648 2459 24706 2465
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 25130 2292 25136 2304
rect 25091 2264 25136 2292
rect 25130 2252 25136 2264
rect 25188 2252 25194 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 19426 76 19432 128
rect 19484 116 19490 128
rect 20070 116 20076 128
rect 19484 88 20076 116
rect 19484 76 19490 88
rect 20070 76 20076 88
rect 20128 76 20134 128
<< via1 >>
rect 4804 27480 4856 27532
rect 6460 27480 6512 27532
rect 9680 27480 9732 27532
rect 10416 27480 10468 27532
rect 13636 27480 13688 27532
rect 16028 27480 16080 27532
rect 2044 27072 2096 27124
rect 6000 27072 6052 27124
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 3424 25100 3476 25152
rect 6920 25100 6972 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 24768 24871 24820 24880
rect 24768 24837 24777 24871
rect 24777 24837 24811 24871
rect 24811 24837 24820 24871
rect 24768 24828 24820 24837
rect 24032 24692 24084 24744
rect 664 24556 716 24608
rect 6276 24556 6328 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1584 24395 1636 24404
rect 1584 24361 1593 24395
rect 1593 24361 1627 24395
rect 1627 24361 1636 24395
rect 1584 24352 1636 24361
rect 18788 24352 18840 24404
rect 25504 24352 25556 24404
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 17592 24259 17644 24268
rect 17592 24225 17601 24259
rect 17601 24225 17635 24259
rect 17635 24225 17644 24259
rect 17592 24216 17644 24225
rect 23480 24259 23532 24268
rect 23480 24225 23489 24259
rect 23489 24225 23523 24259
rect 23523 24225 23532 24259
rect 23480 24216 23532 24225
rect 24676 24216 24728 24268
rect 25780 24080 25832 24132
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1400 23808 1452 23860
rect 2044 23808 2096 23860
rect 12992 23851 13044 23860
rect 12992 23817 13001 23851
rect 13001 23817 13035 23851
rect 13035 23817 13044 23851
rect 12992 23808 13044 23817
rect 14556 23851 14608 23860
rect 14556 23817 14565 23851
rect 14565 23817 14599 23851
rect 14599 23817 14608 23851
rect 14556 23808 14608 23817
rect 17408 23808 17460 23860
rect 17592 23851 17644 23860
rect 17592 23817 17601 23851
rect 17601 23817 17635 23851
rect 17635 23817 17644 23851
rect 17592 23808 17644 23817
rect 21640 23808 21692 23860
rect 23020 23808 23072 23860
rect 23480 23808 23532 23860
rect 23848 23851 23900 23860
rect 23848 23817 23857 23851
rect 23857 23817 23891 23851
rect 23891 23817 23900 23851
rect 23848 23808 23900 23817
rect 27160 23808 27212 23860
rect 1492 23740 1544 23792
rect 20168 23740 20220 23792
rect 23480 23672 23532 23724
rect 24676 23672 24728 23724
rect 12992 23604 13044 23656
rect 14556 23604 14608 23656
rect 16396 23647 16448 23656
rect 16396 23613 16405 23647
rect 16405 23613 16439 23647
rect 16439 23613 16448 23647
rect 16396 23604 16448 23613
rect 19248 23647 19300 23656
rect 19248 23613 19257 23647
rect 19257 23613 19291 23647
rect 19291 23613 19300 23647
rect 19248 23604 19300 23613
rect 19524 23604 19576 23656
rect 20260 23536 20312 23588
rect 24032 23536 24084 23588
rect 2964 23468 3016 23520
rect 12348 23468 12400 23520
rect 13544 23468 13596 23520
rect 24216 23468 24268 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1584 23307 1636 23316
rect 1584 23273 1593 23307
rect 1593 23273 1627 23307
rect 1627 23273 1636 23307
rect 1584 23264 1636 23273
rect 15108 23264 15160 23316
rect 16396 23264 16448 23316
rect 24124 23264 24176 23316
rect 25228 23264 25280 23316
rect 1400 23171 1452 23180
rect 1400 23137 1409 23171
rect 1409 23137 1443 23171
rect 1443 23137 1452 23171
rect 1400 23128 1452 23137
rect 11152 23128 11204 23180
rect 15292 23128 15344 23180
rect 23296 23171 23348 23180
rect 23296 23137 23305 23171
rect 23305 23137 23339 23171
rect 23339 23137 23348 23171
rect 23296 23128 23348 23137
rect 24124 23128 24176 23180
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 23296 22763 23348 22772
rect 23296 22729 23305 22763
rect 23305 22729 23339 22763
rect 23339 22729 23348 22763
rect 23296 22720 23348 22729
rect 24768 22763 24820 22772
rect 24768 22729 24777 22763
rect 24777 22729 24811 22763
rect 24811 22729 24820 22763
rect 24768 22720 24820 22729
rect 23388 22516 23440 22568
rect 24124 22516 24176 22568
rect 1400 22380 1452 22432
rect 9036 22380 9088 22432
rect 11152 22380 11204 22432
rect 13912 22380 13964 22432
rect 15292 22423 15344 22432
rect 15292 22389 15301 22423
rect 15301 22389 15335 22423
rect 15335 22389 15344 22423
rect 15292 22380 15344 22389
rect 23296 22380 23348 22432
rect 24032 22380 24084 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1952 22040 2004 22092
rect 2044 22040 2096 22092
rect 3056 22040 3108 22092
rect 3516 21904 3568 21956
rect 1768 21836 1820 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1492 21632 1544 21684
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 3056 21539 3108 21548
rect 3056 21505 3065 21539
rect 3065 21505 3099 21539
rect 3099 21505 3108 21539
rect 3056 21496 3108 21505
rect 24676 21428 24728 21480
rect 4988 21360 5040 21412
rect 1952 21335 2004 21344
rect 1952 21301 1961 21335
rect 1961 21301 1995 21335
rect 1995 21301 2004 21335
rect 1952 21292 2004 21301
rect 2504 21335 2556 21344
rect 2504 21301 2513 21335
rect 2513 21301 2547 21335
rect 2547 21301 2556 21335
rect 2504 21292 2556 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1584 21131 1636 21140
rect 1584 21097 1593 21131
rect 1593 21097 1627 21131
rect 1627 21097 1636 21131
rect 1584 21088 1636 21097
rect 2044 20952 2096 21004
rect 1216 20884 1268 20936
rect 3332 20884 3384 20936
rect 2136 20748 2188 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1308 20544 1360 20596
rect 3332 20587 3384 20596
rect 3332 20553 3341 20587
rect 3341 20553 3375 20587
rect 3375 20553 3384 20587
rect 3332 20544 3384 20553
rect 24860 20544 24912 20596
rect 2964 20340 3016 20392
rect 3792 20408 3844 20460
rect 9680 20408 9732 20460
rect 3976 20383 4028 20392
rect 3976 20349 3985 20383
rect 3985 20349 4019 20383
rect 4019 20349 4028 20383
rect 3976 20340 4028 20349
rect 3148 20272 3200 20324
rect 24124 20340 24176 20392
rect 2044 20247 2096 20256
rect 2044 20213 2053 20247
rect 2053 20213 2087 20247
rect 2087 20213 2096 20247
rect 2044 20204 2096 20213
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 2872 20204 2924 20256
rect 9864 20204 9916 20256
rect 9956 20204 10008 20256
rect 16304 20204 16356 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 204 20000 256 20052
rect 2412 20000 2464 20052
rect 4988 20000 5040 20052
rect 19248 19932 19300 19984
rect 22468 19932 22520 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 2780 19864 2832 19916
rect 4620 19864 4672 19916
rect 5356 19864 5408 19916
rect 6092 19864 6144 19916
rect 7656 19864 7708 19916
rect 8024 19864 8076 19916
rect 8944 19864 8996 19916
rect 11428 19864 11480 19916
rect 14004 19864 14056 19916
rect 15568 19864 15620 19916
rect 18052 19907 18104 19916
rect 18052 19873 18061 19907
rect 18061 19873 18095 19907
rect 18095 19873 18104 19907
rect 18052 19864 18104 19873
rect 18604 19907 18656 19916
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 19432 19864 19484 19916
rect 18788 19839 18840 19848
rect 18788 19805 18797 19839
rect 18797 19805 18831 19839
rect 18831 19805 18840 19839
rect 18788 19796 18840 19805
rect 2688 19771 2740 19780
rect 2688 19737 2697 19771
rect 2697 19737 2731 19771
rect 2731 19737 2740 19771
rect 2688 19728 2740 19737
rect 13728 19728 13780 19780
rect 17868 19728 17920 19780
rect 19248 19728 19300 19780
rect 4620 19703 4672 19712
rect 4620 19669 4629 19703
rect 4629 19669 4663 19703
rect 4663 19669 4672 19703
rect 4620 19660 4672 19669
rect 7932 19660 7984 19712
rect 8484 19660 8536 19712
rect 10140 19660 10192 19712
rect 10968 19660 11020 19712
rect 14188 19660 14240 19712
rect 16212 19703 16264 19712
rect 16212 19669 16221 19703
rect 16221 19669 16255 19703
rect 16255 19669 16264 19703
rect 16212 19660 16264 19669
rect 19984 19660 20036 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 7656 19499 7708 19508
rect 7656 19465 7665 19499
rect 7665 19465 7699 19499
rect 7699 19465 7708 19499
rect 7656 19456 7708 19465
rect 8024 19456 8076 19508
rect 8944 19499 8996 19508
rect 8944 19465 8953 19499
rect 8953 19465 8987 19499
rect 8987 19465 8996 19499
rect 8944 19456 8996 19465
rect 13636 19499 13688 19508
rect 13636 19465 13645 19499
rect 13645 19465 13679 19499
rect 13679 19465 13688 19499
rect 13636 19456 13688 19465
rect 15752 19456 15804 19508
rect 18052 19456 18104 19508
rect 24768 19499 24820 19508
rect 24768 19465 24777 19499
rect 24777 19465 24811 19499
rect 24811 19465 24820 19499
rect 24768 19456 24820 19465
rect 1676 19252 1728 19304
rect 2044 19252 2096 19304
rect 4712 19320 4764 19372
rect 6920 19320 6972 19372
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 19432 19363 19484 19372
rect 19432 19329 19441 19363
rect 19441 19329 19475 19363
rect 19475 19329 19484 19363
rect 19432 19320 19484 19329
rect 1492 19184 1544 19236
rect 2780 19184 2832 19236
rect 204 19116 256 19168
rect 2412 19116 2464 19168
rect 3700 19116 3752 19168
rect 3884 19159 3936 19168
rect 3884 19125 3893 19159
rect 3893 19125 3927 19159
rect 3927 19125 3936 19159
rect 3884 19116 3936 19125
rect 4344 19116 4396 19168
rect 4988 19184 5040 19236
rect 8944 19252 8996 19304
rect 4804 19116 4856 19168
rect 5356 19159 5408 19168
rect 5356 19125 5365 19159
rect 5365 19125 5399 19159
rect 5399 19125 5408 19159
rect 5356 19116 5408 19125
rect 7196 19116 7248 19168
rect 8116 19116 8168 19168
rect 9312 19116 9364 19168
rect 11428 19295 11480 19304
rect 11428 19261 11446 19295
rect 11446 19261 11480 19295
rect 11428 19252 11480 19261
rect 13728 19252 13780 19304
rect 14372 19252 14424 19304
rect 14648 19252 14700 19304
rect 17500 19252 17552 19304
rect 18604 19295 18656 19304
rect 18604 19261 18613 19295
rect 18613 19261 18647 19295
rect 18647 19261 18656 19295
rect 18604 19252 18656 19261
rect 19248 19252 19300 19304
rect 20076 19295 20128 19304
rect 20076 19261 20085 19295
rect 20085 19261 20119 19295
rect 20119 19261 20128 19295
rect 20076 19252 20128 19261
rect 20720 19252 20772 19304
rect 15292 19227 15344 19236
rect 15292 19193 15301 19227
rect 15301 19193 15335 19227
rect 15335 19193 15344 19227
rect 15292 19184 15344 19193
rect 16212 19227 16264 19236
rect 16212 19193 16221 19227
rect 16221 19193 16255 19227
rect 16255 19193 16264 19227
rect 16212 19184 16264 19193
rect 9772 19116 9824 19168
rect 12992 19116 13044 19168
rect 13452 19116 13504 19168
rect 14004 19116 14056 19168
rect 15568 19159 15620 19168
rect 15568 19125 15577 19159
rect 15577 19125 15611 19159
rect 15611 19125 15620 19159
rect 15568 19116 15620 19125
rect 16488 19184 16540 19236
rect 16948 19184 17000 19236
rect 17040 19184 17092 19236
rect 17500 19159 17552 19168
rect 17500 19125 17509 19159
rect 17509 19125 17543 19159
rect 17543 19125 17552 19159
rect 17500 19116 17552 19125
rect 18144 19159 18196 19168
rect 18144 19125 18153 19159
rect 18153 19125 18187 19159
rect 18187 19125 18196 19159
rect 18144 19116 18196 19125
rect 18972 19184 19024 19236
rect 19064 19159 19116 19168
rect 19064 19125 19073 19159
rect 19073 19125 19107 19159
rect 19107 19125 19116 19159
rect 19064 19116 19116 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 3884 18912 3936 18964
rect 4988 18912 5040 18964
rect 6276 18912 6328 18964
rect 7656 18912 7708 18964
rect 12348 18912 12400 18964
rect 18420 18912 18472 18964
rect 2228 18844 2280 18896
rect 3424 18844 3476 18896
rect 4896 18844 4948 18896
rect 6552 18844 6604 18896
rect 16304 18887 16356 18896
rect 16304 18853 16313 18887
rect 16313 18853 16347 18887
rect 16347 18853 16356 18887
rect 16304 18844 16356 18853
rect 16396 18887 16448 18896
rect 16396 18853 16405 18887
rect 16405 18853 16439 18887
rect 16439 18853 16448 18887
rect 16948 18887 17000 18896
rect 16396 18844 16448 18853
rect 16948 18853 16957 18887
rect 16957 18853 16991 18887
rect 16991 18853 17000 18887
rect 16948 18844 17000 18853
rect 17868 18887 17920 18896
rect 17868 18853 17877 18887
rect 17877 18853 17911 18887
rect 17911 18853 17920 18887
rect 17868 18844 17920 18853
rect 18052 18844 18104 18896
rect 19064 18912 19116 18964
rect 20076 18912 20128 18964
rect 23388 18912 23440 18964
rect 21088 18887 21140 18896
rect 21088 18853 21097 18887
rect 21097 18853 21131 18887
rect 21131 18853 21140 18887
rect 21088 18844 21140 18853
rect 6092 18776 6144 18828
rect 8024 18776 8076 18828
rect 9680 18776 9732 18828
rect 11704 18776 11756 18828
rect 12164 18776 12216 18828
rect 13820 18819 13872 18828
rect 13820 18785 13829 18819
rect 13829 18785 13863 18819
rect 13863 18785 13872 18819
rect 13820 18776 13872 18785
rect 14556 18776 14608 18828
rect 19892 18776 19944 18828
rect 23112 18819 23164 18828
rect 23112 18785 23121 18819
rect 23121 18785 23155 18819
rect 23155 18785 23164 18819
rect 23112 18776 23164 18785
rect 2504 18708 2556 18760
rect 2596 18708 2648 18760
rect 3056 18708 3108 18760
rect 4160 18751 4212 18760
rect 4160 18717 4169 18751
rect 4169 18717 4203 18751
rect 4203 18717 4212 18751
rect 4620 18751 4672 18760
rect 4160 18708 4212 18717
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 7564 18708 7616 18760
rect 14832 18708 14884 18760
rect 8300 18640 8352 18692
rect 20812 18708 20864 18760
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 24124 18640 24176 18692
rect 1676 18615 1728 18624
rect 1676 18581 1685 18615
rect 1685 18581 1719 18615
rect 1719 18581 1728 18615
rect 1676 18572 1728 18581
rect 2320 18572 2372 18624
rect 6552 18615 6604 18624
rect 6552 18581 6561 18615
rect 6561 18581 6595 18615
rect 6595 18581 6604 18615
rect 6552 18572 6604 18581
rect 7288 18572 7340 18624
rect 10324 18572 10376 18624
rect 10876 18572 10928 18624
rect 14464 18572 14516 18624
rect 14556 18572 14608 18624
rect 15660 18572 15712 18624
rect 20168 18572 20220 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2504 18368 2556 18420
rect 4160 18368 4212 18420
rect 6092 18368 6144 18420
rect 8024 18368 8076 18420
rect 9680 18411 9732 18420
rect 9680 18377 9689 18411
rect 9689 18377 9723 18411
rect 9723 18377 9732 18411
rect 9680 18368 9732 18377
rect 16396 18368 16448 18420
rect 3424 18343 3476 18352
rect 3424 18309 3433 18343
rect 3433 18309 3467 18343
rect 3467 18309 3476 18343
rect 4896 18343 4948 18352
rect 3424 18300 3476 18309
rect 2412 18275 2464 18284
rect 2412 18241 2421 18275
rect 2421 18241 2455 18275
rect 2455 18241 2464 18275
rect 2412 18232 2464 18241
rect 3056 18275 3108 18284
rect 3056 18241 3065 18275
rect 3065 18241 3099 18275
rect 3099 18241 3108 18275
rect 3056 18232 3108 18241
rect 4896 18309 4905 18343
rect 4905 18309 4939 18343
rect 4939 18309 4948 18343
rect 4896 18300 4948 18309
rect 6460 18300 6512 18352
rect 7840 18300 7892 18352
rect 17868 18368 17920 18420
rect 17960 18368 18012 18420
rect 21088 18368 21140 18420
rect 22744 18368 22796 18420
rect 24860 18368 24912 18420
rect 20444 18300 20496 18352
rect 20812 18300 20864 18352
rect 10324 18275 10376 18284
rect 1860 18139 1912 18148
rect 1860 18105 1869 18139
rect 1869 18105 1903 18139
rect 1903 18105 1912 18139
rect 1860 18096 1912 18105
rect 3976 18139 4028 18148
rect 3976 18105 3985 18139
rect 3985 18105 4019 18139
rect 4019 18105 4028 18139
rect 3976 18096 4028 18105
rect 4068 18139 4120 18148
rect 4068 18105 4077 18139
rect 4077 18105 4111 18139
rect 4111 18105 4120 18139
rect 4620 18139 4672 18148
rect 4068 18096 4120 18105
rect 4620 18105 4629 18139
rect 4629 18105 4663 18139
rect 4663 18105 4672 18139
rect 4620 18096 4672 18105
rect 3884 18028 3936 18080
rect 6000 18164 6052 18216
rect 6276 18207 6328 18216
rect 6276 18173 6285 18207
rect 6285 18173 6319 18207
rect 6319 18173 6328 18207
rect 6276 18164 6328 18173
rect 8300 18164 8352 18216
rect 10324 18241 10333 18275
rect 10333 18241 10367 18275
rect 10367 18241 10376 18275
rect 10324 18232 10376 18241
rect 10692 18275 10744 18284
rect 10692 18241 10701 18275
rect 10701 18241 10735 18275
rect 10735 18241 10744 18275
rect 10692 18232 10744 18241
rect 12348 18232 12400 18284
rect 6920 18139 6972 18148
rect 6920 18105 6929 18139
rect 6929 18105 6963 18139
rect 6963 18105 6972 18139
rect 6920 18096 6972 18105
rect 7564 18139 7616 18148
rect 7564 18105 7573 18139
rect 7573 18105 7607 18139
rect 7607 18105 7616 18139
rect 7564 18096 7616 18105
rect 11612 18164 11664 18216
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 13268 18164 13320 18216
rect 14372 18207 14424 18216
rect 14372 18173 14381 18207
rect 14381 18173 14415 18207
rect 14415 18173 14424 18207
rect 14372 18164 14424 18173
rect 14464 18164 14516 18216
rect 15844 18232 15896 18284
rect 17040 18232 17092 18284
rect 18420 18275 18472 18284
rect 18420 18241 18429 18275
rect 18429 18241 18463 18275
rect 18463 18241 18472 18275
rect 18420 18232 18472 18241
rect 21456 18275 21508 18284
rect 15660 18164 15712 18216
rect 21456 18241 21465 18275
rect 21465 18241 21499 18275
rect 21499 18241 21508 18275
rect 23112 18275 23164 18284
rect 21456 18232 21508 18241
rect 23112 18241 23121 18275
rect 23121 18241 23155 18275
rect 23155 18241 23164 18275
rect 23112 18232 23164 18241
rect 23572 18164 23624 18216
rect 7104 18028 7156 18080
rect 7932 18071 7984 18080
rect 7932 18037 7941 18071
rect 7941 18037 7975 18071
rect 7975 18037 7984 18071
rect 12532 18096 12584 18148
rect 13360 18096 13412 18148
rect 14556 18096 14608 18148
rect 15476 18096 15528 18148
rect 18512 18139 18564 18148
rect 18512 18105 18521 18139
rect 18521 18105 18555 18139
rect 18555 18105 18564 18139
rect 19892 18139 19944 18148
rect 18512 18096 18564 18105
rect 19892 18105 19901 18139
rect 19901 18105 19935 18139
rect 19935 18105 19944 18139
rect 19892 18096 19944 18105
rect 20352 18096 20404 18148
rect 21180 18139 21232 18148
rect 21180 18105 21189 18139
rect 21189 18105 21223 18139
rect 21223 18105 21232 18139
rect 21180 18096 21232 18105
rect 7932 18028 7984 18037
rect 11704 18028 11756 18080
rect 15568 18071 15620 18080
rect 15568 18037 15577 18071
rect 15577 18037 15611 18071
rect 15611 18037 15620 18071
rect 15568 18028 15620 18037
rect 17224 18028 17276 18080
rect 18052 18028 18104 18080
rect 20076 18071 20128 18080
rect 20076 18037 20085 18071
rect 20085 18037 20119 18071
rect 20119 18037 20128 18071
rect 20076 18028 20128 18037
rect 20536 18071 20588 18080
rect 20536 18037 20545 18071
rect 20545 18037 20579 18071
rect 20579 18037 20588 18071
rect 20536 18028 20588 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2412 17824 2464 17876
rect 3884 17824 3936 17876
rect 4068 17824 4120 17876
rect 6460 17867 6512 17876
rect 6460 17833 6469 17867
rect 6469 17833 6503 17867
rect 6503 17833 6512 17867
rect 6460 17824 6512 17833
rect 6920 17824 6972 17876
rect 9772 17867 9824 17876
rect 9772 17833 9781 17867
rect 9781 17833 9815 17867
rect 9815 17833 9824 17867
rect 9772 17824 9824 17833
rect 10876 17867 10928 17876
rect 10876 17833 10885 17867
rect 10885 17833 10919 17867
rect 10919 17833 10928 17867
rect 10876 17824 10928 17833
rect 14464 17867 14516 17876
rect 14464 17833 14473 17867
rect 14473 17833 14507 17867
rect 14507 17833 14516 17867
rect 14464 17824 14516 17833
rect 16304 17824 16356 17876
rect 17684 17867 17736 17876
rect 17684 17833 17693 17867
rect 17693 17833 17727 17867
rect 17727 17833 17736 17867
rect 17684 17824 17736 17833
rect 18512 17867 18564 17876
rect 18512 17833 18521 17867
rect 18521 17833 18555 17867
rect 18555 17833 18564 17867
rect 18512 17824 18564 17833
rect 18972 17867 19024 17876
rect 18972 17833 18981 17867
rect 18981 17833 19015 17867
rect 19015 17833 19024 17867
rect 19432 17867 19484 17876
rect 18972 17824 19024 17833
rect 2044 17756 2096 17808
rect 4160 17756 4212 17808
rect 7104 17756 7156 17808
rect 8208 17799 8260 17808
rect 8208 17765 8217 17799
rect 8217 17765 8251 17799
rect 8251 17765 8260 17799
rect 8208 17756 8260 17765
rect 6552 17688 6604 17740
rect 10048 17756 10100 17808
rect 11888 17756 11940 17808
rect 13176 17799 13228 17808
rect 13176 17765 13185 17799
rect 13185 17765 13219 17799
rect 13219 17765 13228 17799
rect 13176 17756 13228 17765
rect 15568 17756 15620 17808
rect 9864 17688 9916 17740
rect 17224 17688 17276 17740
rect 18144 17688 18196 17740
rect 19432 17833 19441 17867
rect 19441 17833 19475 17867
rect 19475 17833 19484 17867
rect 19432 17824 19484 17833
rect 21180 17824 21232 17876
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 21088 17799 21140 17808
rect 21088 17765 21097 17799
rect 21097 17765 21131 17799
rect 21131 17765 21140 17799
rect 21088 17756 21140 17765
rect 22376 17756 22428 17808
rect 23204 17799 23256 17808
rect 23204 17765 23213 17799
rect 23213 17765 23247 17799
rect 23247 17765 23256 17799
rect 23204 17756 23256 17765
rect 24124 17688 24176 17740
rect 3148 17620 3200 17672
rect 3424 17620 3476 17672
rect 5172 17620 5224 17672
rect 6000 17620 6052 17672
rect 7564 17620 7616 17672
rect 10692 17620 10744 17672
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 13360 17620 13412 17672
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 15384 17663 15436 17672
rect 15384 17629 15393 17663
rect 15393 17629 15427 17663
rect 15427 17629 15436 17663
rect 15384 17620 15436 17629
rect 21272 17620 21324 17672
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 22560 17663 22612 17672
rect 22560 17629 22569 17663
rect 22569 17629 22603 17663
rect 22603 17629 22612 17663
rect 22560 17620 22612 17629
rect 2596 17595 2648 17604
rect 2596 17561 2605 17595
rect 2605 17561 2639 17595
rect 2639 17561 2648 17595
rect 2596 17552 2648 17561
rect 3976 17552 4028 17604
rect 4620 17552 4672 17604
rect 11060 17552 11112 17604
rect 13820 17552 13872 17604
rect 20628 17552 20680 17604
rect 23480 17552 23532 17604
rect 11336 17484 11388 17536
rect 12532 17484 12584 17536
rect 12624 17484 12676 17536
rect 15568 17484 15620 17536
rect 18052 17484 18104 17536
rect 20904 17484 20956 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2044 17323 2096 17332
rect 2044 17289 2053 17323
rect 2053 17289 2087 17323
rect 2087 17289 2096 17323
rect 2044 17280 2096 17289
rect 3424 17323 3476 17332
rect 3424 17289 3433 17323
rect 3433 17289 3467 17323
rect 3467 17289 3476 17323
rect 3424 17280 3476 17289
rect 4896 17280 4948 17332
rect 7104 17280 7156 17332
rect 9864 17280 9916 17332
rect 13176 17280 13228 17332
rect 16488 17280 16540 17332
rect 8208 17212 8260 17264
rect 2872 17144 2924 17196
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 4252 17119 4304 17128
rect 4252 17085 4261 17119
rect 4261 17085 4295 17119
rect 4295 17085 4304 17119
rect 4252 17076 4304 17085
rect 6460 17144 6512 17196
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 2044 16940 2096 16992
rect 4160 16983 4212 16992
rect 4160 16949 4169 16983
rect 4169 16949 4203 16983
rect 4203 16949 4212 16983
rect 6000 17008 6052 17060
rect 6920 17008 6972 17060
rect 7656 17144 7708 17196
rect 10876 17187 10928 17196
rect 10876 17153 10885 17187
rect 10885 17153 10919 17187
rect 10919 17153 10928 17187
rect 10876 17144 10928 17153
rect 13452 17212 13504 17264
rect 18144 17280 18196 17332
rect 20076 17280 20128 17332
rect 15384 17144 15436 17196
rect 9772 17076 9824 17128
rect 11980 17076 12032 17128
rect 12624 17076 12676 17128
rect 15476 17119 15528 17128
rect 7932 17008 7984 17060
rect 4160 16940 4212 16949
rect 10048 16940 10100 16992
rect 11336 17008 11388 17060
rect 11520 17051 11572 17060
rect 11520 17017 11529 17051
rect 11529 17017 11563 17051
rect 11563 17017 11572 17051
rect 11520 17008 11572 17017
rect 11888 17051 11940 17060
rect 11888 17017 11897 17051
rect 11897 17017 11931 17051
rect 11931 17017 11940 17051
rect 11888 17008 11940 17017
rect 15476 17085 15485 17119
rect 15485 17085 15519 17119
rect 15519 17085 15528 17119
rect 15476 17076 15528 17085
rect 17960 17212 18012 17264
rect 20536 17212 20588 17264
rect 18788 17144 18840 17196
rect 20076 17144 20128 17196
rect 20444 17187 20496 17196
rect 20444 17153 20453 17187
rect 20453 17153 20487 17187
rect 20487 17153 20496 17187
rect 20444 17144 20496 17153
rect 21088 17280 21140 17332
rect 23112 17323 23164 17332
rect 23112 17289 23121 17323
rect 23121 17289 23155 17323
rect 23155 17289 23164 17323
rect 23112 17280 23164 17289
rect 20904 17212 20956 17264
rect 23848 17212 23900 17264
rect 21272 17144 21324 17196
rect 23204 17144 23256 17196
rect 17684 17008 17736 17060
rect 19432 17008 19484 17060
rect 23112 17076 23164 17128
rect 22376 17051 22428 17060
rect 22376 17017 22385 17051
rect 22385 17017 22419 17051
rect 22419 17017 22428 17051
rect 22376 17008 22428 17017
rect 23756 17051 23808 17060
rect 23756 17017 23765 17051
rect 23765 17017 23799 17051
rect 23799 17017 23808 17051
rect 23756 17008 23808 17017
rect 23848 17051 23900 17060
rect 23848 17017 23857 17051
rect 23857 17017 23891 17051
rect 23891 17017 23900 17051
rect 23848 17008 23900 17017
rect 13452 16940 13504 16992
rect 13728 16940 13780 16992
rect 17776 16940 17828 16992
rect 19064 16983 19116 16992
rect 19064 16949 19073 16983
rect 19073 16949 19107 16983
rect 19107 16949 19116 16983
rect 19064 16940 19116 16949
rect 22560 16940 22612 16992
rect 24124 16940 24176 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2872 16736 2924 16788
rect 3516 16779 3568 16788
rect 3516 16745 3525 16779
rect 3525 16745 3559 16779
rect 3559 16745 3568 16779
rect 3516 16736 3568 16745
rect 4252 16736 4304 16788
rect 7564 16736 7616 16788
rect 8300 16779 8352 16788
rect 8300 16745 8309 16779
rect 8309 16745 8343 16779
rect 8343 16745 8352 16779
rect 8300 16736 8352 16745
rect 9772 16736 9824 16788
rect 11244 16779 11296 16788
rect 11244 16745 11253 16779
rect 11253 16745 11287 16779
rect 11287 16745 11296 16779
rect 11244 16736 11296 16745
rect 11520 16736 11572 16788
rect 12716 16736 12768 16788
rect 15384 16779 15436 16788
rect 15384 16745 15393 16779
rect 15393 16745 15427 16779
rect 15427 16745 15436 16779
rect 15384 16736 15436 16745
rect 15476 16736 15528 16788
rect 16488 16736 16540 16788
rect 17776 16736 17828 16788
rect 20812 16736 20864 16788
rect 20904 16736 20956 16788
rect 2228 16711 2280 16720
rect 2228 16677 2237 16711
rect 2237 16677 2271 16711
rect 2271 16677 2280 16711
rect 2228 16668 2280 16677
rect 3056 16668 3108 16720
rect 6828 16668 6880 16720
rect 11980 16668 12032 16720
rect 4620 16643 4672 16652
rect 4620 16609 4629 16643
rect 4629 16609 4663 16643
rect 4663 16609 4672 16643
rect 4620 16600 4672 16609
rect 4988 16643 5040 16652
rect 4988 16609 4997 16643
rect 4997 16609 5031 16643
rect 5031 16609 5040 16643
rect 4988 16600 5040 16609
rect 1584 16396 1636 16448
rect 6092 16464 6144 16516
rect 7104 16600 7156 16652
rect 8024 16643 8076 16652
rect 8024 16609 8033 16643
rect 8033 16609 8067 16643
rect 8067 16609 8076 16643
rect 8024 16600 8076 16609
rect 8300 16600 8352 16652
rect 9864 16600 9916 16652
rect 10048 16600 10100 16652
rect 10232 16643 10284 16652
rect 10232 16609 10241 16643
rect 10241 16609 10275 16643
rect 10275 16609 10284 16643
rect 10232 16600 10284 16609
rect 10784 16643 10836 16652
rect 10784 16609 10793 16643
rect 10793 16609 10827 16643
rect 10827 16609 10836 16643
rect 10784 16600 10836 16609
rect 11888 16600 11940 16652
rect 15660 16668 15712 16720
rect 13912 16643 13964 16652
rect 13912 16609 13921 16643
rect 13921 16609 13955 16643
rect 13955 16609 13964 16643
rect 13912 16600 13964 16609
rect 14464 16600 14516 16652
rect 15476 16643 15528 16652
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 15844 16643 15896 16652
rect 15844 16609 15853 16643
rect 15853 16609 15887 16643
rect 15887 16609 15896 16643
rect 15844 16600 15896 16609
rect 17776 16600 17828 16652
rect 19248 16668 19300 16720
rect 20076 16668 20128 16720
rect 20168 16668 20220 16720
rect 22560 16736 22612 16788
rect 24676 16736 24728 16788
rect 22744 16668 22796 16720
rect 23204 16711 23256 16720
rect 23204 16677 23213 16711
rect 23213 16677 23247 16711
rect 23247 16677 23256 16711
rect 23204 16668 23256 16677
rect 18604 16643 18656 16652
rect 18604 16609 18613 16643
rect 18613 16609 18647 16643
rect 18647 16609 18656 16643
rect 18604 16600 18656 16609
rect 19800 16643 19852 16652
rect 19800 16609 19809 16643
rect 19809 16609 19843 16643
rect 19843 16609 19852 16643
rect 19800 16600 19852 16609
rect 20628 16600 20680 16652
rect 23940 16643 23992 16652
rect 23940 16609 23949 16643
rect 23949 16609 23983 16643
rect 23983 16609 23992 16643
rect 23940 16600 23992 16609
rect 25596 16600 25648 16652
rect 11060 16532 11112 16584
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 14280 16532 14332 16584
rect 19432 16532 19484 16584
rect 21272 16575 21324 16584
rect 21272 16541 21281 16575
rect 21281 16541 21315 16575
rect 21315 16541 21324 16575
rect 21272 16532 21324 16541
rect 22560 16575 22612 16584
rect 22560 16541 22569 16575
rect 22569 16541 22603 16575
rect 22603 16541 22612 16575
rect 22560 16532 22612 16541
rect 23756 16575 23808 16584
rect 23756 16541 23765 16575
rect 23765 16541 23799 16575
rect 23799 16541 23808 16575
rect 23756 16532 23808 16541
rect 10140 16464 10192 16516
rect 17040 16464 17092 16516
rect 4160 16396 4212 16448
rect 4528 16396 4580 16448
rect 12808 16396 12860 16448
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 17592 16396 17644 16448
rect 18236 16396 18288 16448
rect 19064 16396 19116 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1860 16235 1912 16244
rect 1860 16201 1869 16235
rect 1869 16201 1903 16235
rect 1903 16201 1912 16235
rect 1860 16192 1912 16201
rect 2228 16192 2280 16244
rect 6092 16235 6144 16244
rect 6092 16201 6101 16235
rect 6101 16201 6135 16235
rect 6135 16201 6144 16235
rect 6092 16192 6144 16201
rect 8024 16235 8076 16244
rect 8024 16201 8033 16235
rect 8033 16201 8067 16235
rect 8067 16201 8076 16235
rect 8024 16192 8076 16201
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 14464 16192 14516 16244
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 20904 16192 20956 16244
rect 22560 16192 22612 16244
rect 2596 16167 2648 16176
rect 2596 16133 2605 16167
rect 2605 16133 2639 16167
rect 2639 16133 2648 16167
rect 2596 16124 2648 16133
rect 4620 16124 4672 16176
rect 10692 16124 10744 16176
rect 11244 16124 11296 16176
rect 2136 16056 2188 16108
rect 3056 16056 3108 16108
rect 4988 16099 5040 16108
rect 4988 16065 4997 16099
rect 4997 16065 5031 16099
rect 5031 16065 5040 16099
rect 10232 16099 10284 16108
rect 4988 16056 5040 16065
rect 5264 16031 5316 16040
rect 5264 15997 5273 16031
rect 5273 15997 5307 16031
rect 5307 15997 5316 16031
rect 5264 15988 5316 15997
rect 1860 15920 1912 15972
rect 3608 15963 3660 15972
rect 3608 15929 3617 15963
rect 3617 15929 3651 15963
rect 3651 15929 3660 15963
rect 3608 15920 3660 15929
rect 3424 15895 3476 15904
rect 3424 15861 3433 15895
rect 3433 15861 3467 15895
rect 3467 15861 3476 15895
rect 4620 15895 4672 15904
rect 3424 15852 3476 15861
rect 4620 15861 4629 15895
rect 4629 15861 4663 15895
rect 4663 15861 4672 15895
rect 4620 15852 4672 15861
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 6368 15852 6420 15904
rect 7104 15988 7156 16040
rect 8300 15988 8352 16040
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 6920 15895 6972 15904
rect 6920 15861 6929 15895
rect 6929 15861 6963 15895
rect 6963 15861 6972 15895
rect 6920 15852 6972 15861
rect 8392 15852 8444 15904
rect 9680 15988 9732 16040
rect 11060 16031 11112 16040
rect 11060 15997 11069 16031
rect 11069 15997 11103 16031
rect 11103 15997 11112 16031
rect 11060 15988 11112 15997
rect 14924 15988 14976 16040
rect 15752 16056 15804 16108
rect 18604 16124 18656 16176
rect 21364 16167 21416 16176
rect 21364 16133 21373 16167
rect 21373 16133 21407 16167
rect 21407 16133 21416 16167
rect 21364 16124 21416 16133
rect 22744 16167 22796 16176
rect 22744 16133 22753 16167
rect 22753 16133 22787 16167
rect 22787 16133 22796 16167
rect 22744 16124 22796 16133
rect 23940 16192 23992 16244
rect 24584 16124 24636 16176
rect 16488 16099 16540 16108
rect 16488 16065 16497 16099
rect 16497 16065 16531 16099
rect 16531 16065 16540 16099
rect 16488 16056 16540 16065
rect 17960 16056 18012 16108
rect 19800 16099 19852 16108
rect 19800 16065 19809 16099
rect 19809 16065 19843 16099
rect 19843 16065 19852 16099
rect 19800 16056 19852 16065
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 24860 16056 24912 16108
rect 27620 16056 27672 16108
rect 12808 15963 12860 15972
rect 12808 15929 12817 15963
rect 12817 15929 12851 15963
rect 12851 15929 12860 15963
rect 12808 15920 12860 15929
rect 13452 15920 13504 15972
rect 15568 15963 15620 15972
rect 8852 15895 8904 15904
rect 8852 15861 8861 15895
rect 8861 15861 8895 15895
rect 8895 15861 8904 15895
rect 8852 15852 8904 15861
rect 10784 15852 10836 15904
rect 11060 15852 11112 15904
rect 13912 15852 13964 15904
rect 14556 15852 14608 15904
rect 15568 15929 15577 15963
rect 15577 15929 15611 15963
rect 15611 15929 15620 15963
rect 15568 15920 15620 15929
rect 16580 15963 16632 15972
rect 16580 15929 16589 15963
rect 16589 15929 16623 15963
rect 16623 15929 16632 15963
rect 16580 15920 16632 15929
rect 17592 15920 17644 15972
rect 18696 15963 18748 15972
rect 18696 15929 18705 15963
rect 18705 15929 18739 15963
rect 18739 15929 18748 15963
rect 19248 15963 19300 15972
rect 18696 15920 18748 15929
rect 19248 15929 19257 15963
rect 19257 15929 19291 15963
rect 19291 15929 19300 15963
rect 19248 15920 19300 15929
rect 15476 15852 15528 15904
rect 15936 15895 15988 15904
rect 15936 15861 15945 15895
rect 15945 15861 15979 15895
rect 15979 15861 15988 15895
rect 15936 15852 15988 15861
rect 17776 15895 17828 15904
rect 17776 15861 17785 15895
rect 17785 15861 17819 15895
rect 17819 15861 17828 15895
rect 17776 15852 17828 15861
rect 20536 15895 20588 15904
rect 20536 15861 20545 15895
rect 20545 15861 20579 15895
rect 20579 15861 20588 15895
rect 22284 15895 22336 15904
rect 20536 15852 20588 15861
rect 22284 15861 22293 15895
rect 22293 15861 22327 15895
rect 22327 15861 22336 15895
rect 22284 15852 22336 15861
rect 23940 15852 23992 15904
rect 24676 15852 24728 15904
rect 25596 15895 25648 15904
rect 25596 15861 25605 15895
rect 25605 15861 25639 15895
rect 25639 15861 25648 15895
rect 25596 15852 25648 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2044 15648 2096 15700
rect 3056 15691 3108 15700
rect 3056 15657 3065 15691
rect 3065 15657 3099 15691
rect 3099 15657 3108 15691
rect 3056 15648 3108 15657
rect 3424 15648 3476 15700
rect 8300 15691 8352 15700
rect 2504 15580 2556 15632
rect 2688 15623 2740 15632
rect 2688 15589 2697 15623
rect 2697 15589 2731 15623
rect 2731 15589 2740 15623
rect 2688 15580 2740 15589
rect 3976 15580 4028 15632
rect 4988 15580 5040 15632
rect 5448 15580 5500 15632
rect 7104 15623 7156 15632
rect 7104 15589 7113 15623
rect 7113 15589 7147 15623
rect 7147 15589 7156 15623
rect 7104 15580 7156 15589
rect 7288 15623 7340 15632
rect 7288 15589 7297 15623
rect 7297 15589 7331 15623
rect 7331 15589 7340 15623
rect 7288 15580 7340 15589
rect 8300 15657 8309 15691
rect 8309 15657 8343 15691
rect 8343 15657 8352 15691
rect 8300 15648 8352 15657
rect 9680 15648 9732 15700
rect 14924 15691 14976 15700
rect 14924 15657 14933 15691
rect 14933 15657 14967 15691
rect 14967 15657 14976 15691
rect 14924 15648 14976 15657
rect 15844 15648 15896 15700
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 18236 15691 18288 15700
rect 16120 15648 16172 15657
rect 18236 15657 18245 15691
rect 18245 15657 18279 15691
rect 18279 15657 18288 15691
rect 18236 15648 18288 15657
rect 18696 15648 18748 15700
rect 19432 15691 19484 15700
rect 19432 15657 19441 15691
rect 19441 15657 19475 15691
rect 19475 15657 19484 15691
rect 19432 15648 19484 15657
rect 20812 15648 20864 15700
rect 23940 15691 23992 15700
rect 23940 15657 23949 15691
rect 23949 15657 23983 15691
rect 23983 15657 23992 15691
rect 23940 15648 23992 15657
rect 24584 15648 24636 15700
rect 7748 15580 7800 15632
rect 9864 15623 9916 15632
rect 9864 15589 9873 15623
rect 9873 15589 9907 15623
rect 9907 15589 9916 15623
rect 9864 15580 9916 15589
rect 11060 15580 11112 15632
rect 13084 15623 13136 15632
rect 5264 15512 5316 15564
rect 2412 15444 2464 15496
rect 3516 15444 3568 15496
rect 10692 15512 10744 15564
rect 11244 15555 11296 15564
rect 11244 15521 11253 15555
rect 11253 15521 11287 15555
rect 11287 15521 11296 15555
rect 11244 15512 11296 15521
rect 13084 15589 13093 15623
rect 13093 15589 13127 15623
rect 13127 15589 13136 15623
rect 13084 15580 13136 15589
rect 13452 15580 13504 15632
rect 21088 15623 21140 15632
rect 21088 15589 21097 15623
rect 21097 15589 21131 15623
rect 21131 15589 21140 15623
rect 21088 15580 21140 15589
rect 23112 15623 23164 15632
rect 23112 15589 23121 15623
rect 23121 15589 23155 15623
rect 23155 15589 23164 15623
rect 23112 15580 23164 15589
rect 18052 15512 18104 15564
rect 20260 15512 20312 15564
rect 3332 15376 3384 15428
rect 5540 15444 5592 15496
rect 8208 15444 8260 15496
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 11796 15487 11848 15496
rect 11796 15453 11805 15487
rect 11805 15453 11839 15487
rect 11839 15453 11848 15487
rect 11796 15444 11848 15453
rect 13820 15444 13872 15496
rect 14280 15444 14332 15496
rect 14372 15444 14424 15496
rect 17224 15444 17276 15496
rect 17868 15487 17920 15496
rect 17868 15453 17877 15487
rect 17877 15453 17911 15487
rect 17911 15453 17920 15487
rect 17868 15444 17920 15453
rect 21364 15444 21416 15496
rect 23480 15444 23532 15496
rect 4436 15308 4488 15360
rect 5356 15308 5408 15360
rect 8576 15308 8628 15360
rect 11060 15308 11112 15360
rect 12716 15351 12768 15360
rect 12716 15317 12725 15351
rect 12725 15317 12759 15351
rect 12759 15317 12768 15351
rect 12716 15308 12768 15317
rect 12900 15308 12952 15360
rect 14924 15376 14976 15428
rect 19248 15376 19300 15428
rect 23848 15580 23900 15632
rect 24768 15512 24820 15564
rect 16672 15351 16724 15360
rect 16672 15317 16681 15351
rect 16681 15317 16715 15351
rect 16715 15317 16724 15351
rect 16672 15308 16724 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 4528 15104 4580 15156
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 9864 15147 9916 15156
rect 9864 15113 9873 15147
rect 9873 15113 9907 15147
rect 9907 15113 9916 15147
rect 9864 15104 9916 15113
rect 11888 15104 11940 15156
rect 13084 15104 13136 15156
rect 13820 15147 13872 15156
rect 13820 15113 13829 15147
rect 13829 15113 13863 15147
rect 13863 15113 13872 15147
rect 17224 15147 17276 15156
rect 13820 15104 13872 15113
rect 17224 15113 17233 15147
rect 17233 15113 17267 15147
rect 17267 15113 17276 15147
rect 17224 15104 17276 15113
rect 20628 15104 20680 15156
rect 21088 15104 21140 15156
rect 23112 15104 23164 15156
rect 2044 15036 2096 15088
rect 5448 15036 5500 15088
rect 9772 15036 9824 15088
rect 15568 15036 15620 15088
rect 2688 15011 2740 15020
rect 2688 14977 2697 15011
rect 2697 14977 2731 15011
rect 2731 14977 2740 15011
rect 2688 14968 2740 14977
rect 3332 15011 3384 15020
rect 3332 14977 3341 15011
rect 3341 14977 3375 15011
rect 3375 14977 3384 15011
rect 3332 14968 3384 14977
rect 1860 14943 1912 14952
rect 1860 14909 1869 14943
rect 1869 14909 1903 14943
rect 1903 14909 1912 14943
rect 1860 14900 1912 14909
rect 1952 14832 2004 14884
rect 2964 14832 3016 14884
rect 4436 14900 4488 14952
rect 8852 14968 8904 15020
rect 10876 14968 10928 15020
rect 11244 14968 11296 15020
rect 12900 14968 12952 15020
rect 14832 14968 14884 15020
rect 18236 14968 18288 15020
rect 6920 14900 6972 14952
rect 12716 14900 12768 14952
rect 13636 14900 13688 14952
rect 19432 14968 19484 15020
rect 20260 14968 20312 15020
rect 23480 15036 23532 15088
rect 23848 15036 23900 15088
rect 23940 14968 23992 15020
rect 24768 15011 24820 15020
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 24768 14968 24820 14977
rect 27620 14968 27672 15020
rect 2412 14764 2464 14816
rect 2504 14764 2556 14816
rect 4068 14832 4120 14884
rect 4252 14832 4304 14884
rect 4528 14807 4580 14816
rect 4528 14773 4537 14807
rect 4537 14773 4571 14807
rect 4571 14773 4580 14807
rect 4528 14764 4580 14773
rect 6460 14832 6512 14884
rect 9864 14832 9916 14884
rect 10692 14764 10744 14816
rect 13452 14832 13504 14884
rect 16120 14832 16172 14884
rect 14556 14764 14608 14816
rect 16580 14807 16632 14816
rect 16580 14773 16589 14807
rect 16589 14773 16623 14807
rect 16623 14773 16632 14807
rect 16580 14764 16632 14773
rect 17684 14764 17736 14816
rect 19432 14832 19484 14884
rect 22836 14900 22888 14952
rect 20076 14832 20128 14884
rect 20720 14764 20772 14816
rect 24492 14832 24544 14884
rect 25780 14807 25832 14816
rect 25780 14773 25789 14807
rect 25789 14773 25823 14807
rect 25823 14773 25832 14807
rect 25780 14764 25832 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2964 14603 3016 14612
rect 2964 14569 2973 14603
rect 2973 14569 3007 14603
rect 3007 14569 3016 14603
rect 2964 14560 3016 14569
rect 3516 14603 3568 14612
rect 3516 14569 3525 14603
rect 3525 14569 3559 14603
rect 3559 14569 3568 14603
rect 3516 14560 3568 14569
rect 4528 14603 4580 14612
rect 4528 14569 4537 14603
rect 4537 14569 4571 14603
rect 4571 14569 4580 14603
rect 4528 14560 4580 14569
rect 6460 14603 6512 14612
rect 6460 14569 6469 14603
rect 6469 14569 6503 14603
rect 6503 14569 6512 14603
rect 6460 14560 6512 14569
rect 7288 14560 7340 14612
rect 7748 14560 7800 14612
rect 1768 14492 1820 14544
rect 2044 14535 2096 14544
rect 2044 14501 2053 14535
rect 2053 14501 2087 14535
rect 2087 14501 2096 14535
rect 2044 14492 2096 14501
rect 2688 14492 2740 14544
rect 7196 14492 7248 14544
rect 7932 14535 7984 14544
rect 7932 14501 7941 14535
rect 7941 14501 7975 14535
rect 7975 14501 7984 14535
rect 7932 14492 7984 14501
rect 8852 14560 8904 14612
rect 10692 14560 10744 14612
rect 10876 14603 10928 14612
rect 10876 14569 10885 14603
rect 10885 14569 10919 14603
rect 10919 14569 10928 14603
rect 10876 14560 10928 14569
rect 13084 14603 13136 14612
rect 13084 14569 13093 14603
rect 13093 14569 13127 14603
rect 13127 14569 13136 14603
rect 13084 14560 13136 14569
rect 13636 14603 13688 14612
rect 13636 14569 13645 14603
rect 13645 14569 13679 14603
rect 13679 14569 13688 14603
rect 13636 14560 13688 14569
rect 18788 14560 18840 14612
rect 19984 14603 20036 14612
rect 19984 14569 19993 14603
rect 19993 14569 20027 14603
rect 20027 14569 20036 14603
rect 19984 14560 20036 14569
rect 20628 14603 20680 14612
rect 20628 14569 20637 14603
rect 20637 14569 20671 14603
rect 20671 14569 20680 14603
rect 20628 14560 20680 14569
rect 9864 14492 9916 14544
rect 11888 14492 11940 14544
rect 12164 14535 12216 14544
rect 12164 14501 12173 14535
rect 12173 14501 12207 14535
rect 12207 14501 12216 14535
rect 12164 14492 12216 14501
rect 16120 14492 16172 14544
rect 16672 14492 16724 14544
rect 17408 14492 17460 14544
rect 17684 14492 17736 14544
rect 20168 14492 20220 14544
rect 22284 14560 22336 14612
rect 21088 14535 21140 14544
rect 21088 14501 21097 14535
rect 21097 14501 21131 14535
rect 21131 14501 21140 14535
rect 21088 14492 21140 14501
rect 22928 14492 22980 14544
rect 23848 14535 23900 14544
rect 23848 14501 23857 14535
rect 23857 14501 23891 14535
rect 23891 14501 23900 14535
rect 23848 14492 23900 14501
rect 24860 14535 24912 14544
rect 24860 14501 24869 14535
rect 24869 14501 24903 14535
rect 24903 14501 24912 14535
rect 24860 14492 24912 14501
rect 4344 14424 4396 14476
rect 5448 14424 5500 14476
rect 7748 14424 7800 14476
rect 13820 14467 13872 14476
rect 13820 14433 13829 14467
rect 13829 14433 13863 14467
rect 13863 14433 13872 14467
rect 14004 14467 14056 14476
rect 13820 14424 13872 14433
rect 14004 14433 14013 14467
rect 14013 14433 14047 14467
rect 14047 14433 14056 14467
rect 14004 14424 14056 14433
rect 15292 14424 15344 14476
rect 18880 14467 18932 14476
rect 18880 14433 18889 14467
rect 18889 14433 18923 14467
rect 18923 14433 18932 14467
rect 18880 14424 18932 14433
rect 19248 14424 19300 14476
rect 2044 14356 2096 14408
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 12348 14356 12400 14408
rect 12716 14399 12768 14408
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 13360 14356 13412 14408
rect 17040 14356 17092 14408
rect 17592 14356 17644 14408
rect 21364 14399 21416 14408
rect 21364 14365 21373 14399
rect 21373 14365 21407 14399
rect 21407 14365 21416 14399
rect 21364 14356 21416 14365
rect 24492 14356 24544 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 25044 14399 25096 14408
rect 25044 14365 25053 14399
rect 25053 14365 25087 14399
rect 25087 14365 25096 14399
rect 25044 14356 25096 14365
rect 3976 14288 4028 14340
rect 10968 14288 11020 14340
rect 13268 14288 13320 14340
rect 20536 14288 20588 14340
rect 22928 14288 22980 14340
rect 4068 14220 4120 14272
rect 5540 14220 5592 14272
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 7288 14220 7340 14229
rect 11060 14220 11112 14272
rect 16488 14263 16540 14272
rect 16488 14229 16497 14263
rect 16497 14229 16531 14263
rect 16531 14229 16540 14263
rect 16488 14220 16540 14229
rect 16856 14220 16908 14272
rect 17868 14220 17920 14272
rect 22652 14263 22704 14272
rect 22652 14229 22661 14263
rect 22661 14229 22695 14263
rect 22695 14229 22704 14263
rect 22652 14220 22704 14229
rect 23296 14220 23348 14272
rect 23848 14220 23900 14272
rect 24952 14220 25004 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1768 14059 1820 14068
rect 1768 14025 1777 14059
rect 1777 14025 1811 14059
rect 1811 14025 1820 14059
rect 1768 14016 1820 14025
rect 7748 14016 7800 14068
rect 8024 14016 8076 14068
rect 9864 14059 9916 14068
rect 1676 13744 1728 13796
rect 3516 13880 3568 13932
rect 6000 13948 6052 14000
rect 6276 13948 6328 14000
rect 9864 14025 9873 14059
rect 9873 14025 9907 14059
rect 9907 14025 9916 14059
rect 9864 14016 9916 14025
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 16120 14016 16172 14068
rect 17040 14016 17092 14068
rect 18880 14059 18932 14068
rect 18880 14025 18889 14059
rect 18889 14025 18923 14059
rect 18923 14025 18932 14059
rect 18880 14016 18932 14025
rect 21088 14016 21140 14068
rect 6092 13880 6144 13932
rect 2136 13744 2188 13796
rect 2596 13744 2648 13796
rect 1492 13676 1544 13728
rect 3516 13787 3568 13796
rect 3516 13753 3525 13787
rect 3525 13753 3559 13787
rect 3559 13753 3568 13787
rect 3516 13744 3568 13753
rect 3424 13676 3476 13728
rect 5172 13744 5224 13796
rect 6368 13812 6420 13864
rect 7104 13812 7156 13864
rect 7288 13855 7340 13864
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 8576 13812 8628 13864
rect 9680 13880 9732 13932
rect 8852 13812 8904 13864
rect 10968 13855 11020 13864
rect 10968 13821 10977 13855
rect 10977 13821 11011 13855
rect 11011 13821 11020 13855
rect 10968 13812 11020 13821
rect 11060 13812 11112 13864
rect 14004 13948 14056 14000
rect 14740 13948 14792 14000
rect 17500 13948 17552 14000
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 16856 13880 16908 13932
rect 17592 13880 17644 13932
rect 19984 13948 20036 14000
rect 20168 13948 20220 14000
rect 20904 13948 20956 14000
rect 21364 13991 21416 14000
rect 21364 13957 21373 13991
rect 21373 13957 21407 13991
rect 21407 13957 21416 13991
rect 21364 13948 21416 13957
rect 22284 14016 22336 14068
rect 24124 14016 24176 14068
rect 24860 14016 24912 14068
rect 24952 14016 25004 14068
rect 22836 13948 22888 14000
rect 22928 13948 22980 14000
rect 19432 13880 19484 13932
rect 20444 13880 20496 13932
rect 23848 13880 23900 13932
rect 23940 13880 23992 13932
rect 24768 13880 24820 13932
rect 13820 13812 13872 13864
rect 14464 13812 14516 13864
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 18512 13855 18564 13864
rect 9864 13744 9916 13796
rect 11428 13744 11480 13796
rect 12532 13787 12584 13796
rect 12532 13753 12541 13787
rect 12541 13753 12575 13787
rect 12575 13753 12584 13787
rect 12532 13744 12584 13753
rect 14556 13787 14608 13796
rect 6000 13676 6052 13728
rect 6368 13676 6420 13728
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 7104 13676 7156 13728
rect 12164 13676 12216 13728
rect 14556 13753 14565 13787
rect 14565 13753 14599 13787
rect 14599 13753 14608 13787
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 20260 13812 20312 13864
rect 22652 13812 22704 13864
rect 16396 13787 16448 13796
rect 14556 13744 14608 13753
rect 14280 13676 14332 13728
rect 16396 13753 16405 13787
rect 16405 13753 16439 13787
rect 16439 13753 16448 13787
rect 16396 13744 16448 13753
rect 16488 13787 16540 13796
rect 16488 13753 16497 13787
rect 16497 13753 16531 13787
rect 16531 13753 16540 13787
rect 16488 13744 16540 13753
rect 19708 13744 19760 13796
rect 19984 13744 20036 13796
rect 20904 13787 20956 13796
rect 20904 13753 20913 13787
rect 20913 13753 20947 13787
rect 20947 13753 20956 13787
rect 20904 13744 20956 13753
rect 25780 13787 25832 13796
rect 25780 13753 25789 13787
rect 25789 13753 25823 13787
rect 25823 13753 25832 13787
rect 25780 13744 25832 13753
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17408 13676 17460 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2136 13472 2188 13524
rect 3516 13515 3568 13524
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 4344 13472 4396 13524
rect 5080 13472 5132 13524
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 7932 13515 7984 13524
rect 7932 13481 7941 13515
rect 7941 13481 7975 13515
rect 7975 13481 7984 13515
rect 7932 13472 7984 13481
rect 8024 13472 8076 13524
rect 2504 13404 2556 13456
rect 4252 13447 4304 13456
rect 4252 13413 4261 13447
rect 4261 13413 4295 13447
rect 4295 13413 4304 13447
rect 4252 13404 4304 13413
rect 6644 13447 6696 13456
rect 6644 13413 6653 13447
rect 6653 13413 6687 13447
rect 6687 13413 6696 13447
rect 6644 13404 6696 13413
rect 9404 13472 9456 13524
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 14740 13515 14792 13524
rect 14740 13481 14749 13515
rect 14749 13481 14783 13515
rect 14783 13481 14792 13515
rect 14740 13472 14792 13481
rect 15292 13472 15344 13524
rect 16396 13472 16448 13524
rect 19248 13472 19300 13524
rect 20444 13472 20496 13524
rect 23756 13515 23808 13524
rect 23756 13481 23765 13515
rect 23765 13481 23799 13515
rect 23799 13481 23808 13515
rect 23756 13472 23808 13481
rect 25044 13472 25096 13524
rect 11888 13404 11940 13456
rect 14372 13447 14424 13456
rect 14372 13413 14381 13447
rect 14381 13413 14415 13447
rect 14415 13413 14424 13447
rect 14372 13404 14424 13413
rect 19432 13447 19484 13456
rect 19432 13413 19441 13447
rect 19441 13413 19475 13447
rect 19475 13413 19484 13447
rect 19432 13404 19484 13413
rect 20260 13404 20312 13456
rect 20996 13447 21048 13456
rect 20996 13413 21005 13447
rect 21005 13413 21039 13447
rect 21039 13413 21048 13447
rect 20996 13404 21048 13413
rect 21088 13447 21140 13456
rect 21088 13413 21097 13447
rect 21097 13413 21131 13447
rect 21131 13413 21140 13447
rect 21088 13404 21140 13413
rect 22928 13404 22980 13456
rect 23480 13404 23532 13456
rect 24860 13404 24912 13456
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 2136 13268 2188 13320
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4528 13311 4580 13320
rect 4160 13268 4212 13277
rect 4528 13277 4537 13311
rect 4537 13277 4571 13311
rect 4571 13277 4580 13311
rect 4528 13268 4580 13277
rect 5540 13268 5592 13320
rect 7932 13268 7984 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 9220 13268 9272 13320
rect 12348 13336 12400 13388
rect 11428 13268 11480 13320
rect 13728 13336 13780 13388
rect 14556 13336 14608 13388
rect 15936 13379 15988 13388
rect 15936 13345 15945 13379
rect 15945 13345 15979 13379
rect 15979 13345 15988 13379
rect 15936 13336 15988 13345
rect 17868 13379 17920 13388
rect 17868 13345 17877 13379
rect 17877 13345 17911 13379
rect 17911 13345 17920 13379
rect 17868 13336 17920 13345
rect 14004 13268 14056 13320
rect 17224 13268 17276 13320
rect 18420 13311 18472 13320
rect 18420 13277 18429 13311
rect 18429 13277 18463 13311
rect 18463 13277 18472 13311
rect 18420 13268 18472 13277
rect 11336 13200 11388 13252
rect 12532 13200 12584 13252
rect 12992 13200 13044 13252
rect 22008 13268 22060 13320
rect 24216 13311 24268 13320
rect 19616 13200 19668 13252
rect 24216 13277 24225 13311
rect 24225 13277 24259 13311
rect 24259 13277 24268 13311
rect 24216 13268 24268 13277
rect 23204 13243 23256 13252
rect 23204 13209 23213 13243
rect 23213 13209 23247 13243
rect 23247 13209 23256 13243
rect 23204 13200 23256 13209
rect 6828 13132 6880 13184
rect 11060 13132 11112 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 22652 13132 22704 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 4252 12928 4304 12980
rect 5080 12928 5132 12980
rect 5264 12928 5316 12980
rect 8576 12928 8628 12980
rect 10140 12971 10192 12980
rect 10140 12937 10149 12971
rect 10149 12937 10183 12971
rect 10183 12937 10192 12971
rect 10140 12928 10192 12937
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 13728 12971 13780 12980
rect 13728 12937 13737 12971
rect 13737 12937 13771 12971
rect 13771 12937 13780 12971
rect 13728 12928 13780 12937
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 17132 12928 17184 12980
rect 17776 12971 17828 12980
rect 17776 12937 17785 12971
rect 17785 12937 17819 12971
rect 17819 12937 17828 12971
rect 17776 12928 17828 12937
rect 19616 12971 19668 12980
rect 19616 12937 19625 12971
rect 19625 12937 19659 12971
rect 19659 12937 19668 12971
rect 19616 12928 19668 12937
rect 20076 12971 20128 12980
rect 20076 12937 20085 12971
rect 20085 12937 20119 12971
rect 20119 12937 20128 12971
rect 20076 12928 20128 12937
rect 21088 12928 21140 12980
rect 23480 12971 23532 12980
rect 23480 12937 23489 12971
rect 23489 12937 23523 12971
rect 23523 12937 23532 12971
rect 23480 12928 23532 12937
rect 24216 12928 24268 12980
rect 2504 12860 2556 12912
rect 7012 12860 7064 12912
rect 9864 12903 9916 12912
rect 9864 12869 9873 12903
rect 9873 12869 9907 12903
rect 9907 12869 9916 12903
rect 9864 12860 9916 12869
rect 1952 12835 2004 12844
rect 1952 12801 1961 12835
rect 1961 12801 1995 12835
rect 1995 12801 2004 12835
rect 1952 12792 2004 12801
rect 2964 12792 3016 12844
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 4160 12792 4212 12844
rect 6736 12724 6788 12776
rect 8392 12724 8444 12776
rect 8760 12724 8812 12776
rect 14096 12860 14148 12912
rect 16028 12860 16080 12912
rect 19432 12860 19484 12912
rect 12716 12792 12768 12844
rect 13544 12792 13596 12844
rect 14556 12835 14608 12844
rect 11060 12724 11112 12776
rect 2596 12699 2648 12708
rect 2596 12665 2605 12699
rect 2605 12665 2639 12699
rect 2639 12665 2648 12699
rect 2596 12656 2648 12665
rect 3884 12699 3936 12708
rect 3884 12665 3886 12699
rect 3886 12665 3920 12699
rect 3920 12665 3936 12699
rect 3884 12656 3936 12665
rect 4528 12656 4580 12708
rect 5540 12631 5592 12640
rect 5540 12597 5549 12631
rect 5549 12597 5583 12631
rect 5583 12597 5592 12631
rect 5540 12588 5592 12597
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 6644 12588 6696 12597
rect 6828 12588 6880 12640
rect 7012 12699 7064 12708
rect 7012 12665 7021 12699
rect 7021 12665 7055 12699
rect 7055 12665 7064 12699
rect 7012 12656 7064 12665
rect 9772 12656 9824 12708
rect 11612 12656 11664 12708
rect 12532 12699 12584 12708
rect 12532 12665 12541 12699
rect 12541 12665 12575 12699
rect 12575 12665 12584 12699
rect 12532 12656 12584 12665
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 16304 12792 16356 12844
rect 14280 12699 14332 12708
rect 8024 12631 8076 12640
rect 8024 12597 8033 12631
rect 8033 12597 8067 12631
rect 8067 12597 8076 12631
rect 8024 12588 8076 12597
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 9496 12588 9548 12597
rect 12440 12588 12492 12640
rect 14280 12665 14289 12699
rect 14289 12665 14323 12699
rect 14323 12665 14332 12699
rect 14280 12656 14332 12665
rect 14740 12656 14792 12708
rect 15936 12699 15988 12708
rect 15936 12665 15945 12699
rect 15945 12665 15979 12699
rect 15979 12665 15988 12699
rect 15936 12656 15988 12665
rect 16212 12656 16264 12708
rect 20352 12792 20404 12844
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 23204 12792 23256 12844
rect 17776 12724 17828 12776
rect 20260 12724 20312 12776
rect 14832 12588 14884 12640
rect 20352 12656 20404 12708
rect 17224 12588 17276 12640
rect 17776 12588 17828 12640
rect 20076 12588 20128 12640
rect 21548 12588 21600 12640
rect 23756 12699 23808 12708
rect 23756 12665 23765 12699
rect 23765 12665 23799 12699
rect 23799 12665 23808 12699
rect 23756 12656 23808 12665
rect 23848 12699 23900 12708
rect 23848 12665 23857 12699
rect 23857 12665 23891 12699
rect 23891 12665 23900 12699
rect 23848 12656 23900 12665
rect 22928 12631 22980 12640
rect 22928 12597 22937 12631
rect 22937 12597 22971 12631
rect 22971 12597 22980 12631
rect 22928 12588 22980 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1952 12384 2004 12436
rect 2136 12384 2188 12436
rect 3148 12384 3200 12436
rect 3792 12427 3844 12436
rect 3792 12393 3801 12427
rect 3801 12393 3835 12427
rect 3835 12393 3844 12427
rect 3792 12384 3844 12393
rect 5080 12427 5132 12436
rect 5080 12393 5089 12427
rect 5089 12393 5123 12427
rect 5123 12393 5132 12427
rect 5080 12384 5132 12393
rect 7012 12384 7064 12436
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 11888 12384 11940 12436
rect 12440 12384 12492 12436
rect 14280 12384 14332 12436
rect 16304 12427 16356 12436
rect 16304 12393 16313 12427
rect 16313 12393 16347 12427
rect 16347 12393 16356 12427
rect 16304 12384 16356 12393
rect 19432 12384 19484 12436
rect 20996 12384 21048 12436
rect 21548 12427 21600 12436
rect 21548 12393 21557 12427
rect 21557 12393 21591 12427
rect 21591 12393 21600 12427
rect 21548 12384 21600 12393
rect 22928 12384 22980 12436
rect 23848 12384 23900 12436
rect 2228 12316 2280 12368
rect 2596 12316 2648 12368
rect 4160 12316 4212 12368
rect 4344 12316 4396 12368
rect 6000 12316 6052 12368
rect 9496 12316 9548 12368
rect 13912 12316 13964 12368
rect 14556 12316 14608 12368
rect 15568 12316 15620 12368
rect 16028 12359 16080 12368
rect 16028 12325 16037 12359
rect 16037 12325 16071 12359
rect 16071 12325 16080 12359
rect 16028 12316 16080 12325
rect 18788 12316 18840 12368
rect 21088 12316 21140 12368
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 16948 12291 17000 12300
rect 16948 12257 16957 12291
rect 16957 12257 16991 12291
rect 16991 12257 17000 12291
rect 16948 12248 17000 12257
rect 18420 12248 18472 12300
rect 20352 12248 20404 12300
rect 23204 12248 23256 12300
rect 25044 12316 25096 12368
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 5448 12180 5500 12232
rect 6552 12180 6604 12232
rect 8392 12180 8444 12232
rect 11612 12223 11664 12232
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 13820 12180 13872 12232
rect 15752 12180 15804 12232
rect 16856 12223 16908 12232
rect 16856 12189 16865 12223
rect 16865 12189 16899 12223
rect 16899 12189 16908 12223
rect 16856 12180 16908 12189
rect 17040 12180 17092 12232
rect 24216 12223 24268 12232
rect 24216 12189 24225 12223
rect 24225 12189 24259 12223
rect 24259 12189 24268 12223
rect 24216 12180 24268 12189
rect 3056 12112 3108 12164
rect 3332 12112 3384 12164
rect 4528 12112 4580 12164
rect 17776 12112 17828 12164
rect 18972 12112 19024 12164
rect 20996 12112 21048 12164
rect 2044 12044 2096 12096
rect 2780 12044 2832 12096
rect 8760 12044 8812 12096
rect 10508 12087 10560 12096
rect 10508 12053 10517 12087
rect 10517 12053 10551 12087
rect 10551 12053 10560 12087
rect 10508 12044 10560 12053
rect 11060 12087 11112 12096
rect 11060 12053 11069 12087
rect 11069 12053 11103 12087
rect 11103 12053 11112 12087
rect 11060 12044 11112 12053
rect 12532 12044 12584 12096
rect 12900 12087 12952 12096
rect 12900 12053 12909 12087
rect 12909 12053 12943 12087
rect 12943 12053 12952 12087
rect 12900 12044 12952 12053
rect 13636 12044 13688 12096
rect 14740 12087 14792 12096
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 15384 12044 15436 12096
rect 19156 12044 19208 12096
rect 20260 12087 20312 12096
rect 20260 12053 20269 12087
rect 20269 12053 20303 12087
rect 20303 12053 20312 12087
rect 20260 12044 20312 12053
rect 22652 12087 22704 12096
rect 22652 12053 22661 12087
rect 22661 12053 22695 12087
rect 22695 12053 22704 12087
rect 22652 12044 22704 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2228 11840 2280 11892
rect 2596 11815 2648 11824
rect 2596 11781 2605 11815
rect 2605 11781 2639 11815
rect 2639 11781 2648 11815
rect 2596 11772 2648 11781
rect 3884 11840 3936 11892
rect 5448 11883 5500 11892
rect 5448 11849 5457 11883
rect 5457 11849 5491 11883
rect 5491 11849 5500 11883
rect 5448 11840 5500 11849
rect 9220 11840 9272 11892
rect 9404 11883 9456 11892
rect 9404 11849 9413 11883
rect 9413 11849 9447 11883
rect 9447 11849 9456 11883
rect 9404 11840 9456 11849
rect 9496 11840 9548 11892
rect 10508 11840 10560 11892
rect 10968 11840 11020 11892
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 13268 11840 13320 11892
rect 14832 11840 14884 11892
rect 15568 11840 15620 11892
rect 18420 11840 18472 11892
rect 21088 11840 21140 11892
rect 21548 11840 21600 11892
rect 23848 11840 23900 11892
rect 24216 11840 24268 11892
rect 24860 11840 24912 11892
rect 8024 11772 8076 11824
rect 1860 11568 1912 11620
rect 6644 11704 6696 11756
rect 7012 11704 7064 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 4252 11679 4304 11688
rect 4252 11645 4261 11679
rect 4261 11645 4295 11679
rect 4295 11645 4304 11679
rect 4252 11636 4304 11645
rect 4804 11636 4856 11688
rect 7564 11679 7616 11688
rect 7564 11645 7573 11679
rect 7573 11645 7607 11679
rect 7607 11645 7616 11679
rect 7564 11636 7616 11645
rect 15384 11772 15436 11824
rect 13912 11704 13964 11756
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 1952 11500 2004 11552
rect 4344 11568 4396 11620
rect 6000 11568 6052 11620
rect 8668 11568 8720 11620
rect 3056 11543 3108 11552
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3056 11500 3108 11509
rect 6184 11500 6236 11552
rect 6552 11500 6604 11552
rect 10048 11500 10100 11552
rect 10968 11611 11020 11620
rect 10968 11577 10977 11611
rect 10977 11577 11011 11611
rect 11011 11577 11020 11611
rect 10968 11568 11020 11577
rect 11244 11568 11296 11620
rect 11888 11568 11940 11620
rect 13728 11568 13780 11620
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 16948 11772 17000 11824
rect 17132 11815 17184 11824
rect 17132 11781 17141 11815
rect 17141 11781 17175 11815
rect 17175 11781 17184 11815
rect 17132 11772 17184 11781
rect 19984 11772 20036 11824
rect 17040 11704 17092 11756
rect 18880 11747 18932 11756
rect 18880 11713 18889 11747
rect 18889 11713 18923 11747
rect 18923 11713 18932 11747
rect 18880 11704 18932 11713
rect 17224 11636 17276 11688
rect 16856 11568 16908 11620
rect 20076 11704 20128 11756
rect 21824 11679 21876 11688
rect 21824 11645 21833 11679
rect 21833 11645 21867 11679
rect 21867 11645 21876 11679
rect 21824 11636 21876 11645
rect 23940 11772 23992 11824
rect 24216 11704 24268 11756
rect 25044 11704 25096 11756
rect 23572 11636 23624 11688
rect 21548 11568 21600 11620
rect 17500 11543 17552 11552
rect 17500 11509 17509 11543
rect 17509 11509 17543 11543
rect 17543 11509 17552 11543
rect 17500 11500 17552 11509
rect 18788 11543 18840 11552
rect 18788 11509 18797 11543
rect 18797 11509 18831 11543
rect 18831 11509 18840 11543
rect 18788 11500 18840 11509
rect 20444 11543 20496 11552
rect 20444 11509 20453 11543
rect 20453 11509 20487 11543
rect 20487 11509 20496 11543
rect 20444 11500 20496 11509
rect 20996 11500 21048 11552
rect 25136 11500 25188 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 4252 11296 4304 11348
rect 7012 11339 7064 11348
rect 7012 11305 7021 11339
rect 7021 11305 7055 11339
rect 7055 11305 7064 11339
rect 7012 11296 7064 11305
rect 8392 11296 8444 11348
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 11612 11339 11664 11348
rect 10140 11296 10192 11305
rect 1768 11228 1820 11280
rect 2228 11271 2280 11280
rect 2228 11237 2237 11271
rect 2237 11237 2271 11271
rect 2271 11237 2280 11271
rect 2228 11228 2280 11237
rect 2964 11228 3016 11280
rect 4344 11271 4396 11280
rect 4344 11237 4353 11271
rect 4353 11237 4387 11271
rect 4387 11237 4396 11271
rect 4344 11228 4396 11237
rect 6184 11228 6236 11280
rect 8760 11271 8812 11280
rect 8760 11237 8769 11271
rect 8769 11237 8803 11271
rect 8803 11237 8812 11271
rect 8760 11228 8812 11237
rect 11612 11305 11621 11339
rect 11621 11305 11655 11339
rect 11655 11305 11664 11339
rect 11612 11296 11664 11305
rect 13820 11296 13872 11348
rect 19984 11339 20036 11348
rect 19984 11305 19993 11339
rect 19993 11305 20027 11339
rect 20027 11305 20036 11339
rect 19984 11296 20036 11305
rect 20260 11296 20312 11348
rect 24400 11296 24452 11348
rect 11152 11228 11204 11280
rect 13728 11271 13780 11280
rect 13728 11237 13731 11271
rect 13731 11237 13765 11271
rect 13765 11237 13780 11271
rect 13728 11228 13780 11237
rect 4252 11160 4304 11212
rect 4620 11160 4672 11212
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 8300 11203 8352 11212
rect 8300 11169 8309 11203
rect 8309 11169 8343 11203
rect 8343 11169 8352 11203
rect 8300 11160 8352 11169
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 8760 10956 8812 11008
rect 11336 11092 11388 11144
rect 12624 11160 12676 11212
rect 14740 11228 14792 11280
rect 16948 11228 17000 11280
rect 18788 11228 18840 11280
rect 17776 11203 17828 11212
rect 17776 11169 17785 11203
rect 17785 11169 17819 11203
rect 17819 11169 17828 11203
rect 17776 11160 17828 11169
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 21824 11228 21876 11280
rect 23204 11271 23256 11280
rect 23204 11237 23213 11271
rect 23213 11237 23247 11271
rect 23247 11237 23256 11271
rect 23204 11228 23256 11237
rect 20996 11203 21048 11212
rect 20996 11169 21005 11203
rect 21005 11169 21039 11203
rect 21039 11169 21048 11203
rect 20996 11160 21048 11169
rect 21272 11160 21324 11212
rect 24768 11160 24820 11212
rect 13820 11092 13872 11144
rect 15752 11135 15804 11144
rect 11888 11024 11940 11076
rect 15292 11024 15344 11076
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 19064 11135 19116 11144
rect 19064 11101 19073 11135
rect 19073 11101 19107 11135
rect 19107 11101 19116 11135
rect 19064 11092 19116 11101
rect 20352 11092 20404 11144
rect 23112 11135 23164 11144
rect 23112 11101 23121 11135
rect 23121 11101 23155 11135
rect 23155 11101 23164 11135
rect 23112 11092 23164 11101
rect 25136 11092 25188 11144
rect 22652 11024 22704 11076
rect 24032 11024 24084 11076
rect 12716 10956 12768 11008
rect 16396 10999 16448 11008
rect 16396 10965 16405 10999
rect 16405 10965 16439 10999
rect 16439 10965 16448 10999
rect 16396 10956 16448 10965
rect 18788 10956 18840 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1768 10795 1820 10804
rect 1768 10761 1777 10795
rect 1777 10761 1811 10795
rect 1811 10761 1820 10795
rect 1768 10752 1820 10761
rect 1952 10752 2004 10804
rect 2504 10752 2556 10804
rect 4252 10795 4304 10804
rect 4252 10761 4261 10795
rect 4261 10761 4295 10795
rect 4295 10761 4304 10795
rect 4252 10752 4304 10761
rect 5264 10752 5316 10804
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 8300 10752 8352 10804
rect 10140 10752 10192 10804
rect 12624 10795 12676 10804
rect 12624 10761 12633 10795
rect 12633 10761 12667 10795
rect 12667 10761 12676 10795
rect 12624 10752 12676 10761
rect 13728 10795 13780 10804
rect 13728 10761 13737 10795
rect 13737 10761 13771 10795
rect 13771 10761 13780 10795
rect 13728 10752 13780 10761
rect 15660 10752 15712 10804
rect 17776 10752 17828 10804
rect 23112 10752 23164 10804
rect 23572 10752 23624 10804
rect 25412 10795 25464 10804
rect 25412 10761 25421 10795
rect 25421 10761 25455 10795
rect 25455 10761 25464 10795
rect 25412 10752 25464 10761
rect 2964 10659 3016 10668
rect 2964 10625 2973 10659
rect 2973 10625 3007 10659
rect 3007 10625 3016 10659
rect 2964 10616 3016 10625
rect 4620 10548 4672 10600
rect 11060 10684 11112 10736
rect 15384 10684 15436 10736
rect 16948 10684 17000 10736
rect 19064 10684 19116 10736
rect 22192 10684 22244 10736
rect 5448 10616 5500 10668
rect 6460 10616 6512 10668
rect 8576 10616 8628 10668
rect 20444 10616 20496 10668
rect 21364 10616 21416 10668
rect 23204 10616 23256 10668
rect 24032 10659 24084 10668
rect 24032 10625 24041 10659
rect 24041 10625 24075 10659
rect 24075 10625 24084 10659
rect 24032 10616 24084 10625
rect 4988 10591 5040 10600
rect 4988 10557 4997 10591
rect 4997 10557 5031 10591
rect 5031 10557 5040 10591
rect 4988 10548 5040 10557
rect 2228 10412 2280 10464
rect 2504 10480 2556 10532
rect 8208 10548 8260 10600
rect 9128 10548 9180 10600
rect 10784 10548 10836 10600
rect 12716 10548 12768 10600
rect 9864 10480 9916 10532
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 8668 10412 8720 10464
rect 11244 10480 11296 10532
rect 11336 10480 11388 10532
rect 12900 10523 12952 10532
rect 12900 10489 12909 10523
rect 12909 10489 12943 10523
rect 12943 10489 12952 10523
rect 12900 10480 12952 10489
rect 15476 10548 15528 10600
rect 10876 10412 10928 10464
rect 14188 10412 14240 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 18880 10548 18932 10600
rect 19340 10480 19392 10532
rect 20168 10480 20220 10532
rect 17224 10412 17276 10464
rect 18788 10455 18840 10464
rect 18788 10421 18797 10455
rect 18797 10421 18831 10455
rect 18831 10421 18840 10455
rect 18788 10412 18840 10421
rect 19248 10412 19300 10464
rect 21272 10480 21324 10532
rect 21916 10523 21968 10532
rect 20996 10455 21048 10464
rect 20996 10421 21005 10455
rect 21005 10421 21039 10455
rect 21039 10421 21048 10455
rect 20996 10412 21048 10421
rect 21088 10412 21140 10464
rect 21916 10489 21925 10523
rect 21925 10489 21959 10523
rect 21959 10489 21968 10523
rect 21916 10480 21968 10489
rect 23756 10523 23808 10532
rect 23756 10489 23765 10523
rect 23765 10489 23799 10523
rect 23799 10489 23808 10523
rect 23756 10480 23808 10489
rect 23572 10412 23624 10464
rect 24032 10480 24084 10532
rect 24768 10455 24820 10464
rect 24768 10421 24777 10455
rect 24777 10421 24811 10455
rect 24811 10421 24820 10455
rect 24768 10412 24820 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1860 10208 1912 10260
rect 2320 10208 2372 10260
rect 4436 10251 4488 10260
rect 4436 10217 4445 10251
rect 4445 10217 4479 10251
rect 4479 10217 4488 10251
rect 4436 10208 4488 10217
rect 6092 10208 6144 10260
rect 10784 10251 10836 10260
rect 10784 10217 10793 10251
rect 10793 10217 10827 10251
rect 10827 10217 10836 10251
rect 10784 10208 10836 10217
rect 13636 10208 13688 10260
rect 15292 10208 15344 10260
rect 8208 10183 8260 10192
rect 8208 10149 8217 10183
rect 8217 10149 8251 10183
rect 8251 10149 8260 10183
rect 8208 10140 8260 10149
rect 1308 10072 1360 10124
rect 3332 10072 3384 10124
rect 3976 10072 4028 10124
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 5172 10072 5224 10124
rect 6276 10072 6328 10124
rect 6460 10115 6512 10124
rect 6460 10081 6469 10115
rect 6469 10081 6503 10115
rect 6503 10081 6512 10115
rect 6460 10072 6512 10081
rect 10140 10072 10192 10124
rect 10692 10115 10744 10124
rect 10692 10081 10701 10115
rect 10701 10081 10735 10115
rect 10735 10081 10744 10115
rect 10692 10072 10744 10081
rect 10876 10072 10928 10124
rect 11612 10115 11664 10124
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 12716 10072 12768 10124
rect 14188 10140 14240 10192
rect 16856 10140 16908 10192
rect 18788 10140 18840 10192
rect 21180 10183 21232 10192
rect 21180 10149 21189 10183
rect 21189 10149 21223 10183
rect 21223 10149 21232 10183
rect 21180 10140 21232 10149
rect 21916 10208 21968 10260
rect 22192 10208 22244 10260
rect 23756 10251 23808 10260
rect 23756 10217 23765 10251
rect 23765 10217 23799 10251
rect 23799 10217 23808 10251
rect 23756 10208 23808 10217
rect 24124 10208 24176 10260
rect 25228 10208 25280 10260
rect 22376 10140 22428 10192
rect 15384 10115 15436 10124
rect 7932 10004 7984 10056
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 15476 10072 15528 10124
rect 19248 10115 19300 10124
rect 19248 10081 19257 10115
rect 19257 10081 19291 10115
rect 19291 10081 19300 10115
rect 19248 10072 19300 10081
rect 19340 10072 19392 10124
rect 20996 10072 21048 10124
rect 22928 10115 22980 10124
rect 22928 10081 22937 10115
rect 22937 10081 22971 10115
rect 22971 10081 22980 10115
rect 22928 10072 22980 10081
rect 23112 10115 23164 10124
rect 23112 10081 23121 10115
rect 23121 10081 23155 10115
rect 23155 10081 23164 10115
rect 23112 10072 23164 10081
rect 24032 10072 24084 10124
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 19984 10047 20036 10056
rect 19984 10013 19993 10047
rect 19993 10013 20027 10047
rect 20027 10013 20036 10047
rect 19984 10004 20036 10013
rect 20720 10004 20772 10056
rect 8760 9936 8812 9988
rect 17224 9936 17276 9988
rect 17960 9936 18012 9988
rect 22284 9936 22336 9988
rect 24124 10004 24176 10056
rect 25320 10072 25372 10124
rect 2228 9911 2280 9920
rect 2228 9877 2237 9911
rect 2237 9877 2271 9911
rect 2271 9877 2280 9911
rect 2228 9868 2280 9877
rect 2872 9911 2924 9920
rect 2872 9877 2881 9911
rect 2881 9877 2915 9911
rect 2915 9877 2924 9911
rect 2872 9868 2924 9877
rect 9220 9868 9272 9920
rect 9496 9911 9548 9920
rect 9496 9877 9505 9911
rect 9505 9877 9539 9911
rect 9539 9877 9548 9911
rect 9496 9868 9548 9877
rect 12716 9911 12768 9920
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 14740 9868 14792 9920
rect 15844 9868 15896 9920
rect 17868 9911 17920 9920
rect 17868 9877 17877 9911
rect 17877 9877 17911 9911
rect 17911 9877 17920 9911
rect 17868 9868 17920 9877
rect 18880 9868 18932 9920
rect 21364 9868 21416 9920
rect 21824 9911 21876 9920
rect 21824 9877 21833 9911
rect 21833 9877 21867 9911
rect 21867 9877 21876 9911
rect 21824 9868 21876 9877
rect 23388 9868 23440 9920
rect 23756 9868 23808 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1308 9664 1360 9716
rect 3332 9707 3384 9716
rect 3332 9673 3341 9707
rect 3341 9673 3375 9707
rect 3375 9673 3384 9707
rect 3332 9664 3384 9673
rect 3976 9707 4028 9716
rect 3976 9673 3985 9707
rect 3985 9673 4019 9707
rect 4019 9673 4028 9707
rect 3976 9664 4028 9673
rect 5172 9664 5224 9716
rect 5540 9664 5592 9716
rect 6184 9664 6236 9716
rect 8208 9664 8260 9716
rect 9128 9707 9180 9716
rect 9128 9673 9137 9707
rect 9137 9673 9171 9707
rect 9171 9673 9180 9707
rect 9128 9664 9180 9673
rect 9772 9707 9824 9716
rect 9772 9673 9781 9707
rect 9781 9673 9815 9707
rect 9815 9673 9824 9707
rect 9772 9664 9824 9673
rect 10140 9664 10192 9716
rect 13820 9707 13872 9716
rect 13820 9673 13829 9707
rect 13829 9673 13863 9707
rect 13863 9673 13872 9707
rect 15384 9707 15436 9716
rect 13820 9664 13872 9673
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 17868 9664 17920 9716
rect 18512 9664 18564 9716
rect 19248 9664 19300 9716
rect 21088 9707 21140 9716
rect 21088 9673 21097 9707
rect 21097 9673 21131 9707
rect 21131 9673 21140 9707
rect 21088 9664 21140 9673
rect 112 9596 164 9648
rect 2136 9596 2188 9648
rect 2872 9596 2924 9648
rect 3148 9596 3200 9648
rect 3056 9528 3108 9580
rect 2044 9460 2096 9512
rect 1584 9392 1636 9444
rect 7656 9596 7708 9648
rect 10048 9528 10100 9580
rect 9220 9460 9272 9512
rect 9496 9460 9548 9512
rect 11336 9528 11388 9580
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 11704 9528 11756 9580
rect 14464 9596 14516 9648
rect 15844 9596 15896 9648
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 16212 9528 16264 9580
rect 16948 9528 17000 9580
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 12716 9503 12768 9512
rect 6460 9392 6512 9444
rect 8668 9392 8720 9444
rect 9128 9324 9180 9376
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 10692 9324 10744 9333
rect 11612 9324 11664 9376
rect 12256 9367 12308 9376
rect 12256 9333 12265 9367
rect 12265 9333 12299 9367
rect 12299 9333 12308 9367
rect 12256 9324 12308 9333
rect 14280 9460 14332 9512
rect 14464 9460 14516 9512
rect 15568 9460 15620 9512
rect 15844 9503 15896 9512
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 15844 9460 15896 9469
rect 15936 9460 15988 9512
rect 21916 9596 21968 9648
rect 18604 9571 18656 9580
rect 18604 9537 18613 9571
rect 18613 9537 18647 9571
rect 18647 9537 18656 9571
rect 18604 9528 18656 9537
rect 18788 9528 18840 9580
rect 20168 9571 20220 9580
rect 20168 9537 20177 9571
rect 20177 9537 20211 9571
rect 20211 9537 20220 9571
rect 20168 9528 20220 9537
rect 22928 9664 22980 9716
rect 24124 9707 24176 9716
rect 24124 9673 24133 9707
rect 24133 9673 24167 9707
rect 24167 9673 24176 9707
rect 24124 9664 24176 9673
rect 24676 9664 24728 9716
rect 24860 9707 24912 9716
rect 24860 9673 24869 9707
rect 24869 9673 24903 9707
rect 24903 9673 24912 9707
rect 24860 9664 24912 9673
rect 22376 9596 22428 9648
rect 23848 9596 23900 9648
rect 25320 9639 25372 9648
rect 25320 9605 25329 9639
rect 25329 9605 25363 9639
rect 25363 9605 25372 9639
rect 25320 9596 25372 9605
rect 27620 9596 27672 9648
rect 22284 9571 22336 9580
rect 22284 9537 22293 9571
rect 22293 9537 22327 9571
rect 22327 9537 22336 9571
rect 22284 9528 22336 9537
rect 23296 9528 23348 9580
rect 18880 9460 18932 9512
rect 14372 9324 14424 9376
rect 14740 9324 14792 9376
rect 18144 9435 18196 9444
rect 18144 9401 18153 9435
rect 18153 9401 18187 9435
rect 18187 9401 18196 9435
rect 18144 9392 18196 9401
rect 15844 9324 15896 9376
rect 16856 9324 16908 9376
rect 17868 9324 17920 9376
rect 19248 9367 19300 9376
rect 19248 9333 19257 9367
rect 19257 9333 19291 9367
rect 19291 9333 19300 9367
rect 19248 9324 19300 9333
rect 20720 9392 20772 9444
rect 20996 9324 21048 9376
rect 21180 9324 21232 9376
rect 22100 9435 22152 9444
rect 22100 9401 22109 9435
rect 22109 9401 22143 9435
rect 22143 9401 22152 9435
rect 22100 9392 22152 9401
rect 23112 9324 23164 9376
rect 23664 9367 23716 9376
rect 23664 9333 23673 9367
rect 23673 9333 23707 9367
rect 23707 9333 23716 9367
rect 23664 9324 23716 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 7932 9163 7984 9172
rect 7932 9129 7941 9163
rect 7941 9129 7975 9163
rect 7975 9129 7984 9163
rect 7932 9120 7984 9129
rect 9220 9120 9272 9172
rect 14464 9163 14516 9172
rect 14464 9129 14473 9163
rect 14473 9129 14507 9163
rect 14507 9129 14516 9163
rect 14464 9120 14516 9129
rect 15476 9120 15528 9172
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 20168 9163 20220 9172
rect 20168 9129 20177 9163
rect 20177 9129 20211 9163
rect 20211 9129 20220 9163
rect 20168 9120 20220 9129
rect 22100 9163 22152 9172
rect 22100 9129 22109 9163
rect 22109 9129 22143 9163
rect 22143 9129 22152 9163
rect 22100 9120 22152 9129
rect 23388 9120 23440 9172
rect 6368 9052 6420 9104
rect 6552 9095 6604 9104
rect 6552 9061 6561 9095
rect 6561 9061 6595 9095
rect 6595 9061 6604 9095
rect 6552 9052 6604 9061
rect 8300 9052 8352 9104
rect 8760 9095 8812 9104
rect 8760 9061 8769 9095
rect 8769 9061 8803 9095
rect 8803 9061 8812 9095
rect 8760 9052 8812 9061
rect 8944 9052 8996 9104
rect 10876 9052 10928 9104
rect 112 8984 164 9036
rect 1584 8984 1636 9036
rect 6000 9027 6052 9036
rect 6000 8993 6009 9027
rect 6009 8993 6043 9027
rect 6043 8993 6052 9027
rect 6000 8984 6052 8993
rect 6460 8984 6512 9036
rect 10508 8984 10560 9036
rect 10600 8984 10652 9036
rect 12440 9052 12492 9104
rect 12716 9052 12768 9104
rect 20720 9052 20772 9104
rect 20996 9052 21048 9104
rect 21364 9052 21416 9104
rect 8024 8848 8076 8900
rect 6736 8780 6788 8832
rect 11704 8916 11756 8968
rect 12808 8984 12860 9036
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 17224 8984 17276 9036
rect 17776 9027 17828 9036
rect 17776 8993 17785 9027
rect 17785 8993 17819 9027
rect 17819 8993 17828 9027
rect 17776 8984 17828 8993
rect 19156 9027 19208 9036
rect 19156 8993 19165 9027
rect 19165 8993 19199 9027
rect 19199 8993 19208 9027
rect 19156 8984 19208 8993
rect 19248 8984 19300 9036
rect 19984 8984 20036 9036
rect 22652 9027 22704 9036
rect 22652 8993 22661 9027
rect 22661 8993 22695 9027
rect 22695 8993 22704 9027
rect 22652 8984 22704 8993
rect 23848 8984 23900 9036
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 12256 8848 12308 8900
rect 14280 8848 14332 8900
rect 10692 8780 10744 8832
rect 13268 8823 13320 8832
rect 13268 8789 13277 8823
rect 13277 8789 13311 8823
rect 13311 8789 13320 8823
rect 13268 8780 13320 8789
rect 14372 8780 14424 8832
rect 16212 8780 16264 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2228 8576 2280 8628
rect 2780 8576 2832 8628
rect 6000 8576 6052 8628
rect 6460 8576 6512 8628
rect 6828 8576 6880 8628
rect 8300 8576 8352 8628
rect 8944 8619 8996 8628
rect 8944 8585 8953 8619
rect 8953 8585 8987 8619
rect 8987 8585 8996 8619
rect 8944 8576 8996 8585
rect 9312 8619 9364 8628
rect 9312 8585 9321 8619
rect 9321 8585 9355 8619
rect 9355 8585 9364 8619
rect 9312 8576 9364 8585
rect 9956 8576 10008 8628
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 12256 8576 12308 8628
rect 12716 8619 12768 8628
rect 12716 8585 12725 8619
rect 12725 8585 12759 8619
rect 12759 8585 12768 8619
rect 12716 8576 12768 8585
rect 12808 8576 12860 8628
rect 14372 8576 14424 8628
rect 15844 8576 15896 8628
rect 17776 8576 17828 8628
rect 19156 8576 19208 8628
rect 19984 8619 20036 8628
rect 19984 8585 19993 8619
rect 19993 8585 20027 8619
rect 20027 8585 20036 8619
rect 19984 8576 20036 8585
rect 10048 8508 10100 8560
rect 14832 8551 14884 8560
rect 14832 8517 14841 8551
rect 14841 8517 14875 8551
rect 14875 8517 14884 8551
rect 14832 8508 14884 8517
rect 15384 8508 15436 8560
rect 19248 8551 19300 8560
rect 19248 8517 19257 8551
rect 19257 8517 19291 8551
rect 19291 8517 19300 8551
rect 19248 8508 19300 8517
rect 1400 8372 1452 8424
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 2688 8372 2740 8424
rect 7840 8440 7892 8492
rect 9588 8440 9640 8492
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 13176 8440 13228 8492
rect 16120 8440 16172 8492
rect 16856 8440 16908 8492
rect 18052 8483 18104 8492
rect 10692 8372 10744 8424
rect 9036 8304 9088 8356
rect 10508 8304 10560 8356
rect 12440 8347 12492 8356
rect 12440 8313 12449 8347
rect 12449 8313 12483 8347
rect 12483 8313 12492 8347
rect 12440 8304 12492 8313
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 14372 8372 14424 8424
rect 14924 8372 14976 8424
rect 15660 8372 15712 8424
rect 16212 8372 16264 8424
rect 16488 8372 16540 8424
rect 18052 8449 18061 8483
rect 18061 8449 18095 8483
rect 18095 8449 18104 8483
rect 18052 8440 18104 8449
rect 19340 8372 19392 8424
rect 20812 8576 20864 8628
rect 20996 8619 21048 8628
rect 20996 8585 21005 8619
rect 21005 8585 21039 8619
rect 21039 8585 21048 8619
rect 20996 8576 21048 8585
rect 21824 8576 21876 8628
rect 23848 8619 23900 8628
rect 23848 8585 23857 8619
rect 23857 8585 23891 8619
rect 23891 8585 23900 8619
rect 23848 8576 23900 8585
rect 21916 8483 21968 8492
rect 21916 8449 21925 8483
rect 21925 8449 21959 8483
rect 21959 8449 21968 8483
rect 21916 8440 21968 8449
rect 9680 8279 9732 8288
rect 9680 8245 9689 8279
rect 9689 8245 9723 8279
rect 9723 8245 9732 8279
rect 9680 8236 9732 8245
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 12164 8279 12216 8288
rect 10048 8236 10100 8245
rect 12164 8245 12173 8279
rect 12173 8245 12207 8279
rect 12207 8245 12216 8279
rect 12164 8236 12216 8245
rect 12624 8236 12676 8288
rect 12992 8236 13044 8288
rect 13636 8236 13688 8288
rect 14556 8279 14608 8288
rect 14556 8245 14565 8279
rect 14565 8245 14599 8279
rect 14599 8245 14608 8279
rect 14556 8236 14608 8245
rect 15292 8236 15344 8288
rect 15660 8236 15712 8288
rect 16304 8236 16356 8288
rect 21732 8304 21784 8356
rect 18972 8279 19024 8288
rect 18972 8245 18981 8279
rect 18981 8245 19015 8279
rect 19015 8245 19024 8279
rect 18972 8236 19024 8245
rect 20536 8236 20588 8288
rect 22652 8279 22704 8288
rect 22652 8245 22661 8279
rect 22661 8245 22695 8279
rect 22695 8245 22704 8279
rect 22652 8236 22704 8245
rect 27712 8236 27764 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 8944 8032 8996 8084
rect 9036 8075 9088 8084
rect 9036 8041 9045 8075
rect 9045 8041 9079 8075
rect 9079 8041 9088 8075
rect 9036 8032 9088 8041
rect 9404 8032 9456 8084
rect 4160 7964 4212 8016
rect 8024 8007 8076 8016
rect 8024 7973 8033 8007
rect 8033 7973 8067 8007
rect 8067 7973 8076 8007
rect 8024 7964 8076 7973
rect 9864 8032 9916 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 12900 8032 12952 8084
rect 14832 8075 14884 8084
rect 14832 8041 14841 8075
rect 14841 8041 14875 8075
rect 14875 8041 14884 8075
rect 14832 8032 14884 8041
rect 17500 8032 17552 8084
rect 19156 8032 19208 8084
rect 19524 8032 19576 8084
rect 20536 8032 20588 8084
rect 17868 7964 17920 8016
rect 18972 7964 19024 8016
rect 20996 7964 21048 8016
rect 2412 7939 2464 7948
rect 112 7760 164 7812
rect 2412 7905 2421 7939
rect 2421 7905 2455 7939
rect 2455 7905 2464 7939
rect 2412 7896 2464 7905
rect 1860 7760 1912 7812
rect 8668 7760 8720 7812
rect 10692 7896 10744 7948
rect 11244 7896 11296 7948
rect 9588 7828 9640 7880
rect 12164 7896 12216 7948
rect 14832 7896 14884 7948
rect 14924 7896 14976 7948
rect 15476 7896 15528 7948
rect 15660 7896 15712 7948
rect 16028 7896 16080 7948
rect 17316 7896 17368 7948
rect 18788 7896 18840 7948
rect 15752 7871 15804 7880
rect 11520 7760 11572 7812
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 18604 7871 18656 7880
rect 16120 7760 16172 7812
rect 8576 7692 8628 7744
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 10048 7735 10100 7744
rect 10048 7701 10057 7735
rect 10057 7701 10091 7735
rect 10091 7701 10100 7735
rect 10048 7692 10100 7701
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 17224 7692 17276 7744
rect 17408 7692 17460 7744
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 20352 7828 20404 7880
rect 18236 7692 18288 7744
rect 21824 7735 21876 7744
rect 21824 7701 21833 7735
rect 21833 7701 21867 7735
rect 21867 7701 21876 7735
rect 21824 7692 21876 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1676 7488 1728 7540
rect 1860 7531 1912 7540
rect 1860 7497 1869 7531
rect 1869 7497 1903 7531
rect 1903 7497 1912 7531
rect 1860 7488 1912 7497
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 9588 7488 9640 7540
rect 11704 7488 11756 7540
rect 16120 7531 16172 7540
rect 16120 7497 16129 7531
rect 16129 7497 16163 7531
rect 16163 7497 16172 7531
rect 16120 7488 16172 7497
rect 17316 7488 17368 7540
rect 17868 7531 17920 7540
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 17868 7488 17920 7497
rect 19064 7531 19116 7540
rect 19064 7497 19073 7531
rect 19073 7497 19107 7531
rect 19107 7497 19116 7531
rect 19064 7488 19116 7497
rect 19248 7488 19300 7540
rect 20996 7531 21048 7540
rect 9496 7420 9548 7472
rect 1216 7352 1268 7404
rect 11060 7420 11112 7472
rect 14832 7463 14884 7472
rect 14832 7429 14841 7463
rect 14841 7429 14875 7463
rect 14875 7429 14884 7463
rect 14832 7420 14884 7429
rect 11244 7352 11296 7404
rect 11520 7352 11572 7404
rect 13636 7352 13688 7404
rect 17500 7352 17552 7404
rect 18236 7352 18288 7404
rect 18788 7395 18840 7404
rect 18788 7361 18797 7395
rect 18797 7361 18831 7395
rect 18831 7361 18840 7395
rect 18788 7352 18840 7361
rect 20996 7497 21005 7531
rect 21005 7497 21039 7531
rect 21039 7497 21048 7531
rect 20996 7488 21048 7497
rect 25964 7488 26016 7540
rect 21916 7395 21968 7404
rect 10048 7327 10100 7336
rect 10048 7293 10057 7327
rect 10057 7293 10091 7327
rect 10091 7293 10100 7327
rect 10048 7284 10100 7293
rect 12900 7284 12952 7336
rect 14740 7327 14792 7336
rect 10692 7216 10744 7268
rect 12440 7216 12492 7268
rect 13176 7216 13228 7268
rect 14740 7293 14749 7327
rect 14749 7293 14783 7327
rect 14783 7293 14792 7327
rect 14740 7284 14792 7293
rect 13820 7259 13872 7268
rect 13820 7225 13829 7259
rect 13829 7225 13863 7259
rect 13863 7225 13872 7259
rect 13820 7216 13872 7225
rect 2412 7148 2464 7200
rect 5540 7148 5592 7200
rect 7564 7148 7616 7200
rect 10048 7148 10100 7200
rect 11888 7148 11940 7200
rect 12164 7148 12216 7200
rect 14556 7191 14608 7200
rect 14556 7157 14565 7191
rect 14565 7157 14599 7191
rect 14599 7157 14608 7191
rect 15660 7284 15712 7336
rect 19064 7284 19116 7336
rect 21916 7361 21925 7395
rect 21925 7361 21959 7395
rect 21959 7361 21968 7395
rect 21916 7352 21968 7361
rect 15476 7259 15528 7268
rect 15476 7225 15485 7259
rect 15485 7225 15519 7259
rect 15519 7225 15528 7259
rect 15476 7216 15528 7225
rect 16488 7259 16540 7268
rect 16488 7225 16497 7259
rect 16497 7225 16531 7259
rect 16531 7225 16540 7259
rect 16488 7216 16540 7225
rect 16672 7216 16724 7268
rect 18236 7259 18288 7268
rect 18236 7225 18245 7259
rect 18245 7225 18279 7259
rect 18279 7225 18288 7259
rect 18236 7216 18288 7225
rect 14556 7148 14608 7157
rect 15384 7148 15436 7200
rect 20352 7259 20404 7268
rect 20352 7225 20361 7259
rect 20361 7225 20395 7259
rect 20395 7225 20404 7259
rect 20352 7216 20404 7225
rect 21824 7216 21876 7268
rect 22376 7191 22428 7200
rect 22376 7157 22385 7191
rect 22385 7157 22419 7191
rect 22419 7157 22428 7191
rect 22376 7148 22428 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1216 6944 1268 6996
rect 9404 6987 9456 6996
rect 9404 6953 9413 6987
rect 9413 6953 9447 6987
rect 9447 6953 9456 6987
rect 9404 6944 9456 6953
rect 14832 6987 14884 6996
rect 14832 6953 14841 6987
rect 14841 6953 14875 6987
rect 14875 6953 14884 6987
rect 14832 6944 14884 6953
rect 15384 6944 15436 6996
rect 15568 6944 15620 6996
rect 16488 6944 16540 6996
rect 21824 6944 21876 6996
rect 9680 6919 9732 6928
rect 9680 6885 9689 6919
rect 9689 6885 9723 6919
rect 9723 6885 9732 6919
rect 9680 6876 9732 6885
rect 10324 6851 10376 6860
rect 10324 6817 10333 6851
rect 10333 6817 10367 6851
rect 10367 6817 10376 6851
rect 10324 6808 10376 6817
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 14740 6876 14792 6928
rect 16212 6876 16264 6928
rect 16856 6876 16908 6928
rect 18328 6919 18380 6928
rect 18328 6885 18337 6919
rect 18337 6885 18371 6919
rect 18371 6885 18380 6919
rect 18328 6876 18380 6885
rect 20352 6876 20404 6928
rect 12992 6740 13044 6792
rect 14280 6851 14332 6860
rect 14280 6817 14289 6851
rect 14289 6817 14323 6851
rect 14323 6817 14332 6851
rect 14280 6808 14332 6817
rect 15476 6808 15528 6860
rect 19524 6808 19576 6860
rect 16580 6740 16632 6792
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 18788 6715 18840 6724
rect 10876 6647 10928 6656
rect 10876 6613 10885 6647
rect 10885 6613 10919 6647
rect 10919 6613 10928 6647
rect 10876 6604 10928 6613
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 18788 6681 18797 6715
rect 18797 6681 18831 6715
rect 18831 6681 18840 6715
rect 18788 6672 18840 6681
rect 18144 6604 18196 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 9404 6400 9456 6452
rect 10324 6443 10376 6452
rect 10324 6409 10333 6443
rect 10333 6409 10367 6443
rect 10367 6409 10376 6443
rect 10324 6400 10376 6409
rect 12164 6400 12216 6452
rect 12808 6400 12860 6452
rect 13268 6400 13320 6452
rect 10876 6375 10928 6384
rect 10876 6341 10885 6375
rect 10885 6341 10919 6375
rect 10919 6341 10928 6375
rect 10876 6332 10928 6341
rect 4804 6264 4856 6316
rect 11336 6332 11388 6384
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 9404 6171 9456 6180
rect 9404 6137 9413 6171
rect 9413 6137 9447 6171
rect 9447 6137 9456 6171
rect 9404 6128 9456 6137
rect 10692 6196 10744 6248
rect 11152 6196 11204 6248
rect 16672 6400 16724 6452
rect 16856 6443 16908 6452
rect 16856 6409 16865 6443
rect 16865 6409 16899 6443
rect 16899 6409 16908 6443
rect 16856 6400 16908 6409
rect 19524 6400 19576 6452
rect 14372 6264 14424 6316
rect 15568 6239 15620 6248
rect 12808 6128 12860 6180
rect 14004 6128 14056 6180
rect 15568 6205 15577 6239
rect 15577 6205 15611 6239
rect 15611 6205 15620 6239
rect 15568 6196 15620 6205
rect 18328 6264 18380 6316
rect 18144 6239 18196 6248
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 18144 6196 18196 6205
rect 10692 6103 10744 6112
rect 10692 6069 10701 6103
rect 10701 6069 10735 6103
rect 10735 6069 10744 6103
rect 10692 6060 10744 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 9404 5899 9456 5908
rect 9404 5865 9413 5899
rect 9413 5865 9447 5899
rect 9447 5865 9456 5899
rect 9404 5856 9456 5865
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 13452 5899 13504 5908
rect 13452 5865 13461 5899
rect 13461 5865 13495 5899
rect 13495 5865 13504 5899
rect 13452 5856 13504 5865
rect 14372 5899 14424 5908
rect 14372 5865 14381 5899
rect 14381 5865 14415 5899
rect 14415 5865 14424 5899
rect 14372 5856 14424 5865
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 15568 5856 15620 5908
rect 16580 5899 16632 5908
rect 16580 5865 16589 5899
rect 16589 5865 16623 5899
rect 16623 5865 16632 5899
rect 16580 5856 16632 5865
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 18236 5856 18288 5865
rect 10968 5788 11020 5840
rect 10692 5720 10744 5772
rect 12900 5788 12952 5840
rect 13268 5788 13320 5840
rect 16948 5831 17000 5840
rect 16948 5797 16957 5831
rect 16957 5797 16991 5831
rect 16991 5797 17000 5831
rect 16948 5788 17000 5797
rect 17500 5831 17552 5840
rect 17500 5797 17509 5831
rect 17509 5797 17543 5831
rect 17543 5797 17552 5831
rect 17500 5788 17552 5797
rect 11428 5763 11480 5772
rect 11428 5729 11437 5763
rect 11437 5729 11471 5763
rect 11471 5729 11480 5763
rect 11428 5720 11480 5729
rect 13544 5720 13596 5772
rect 15752 5763 15804 5772
rect 15752 5729 15761 5763
rect 15761 5729 15795 5763
rect 15795 5729 15804 5763
rect 15752 5720 15804 5729
rect 11520 5652 11572 5704
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 13176 5584 13228 5636
rect 16764 5584 16816 5636
rect 17224 5516 17276 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 10968 5312 11020 5364
rect 13268 5355 13320 5364
rect 13268 5321 13277 5355
rect 13277 5321 13311 5355
rect 13311 5321 13320 5355
rect 13268 5312 13320 5321
rect 13544 5355 13596 5364
rect 13544 5321 13553 5355
rect 13553 5321 13587 5355
rect 13587 5321 13596 5355
rect 13544 5312 13596 5321
rect 14004 5355 14056 5364
rect 14004 5321 14013 5355
rect 14013 5321 14047 5355
rect 14047 5321 14056 5355
rect 14004 5312 14056 5321
rect 15752 5312 15804 5364
rect 15844 5244 15896 5296
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 16948 5176 17000 5228
rect 9864 5151 9916 5160
rect 9864 5117 9873 5151
rect 9873 5117 9907 5151
rect 9907 5117 9916 5151
rect 9864 5108 9916 5117
rect 11428 5108 11480 5160
rect 13820 5108 13872 5160
rect 15292 5151 15344 5160
rect 15292 5117 15301 5151
rect 15301 5117 15335 5151
rect 15335 5117 15344 5151
rect 15292 5108 15344 5117
rect 16672 5151 16724 5160
rect 16672 5117 16681 5151
rect 16681 5117 16715 5151
rect 16715 5117 16724 5151
rect 16672 5108 16724 5117
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 18880 4972 18932 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 10968 4811 11020 4820
rect 10968 4777 10977 4811
rect 10977 4777 11011 4811
rect 11011 4777 11020 4811
rect 10968 4768 11020 4777
rect 16856 4768 16908 4820
rect 22376 4768 22428 4820
rect 10876 4675 10928 4684
rect 10876 4641 10885 4675
rect 10885 4641 10919 4675
rect 10919 4641 10928 4675
rect 10876 4632 10928 4641
rect 16580 4675 16632 4684
rect 16580 4641 16598 4675
rect 16598 4641 16632 4675
rect 16580 4632 16632 4641
rect 17684 4632 17736 4684
rect 21732 4675 21784 4684
rect 21732 4641 21741 4675
rect 21741 4641 21775 4675
rect 21775 4641 21784 4675
rect 21732 4632 21784 4641
rect 16672 4564 16724 4616
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 16580 4267 16632 4276
rect 16580 4233 16589 4267
rect 16589 4233 16623 4267
rect 16623 4233 16632 4267
rect 16580 4224 16632 4233
rect 21732 4224 21784 4276
rect 27620 4224 27672 4276
rect 10784 3927 10836 3936
rect 10784 3893 10793 3927
rect 10793 3893 10827 3927
rect 10827 3893 10836 3927
rect 10784 3884 10836 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 112 3544 164 3596
rect 1400 3587 1452 3596
rect 1400 3553 1444 3587
rect 1444 3553 1452 3587
rect 1400 3544 1452 3553
rect 11336 3476 11388 3528
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1400 3136 1452 3188
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 24124 2592 24176 2644
rect 25136 2456 25188 2508
rect 25136 2295 25188 2304
rect 25136 2261 25145 2295
rect 25145 2261 25179 2295
rect 25179 2261 25188 2295
rect 25136 2252 25188 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 19432 76 19484 128
rect 20076 76 20128 128
<< metal2 >>
rect 662 27520 718 28000
rect 2042 27520 2098 28000
rect 3422 27520 3478 28000
rect 4802 27532 4858 28000
rect 6182 27554 6238 28000
rect 4802 27520 4804 27532
rect 676 24614 704 27520
rect 1306 27160 1362 27169
rect 2056 27130 2084 27520
rect 1306 27095 1362 27104
rect 2044 27124 2096 27130
rect 664 24608 716 24614
rect 664 24550 716 24556
rect 1216 20936 1268 20942
rect 1216 20878 1268 20884
rect 110 20088 166 20097
rect 166 20058 244 20074
rect 166 20052 256 20058
rect 166 20046 204 20052
rect 110 20023 166 20032
rect 204 19994 256 20000
rect 204 19168 256 19174
rect 110 19136 166 19145
rect 166 19116 204 19122
rect 166 19110 256 19116
rect 166 19094 244 19110
rect 110 19071 166 19080
rect 1228 15337 1256 20878
rect 1320 20602 1348 27095
rect 2044 27066 2096 27072
rect 1490 25800 1546 25809
rect 1490 25735 1546 25744
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1412 23866 1440 24210
rect 1400 23860 1452 23866
rect 1400 23802 1452 23808
rect 1504 23798 1532 25735
rect 3436 25158 3464 27520
rect 4856 27520 4858 27532
rect 6104 27526 6238 27554
rect 4804 27474 4856 27480
rect 4816 27443 4844 27474
rect 6000 27124 6052 27130
rect 6000 27066 6052 27072
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 1582 24848 1638 24857
rect 1582 24783 1638 24792
rect 1596 24410 1624 24783
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1582 24032 1638 24041
rect 1582 23967 1638 23976
rect 1492 23792 1544 23798
rect 1492 23734 1544 23740
rect 1596 23322 1624 23967
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 2044 23860 2096 23866
rect 2044 23802 2096 23808
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1400 23180 1452 23186
rect 1400 23122 1452 23128
rect 1412 22438 1440 23122
rect 1490 22672 1546 22681
rect 1490 22607 1546 22616
rect 1400 22432 1452 22438
rect 1400 22374 1452 22380
rect 1504 21690 1532 22607
rect 2056 22098 2084 23802
rect 2964 23520 3016 23526
rect 2964 23462 3016 23468
rect 1952 22092 2004 22098
rect 1952 22034 2004 22040
rect 2044 22092 2096 22098
rect 2044 22034 2096 22040
rect 1768 21888 1820 21894
rect 1768 21830 1820 21836
rect 1582 21720 1638 21729
rect 1492 21684 1544 21690
rect 1582 21655 1638 21664
rect 1492 21626 1544 21632
rect 1596 21146 1624 21655
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1308 20596 1360 20602
rect 1308 20538 1360 20544
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1412 19224 1440 19858
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1492 19236 1544 19242
rect 1412 19196 1492 19224
rect 1214 15328 1270 15337
rect 1214 15263 1270 15272
rect 1306 12336 1362 12345
rect 1306 12271 1362 12280
rect 1214 10296 1270 10305
rect 1214 10231 1270 10240
rect 110 9752 166 9761
rect 110 9687 166 9696
rect 124 9654 152 9687
rect 112 9648 164 9654
rect 112 9590 164 9596
rect 112 9036 164 9042
rect 112 8978 164 8984
rect 124 8809 152 8978
rect 110 8800 166 8809
rect 110 8735 166 8744
rect 112 7812 164 7818
rect 112 7754 164 7760
rect 124 7721 152 7754
rect 110 7712 166 7721
rect 110 7647 166 7656
rect 1228 7410 1256 10231
rect 1320 10130 1348 12271
rect 1308 10124 1360 10130
rect 1308 10066 1360 10072
rect 1320 9722 1348 10066
rect 1308 9716 1360 9722
rect 1308 9658 1360 9664
rect 1412 8430 1440 19196
rect 1492 19178 1544 19184
rect 1688 18630 1716 19246
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1780 17864 1808 21830
rect 1964 21350 1992 22034
rect 1952 21344 2004 21350
rect 1952 21286 2004 21292
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 1860 18148 1912 18154
rect 1860 18090 1912 18096
rect 1504 17836 1808 17864
rect 1504 13734 1532 17836
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1596 9450 1624 16390
rect 1872 16250 1900 18090
rect 1964 17649 1992 21286
rect 2044 21004 2096 21010
rect 2044 20946 2096 20952
rect 2056 20262 2084 20946
rect 2136 20800 2188 20806
rect 2136 20742 2188 20748
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 2056 19310 2084 20198
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 2044 17808 2096 17814
rect 2044 17750 2096 17756
rect 1950 17640 2006 17649
rect 1950 17575 2006 17584
rect 2056 17338 2084 17750
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 2056 16998 2084 17274
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1872 15978 1900 16186
rect 2148 16114 2176 20742
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2424 20058 2452 20198
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2228 18896 2280 18902
rect 2228 18838 2280 18844
rect 2240 16726 2268 18838
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2228 16720 2280 16726
rect 2228 16662 2280 16668
rect 2240 16250 2268 16662
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2136 16108 2188 16114
rect 2056 16068 2136 16096
rect 1860 15972 1912 15978
rect 1860 15914 1912 15920
rect 2056 15706 2084 16068
rect 2136 16050 2188 16056
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 1858 15464 1914 15473
rect 1858 15399 1914 15408
rect 1872 14958 1900 15399
rect 2044 15088 2096 15094
rect 2044 15030 2096 15036
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1780 14074 1808 14486
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1584 9444 1636 9450
rect 1584 9386 1636 9392
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1596 8634 1624 8978
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1688 7546 1716 13738
rect 1964 12850 1992 14826
rect 2056 14550 2084 15030
rect 2044 14544 2096 14550
rect 2044 14486 2096 14492
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1964 12442 1992 12786
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 2056 12102 2084 14350
rect 2136 13796 2188 13802
rect 2136 13738 2188 13744
rect 2148 13530 2176 13738
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2148 12442 2176 13262
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2240 11898 2268 12310
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 1860 11620 1912 11626
rect 1860 11562 1912 11568
rect 1768 11280 1820 11286
rect 1768 11222 1820 11228
rect 1780 10810 1808 11222
rect 1872 11014 1900 11562
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1872 10266 1900 10950
rect 1964 10810 1992 11494
rect 2240 11286 2268 11834
rect 2228 11280 2280 11286
rect 2042 11248 2098 11257
rect 2228 11222 2280 11228
rect 2042 11183 2098 11192
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 2056 9518 2084 11183
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2148 9654 2176 11086
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2240 9926 2268 10406
rect 2332 10266 2360 18566
rect 2424 18290 2452 19110
rect 2516 18766 2544 21286
rect 2686 20632 2742 20641
rect 2686 20567 2742 20576
rect 2700 19786 2728 20567
rect 2976 20398 3004 23462
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 3056 22092 3108 22098
rect 3056 22034 3108 22040
rect 3068 21554 3096 22034
rect 3516 21956 3568 21962
rect 3516 21898 3568 21904
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 3068 21457 3096 21490
rect 3054 21448 3110 21457
rect 3054 21383 3110 21392
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 3344 20602 3372 20878
rect 3332 20596 3384 20602
rect 3332 20538 3384 20544
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 3148 20324 3200 20330
rect 3148 20266 3200 20272
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2688 19780 2740 19786
rect 2688 19722 2740 19728
rect 2792 19242 2820 19858
rect 2780 19236 2832 19242
rect 2780 19178 2832 19184
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2516 18426 2544 18702
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2424 17882 2452 18226
rect 2412 17876 2464 17882
rect 2412 17818 2464 17824
rect 2608 17610 2636 18702
rect 2596 17604 2648 17610
rect 2596 17546 2648 17552
rect 2608 16182 2636 17546
rect 2884 17202 2912 20198
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 3068 18290 3096 18702
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 3068 17202 3096 18226
rect 3160 17678 3188 20266
rect 3424 18896 3476 18902
rect 3424 18838 3476 18844
rect 3436 18358 3464 18838
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3436 17338 3464 17614
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 2884 16794 2912 17138
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 3068 16726 3096 17138
rect 3528 16794 3556 21898
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 4988 21412 5040 21418
rect 4988 21354 5040 21360
rect 3792 20460 3844 20466
rect 3792 20402 3844 20408
rect 3700 19168 3752 19174
rect 3700 19110 3752 19116
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 2596 16176 2648 16182
rect 2596 16118 2648 16124
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 3068 15706 3096 16050
rect 3528 15960 3556 16730
rect 3608 15972 3660 15978
rect 3528 15932 3608 15960
rect 3608 15914 3660 15920
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3436 15706 3464 15846
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 2504 15632 2556 15638
rect 2504 15574 2556 15580
rect 2688 15632 2740 15638
rect 2688 15574 2740 15580
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2424 14822 2452 15438
rect 2516 14822 2544 15574
rect 2700 15026 2728 15574
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 3344 15026 3372 15370
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 2412 14816 2464 14822
rect 2412 14758 2464 14764
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2240 8634 2268 9862
rect 2424 9178 2452 14758
rect 2516 13784 2544 14758
rect 2700 14550 2728 14962
rect 2964 14884 3016 14890
rect 2964 14826 3016 14832
rect 2976 14618 3004 14826
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2596 13796 2648 13802
rect 2516 13756 2596 13784
rect 2596 13738 2648 13744
rect 3436 13734 3464 15642
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3528 14618 3556 15438
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3528 13938 3556 14554
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3712 13814 3740 19110
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 3620 13786 3740 13814
rect 3804 13814 3832 20402
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 3884 19168 3936 19174
rect 3884 19110 3936 19116
rect 3896 18970 3924 19110
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 3988 18601 4016 20334
rect 5000 20058 5028 21354
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 4620 19916 4672 19922
rect 4620 19858 4672 19864
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 4632 19718 4660 19858
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 3974 18592 4030 18601
rect 3974 18527 4030 18536
rect 4172 18426 4200 18702
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 3976 18148 4028 18154
rect 3976 18090 4028 18096
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3896 17882 3924 18022
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3988 17610 4016 18090
rect 4080 17882 4108 18090
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 3976 17604 4028 17610
rect 3976 17546 4028 17552
rect 4172 16998 4200 17750
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16454 4200 16934
rect 4264 16794 4292 17070
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 3988 14346 4016 15574
rect 4068 14884 4120 14890
rect 4252 14884 4304 14890
rect 4120 14844 4252 14872
rect 4068 14826 4120 14832
rect 4252 14826 4304 14832
rect 4356 14482 4384 19110
rect 4632 18766 4660 19654
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4632 18154 4660 18702
rect 4620 18148 4672 18154
rect 4620 18090 4672 18096
rect 4632 17610 4660 18090
rect 4620 17604 4672 17610
rect 4620 17546 4672 17552
rect 4620 16652 4672 16658
rect 4724 16640 4752 19314
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4672 16612 4752 16640
rect 4620 16594 4672 16600
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 4448 14958 4476 15302
rect 4540 15162 4568 16390
rect 4632 16182 4660 16594
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4632 15910 4660 16118
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3804 13786 4016 13814
rect 3424 13728 3476 13734
rect 2686 13696 2742 13705
rect 3424 13670 3476 13676
rect 2686 13631 2742 13640
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2516 12918 2544 13398
rect 2504 12912 2556 12918
rect 2504 12854 2556 12860
rect 2596 12708 2648 12714
rect 2596 12650 2648 12656
rect 2608 12374 2636 12650
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 2608 12238 2636 12310
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2608 11830 2636 12174
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2516 10538 2544 10746
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2700 8430 2728 13631
rect 3528 13530 3556 13738
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2976 12850 3004 13262
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2792 8634 2820 12038
rect 2976 11286 3004 12786
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 3068 11558 3096 12106
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 2976 10674 3004 11222
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9654 2912 9862
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 3068 9586 3096 11494
rect 3160 9654 3188 12378
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3344 10130 3372 12106
rect 3620 11257 3648 13786
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3804 12442 3832 12786
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3896 11898 3924 12650
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3606 11248 3662 11257
rect 3606 11183 3662 11192
rect 3988 10962 4016 13786
rect 4080 12186 4108 14214
rect 4356 13530 4384 14418
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4172 12850 4200 13262
rect 4264 12986 4292 13398
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4172 12374 4200 12786
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4080 12158 4200 12186
rect 3988 10934 4108 10962
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 3344 9722 3372 10066
rect 3988 9722 4016 10066
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1872 7546 1900 7754
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 2332 7449 2360 8366
rect 4080 8129 4108 10934
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 4172 8022 4200 12158
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4264 11354 4292 11630
rect 4356 11626 4384 12310
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4356 11286 4384 11562
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4264 10810 4292 11154
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4448 10266 4476 14894
rect 4540 14822 4568 15098
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 14618 4568 14758
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4540 12714 4568 13262
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4540 12170 4568 12650
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4632 11218 4660 15846
rect 4816 11694 4844 19110
rect 5000 18970 5028 19178
rect 5368 19174 5396 19858
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 4988 18964 5040 18970
rect 5040 18924 5120 18952
rect 4988 18906 5040 18912
rect 4896 18896 4948 18902
rect 4896 18838 4948 18844
rect 4908 18358 4936 18838
rect 4896 18352 4948 18358
rect 4896 18294 4948 18300
rect 4908 17338 4936 18294
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 5000 16114 5028 16594
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5000 15638 5028 16050
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 5092 13784 5120 18924
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5184 15910 5212 17614
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5276 15570 5304 15982
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5276 15473 5304 15506
rect 5262 15464 5318 15473
rect 5262 15399 5318 15408
rect 5172 13796 5224 13802
rect 5092 13756 5172 13784
rect 5092 13530 5120 13756
rect 5172 13738 5224 13744
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5092 12442 5120 12922
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5000 10606 5028 11154
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4632 10130 4660 10542
rect 5184 10130 5212 13738
rect 5276 12986 5304 15399
rect 5368 15366 5396 19110
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18222 6040 27066
rect 6104 19922 6132 27526
rect 6182 27520 6238 27526
rect 6460 27532 6512 27538
rect 7654 27520 7710 28000
rect 7760 27526 8064 27554
rect 7760 27520 7788 27526
rect 7668 27492 7788 27520
rect 6460 27474 6512 27480
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6104 18834 6132 19858
rect 6288 18970 6316 24550
rect 6276 18964 6328 18970
rect 6276 18906 6328 18912
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6104 18426 6132 18770
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 6472 18358 6500 27474
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 6932 19378 6960 25094
rect 8036 19922 8064 27526
rect 9034 27520 9090 28000
rect 9680 27532 9732 27538
rect 9048 23474 9076 27520
rect 10414 27532 10470 28000
rect 10414 27520 10416 27532
rect 9680 27474 9732 27480
rect 10468 27520 10470 27532
rect 11440 27526 11744 27554
rect 10416 27474 10468 27480
rect 8956 23446 9076 23474
rect 8956 19922 8984 23446
rect 9034 22672 9090 22681
rect 9034 22607 9090 22616
rect 9048 22438 9076 22607
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 7668 19514 7696 19858
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7392 19281 7420 19314
rect 7378 19272 7434 19281
rect 7378 19207 7434 19216
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 6552 18896 6604 18902
rect 6552 18838 6604 18844
rect 6564 18630 6592 18838
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 6460 18352 6512 18358
rect 6274 18320 6330 18329
rect 6460 18294 6512 18300
rect 6274 18255 6330 18264
rect 6288 18222 6316 18255
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6012 17066 6040 17614
rect 6472 17202 6500 17818
rect 6564 17746 6592 18566
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6932 17882 6960 18090
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 7116 17814 7144 18022
rect 7104 17808 7156 17814
rect 7104 17750 7156 17756
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 7116 17338 7144 17750
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 6840 16726 6868 17070
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6092 16516 6144 16522
rect 6092 16458 6144 16464
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6104 16250 6132 16458
rect 6092 16244 6144 16250
rect 6012 16204 6092 16232
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5460 15094 5488 15574
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5460 14482 5488 15030
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5552 14278 5580 15438
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6012 14006 6040 16204
rect 6092 16186 6144 16192
rect 6932 15910 6960 17002
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7116 16046 7144 16594
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 6104 13938 6132 14350
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5276 10810 5304 12922
rect 5552 12646 5580 13262
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5460 11898 5488 12174
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5460 10674 5488 11834
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5184 9722 5212 10066
rect 5552 9722 5580 12582
rect 6012 12374 6040 13670
rect 6104 13530 6132 13874
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11626 6040 12310
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 11286 6224 11494
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6104 10266 6132 11086
rect 6196 10810 6224 11222
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6288 10130 6316 13942
rect 6380 13870 6408 15846
rect 7116 15638 7144 15982
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6460 14884 6512 14890
rect 6460 14826 6512 14832
rect 6472 14618 6500 14826
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6472 14489 6500 14554
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6380 13734 6408 13806
rect 6932 13734 6960 14894
rect 7208 14550 7236 19110
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7300 15638 7328 18566
rect 7576 18154 7604 18702
rect 7564 18148 7616 18154
rect 7564 18090 7616 18096
rect 7576 17678 7604 18090
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7576 16794 7604 17614
rect 7668 17202 7696 18906
rect 7944 18873 7972 19654
rect 8036 19514 8064 19858
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 7930 18864 7986 18873
rect 8036 18834 8064 19450
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 7930 18799 7986 18808
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 8036 18426 8064 18770
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 7852 17785 7880 18294
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7838 17776 7894 17785
rect 7838 17711 7894 17720
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7300 14618 7328 15574
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 13870 7328 14214
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7116 13734 7144 13806
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 6184 9716 6236 9722
rect 6288 9704 6316 10066
rect 6236 9676 6316 9704
rect 6184 9658 6236 9664
rect 6380 9110 6408 13670
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6656 12646 6684 13398
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6564 11558 6592 12174
rect 6656 11762 6684 12582
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6472 10130 6500 10610
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6472 9450 6500 10066
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6472 9042 6500 9386
rect 6564 9110 6592 11494
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8634 6040 8978
rect 6472 8634 6500 8978
rect 6748 8838 6776 12718
rect 6840 12646 6868 13126
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7024 12714 7052 12854
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6840 8634 6868 12582
rect 7024 12442 7052 12650
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7024 11354 7052 11698
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2318 7440 2374 7449
rect 1216 7404 1268 7410
rect 2318 7375 2374 7384
rect 1216 7346 1268 7352
rect 1228 7002 1256 7346
rect 2424 7206 2452 7890
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 7576 7206 7604 11630
rect 7668 9654 7696 17138
rect 7748 15632 7800 15638
rect 7748 15574 7800 15580
rect 7760 15162 7788 15574
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7760 14482 7788 14554
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 14074 7788 14418
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7852 8498 7880 17711
rect 7944 17066 7972 18022
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 8036 16250 8064 16594
rect 8024 16244 8076 16250
rect 8024 16186 8076 16192
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7944 13530 7972 14486
rect 8036 14074 8064 16186
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7944 12442 7972 13262
rect 8036 12646 8064 13466
rect 8128 13326 8156 19110
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8312 18222 8340 18634
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8220 17270 8248 17750
rect 8208 17264 8260 17270
rect 8208 17206 8260 17212
rect 8312 16794 8340 18158
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8312 16046 8340 16594
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8312 15706 8340 15982
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 14414 8248 15438
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8298 13968 8354 13977
rect 8404 13954 8432 15846
rect 8354 13926 8432 13954
rect 8298 13903 8354 13912
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 8036 11830 8064 12582
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 8312 11218 8340 13903
rect 8392 13320 8444 13326
rect 8496 13297 8524 19654
rect 8956 19514 8984 19858
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 8956 19310 8984 19450
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8588 13870 8616 15302
rect 8864 15026 8892 15846
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8864 14618 8892 14962
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8576 13864 8628 13870
rect 8852 13864 8904 13870
rect 8628 13824 8852 13852
rect 8576 13806 8628 13812
rect 8852 13806 8904 13812
rect 8392 13262 8444 13268
rect 8482 13288 8538 13297
rect 8404 12782 8432 13262
rect 8482 13223 8538 13232
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8404 12238 8432 12718
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11354 8432 12174
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8588 11218 8616 12922
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8772 12102 8800 12718
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8312 10810 8340 11154
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8588 10674 8616 11154
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8220 10198 8248 10542
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7944 9178 7972 9998
rect 8220 9722 8248 10134
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 8312 9110 8340 10406
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 8036 8022 8064 8842
rect 8312 8634 8340 9046
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8298 8120 8354 8129
rect 8298 8055 8354 8064
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 8312 7313 8340 8055
rect 8588 7750 8616 10610
rect 8680 10470 8708 11562
rect 8772 11286 8800 12038
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8680 9450 8708 10406
rect 8772 9994 8800 10950
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8772 9110 8800 9930
rect 9048 9602 9076 22374
rect 9692 20466 9720 27474
rect 10428 27443 10456 27474
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 11152 23180 11204 23186
rect 11152 23122 11204 23128
rect 11164 22438 11192 23122
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9232 11898 9260 13262
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9140 9722 9168 10542
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9048 9574 9168 9602
rect 9140 9382 9168 9574
rect 9232 9518 9260 9862
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8956 8634 8984 9046
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9048 8090 9076 8298
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8956 7857 8984 8026
rect 8942 7848 8998 7857
rect 8668 7812 8720 7818
rect 8942 7783 8998 7792
rect 8668 7754 8720 7760
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8680 7546 8708 7754
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8298 7304 8354 7313
rect 8298 7239 8354 7248
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 1216 6996 1268 7002
rect 1216 6938 1268 6944
rect 110 6896 166 6905
rect 110 6831 166 6840
rect 124 5681 152 6831
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 110 5672 166 5681
rect 110 5607 166 5616
rect 1766 5264 1822 5273
rect 1766 5199 1822 5208
rect 112 3596 164 3602
rect 112 3538 164 3544
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 124 3505 152 3538
rect 110 3496 166 3505
rect 110 3431 166 3440
rect 1412 3194 1440 3538
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1490 82 1546 480
rect 1780 82 1808 5199
rect 1490 54 1808 82
rect 4526 82 4582 480
rect 4816 82 4844 6258
rect 5552 1465 5580 7142
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 9140 6361 9168 9318
rect 9232 9178 9260 9454
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9324 8634 9352 19110
rect 9692 18834 9720 20402
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9692 18426 9720 18770
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9784 18034 9812 19110
rect 9692 18006 9812 18034
rect 9692 16046 9720 18006
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9784 17134 9812 17818
rect 9876 17746 9904 20198
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9876 17338 9904 17682
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9784 16794 9812 17070
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9876 16658 9904 17274
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9692 15706 9720 15982
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9784 15094 9812 15438
rect 9876 15162 9904 15574
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 9876 14550 9904 14826
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 13938 9720 14350
rect 9876 14074 9904 14486
rect 9864 14068 9916 14074
rect 9784 14028 9864 14056
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9416 11898 9444 13466
rect 9784 12714 9812 14028
rect 9864 14010 9916 14016
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9876 13394 9904 13738
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9876 12918 9904 13330
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9508 12374 9536 12582
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9508 11898 9536 12310
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9518 9536 9862
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9416 7002 9444 8026
rect 9600 7886 9628 8434
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7478 9536 7686
rect 9600 7546 9628 7822
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9416 6458 9444 6938
rect 9692 6934 9720 8230
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9126 6352 9182 6361
rect 9126 6287 9182 6296
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9416 5914 9444 6122
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 7562 5672 7618 5681
rect 7562 5607 7618 5616
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5538 1456 5594 1465
rect 5538 1391 5594 1400
rect 4526 54 4844 82
rect 7576 82 7604 5607
rect 9784 4154 9812 9658
rect 9876 8090 9904 10474
rect 9968 8634 9996 20198
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10048 17808 10100 17814
rect 10048 17750 10100 17756
rect 10060 16998 10088 17750
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10060 16658 10088 16934
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 10152 16522 10180 19654
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10336 18290 10364 18566
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10704 17678 10732 18226
rect 10888 17882 10916 18566
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10888 17202 10916 17818
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 10244 16114 10272 16594
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15570 10732 16118
rect 10796 15910 10824 16594
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10876 15020 10928 15026
rect 10980 15008 11008 19654
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 11072 16590 11100 17546
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11072 16046 11100 16526
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11072 15638 11100 15846
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 11072 15366 11100 15574
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10928 14980 11008 15008
rect 10876 14962 10928 14968
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14618 10732 14758
rect 10888 14618 10916 14962
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10980 13870 11008 14282
rect 11072 14278 11100 15302
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 13870 11100 14214
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10152 12986 10180 13330
rect 11072 13190 11100 13806
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 11072 12782 11100 13126
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 9586 10088 11494
rect 10152 11354 10180 12242
rect 11072 12102 11100 12718
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10520 11898 10548 12038
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10980 11626 11008 11834
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10152 10810 10180 11290
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 11072 10742 11100 12038
rect 11164 11762 11192 22374
rect 11440 19922 11468 27526
rect 11716 27520 11744 27526
rect 11794 27520 11850 28000
rect 13174 27554 13230 28000
rect 14646 27554 14702 28000
rect 13004 27526 13230 27554
rect 11716 27492 11836 27520
rect 13004 23866 13032 27526
rect 13174 27520 13230 27526
rect 13636 27532 13688 27538
rect 13636 27474 13688 27480
rect 14568 27526 14702 27554
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 13004 23662 13032 23802
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 11440 19310 11468 19858
rect 11428 19304 11480 19310
rect 11428 19246 11480 19252
rect 12360 18970 12388 23462
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11256 16794 11284 17614
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11348 17066 11376 17478
rect 11336 17060 11388 17066
rect 11336 17002 11388 17008
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11532 16794 11560 17002
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11256 16182 11284 16730
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11256 15026 11284 15506
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11624 13814 11652 18158
rect 11716 18086 11744 18770
rect 12176 18222 12204 18770
rect 12360 18290 12388 18906
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11532 13786 11652 13814
rect 11440 13326 11468 13738
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11348 12322 11376 13194
rect 11440 12442 11468 13262
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11348 12294 11468 12322
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11164 11286 11192 11698
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11060 10736 11112 10742
rect 10138 10704 10194 10713
rect 11060 10678 11112 10684
rect 10138 10639 10194 10648
rect 10152 10130 10180 10639
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10796 10266 10824 10542
rect 11256 10538 11284 11562
rect 11334 11248 11390 11257
rect 11334 11183 11390 11192
rect 11348 11150 11376 11183
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11244 10532 11296 10538
rect 11244 10474 11296 10480
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10888 10130 10916 10406
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10152 9722 10180 10066
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10704 9382 10732 10066
rect 10888 9518 10916 10066
rect 11348 9586 11376 10474
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10600 9036 10652 9042
rect 10704 9024 10732 9318
rect 10888 9110 10916 9454
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10652 8996 10732 9024
rect 10600 8978 10652 8984
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 10060 8294 10088 8502
rect 10520 8362 10548 8978
rect 10612 8498 10640 8978
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10704 8430 10732 8774
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 10060 7750 10088 8230
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 7954 10732 8366
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 7342 10088 7686
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10704 7274 10732 7890
rect 11256 7750 11284 7890
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 9862 5264 9918 5273
rect 9862 5199 9918 5208
rect 9876 5166 9904 5199
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9784 4126 9904 4154
rect 9876 2689 9904 4126
rect 9862 2680 9918 2689
rect 9862 2615 9918 2624
rect 10060 1329 10088 7142
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10336 6458 10364 6802
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10704 6254 10732 7210
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10888 6390 10916 6598
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10704 6118 10732 6190
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5778 10732 6054
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10888 4690 10916 6326
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 10980 5370 11008 5782
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10980 4826 11008 5306
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10888 4154 10916 4626
rect 10796 4126 10916 4154
rect 10796 3942 10824 4126
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10796 3641 10824 3878
rect 10782 3632 10838 3641
rect 10782 3567 10838 3576
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10046 1320 10102 1329
rect 10046 1255 10102 1264
rect 7654 82 7710 480
rect 7576 54 7710 82
rect 1490 0 1546 54
rect 4526 0 4582 54
rect 7654 0 7710 54
rect 10782 82 10838 480
rect 11072 82 11100 7414
rect 11256 7410 11284 7686
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11256 6322 11284 7346
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11348 6390 11376 6802
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11152 6248 11204 6254
rect 11440 6236 11468 12294
rect 11532 9586 11560 13786
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11624 12238 11652 12650
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11624 11354 11652 12174
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11716 11064 11744 18022
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11900 17066 11928 17750
rect 12544 17542 12572 18090
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12636 17134 12664 17478
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 11900 16658 11928 17002
rect 11992 16726 12020 17070
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11808 15502 11836 16526
rect 11900 16250 11928 16594
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11900 15162 11928 16186
rect 12728 16114 12756 16730
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12728 15858 12756 16050
rect 12820 15978 12848 16390
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12728 15830 12848 15858
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11900 14550 11928 15098
rect 12728 14958 12756 15302
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 11900 13462 11928 14486
rect 12176 14074 12204 14486
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12176 13734 12204 14010
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12176 13530 12204 13670
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11900 12986 11928 13398
rect 12360 13394 12388 14350
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12544 13258 12572 13738
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11900 12442 11928 12922
rect 12728 12850 12756 14350
rect 12820 13938 12848 15830
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12912 15026 12940 15302
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 13004 13258 13032 19110
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13188 17338 13216 17750
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 13096 15162 13124 15574
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13096 14618 13124 15098
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13280 14346 13308 18158
rect 13360 18148 13412 18154
rect 13360 18090 13412 18096
rect 13372 17678 13400 18090
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13372 16454 13400 17614
rect 13464 17270 13492 19110
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 14414 13400 16390
rect 13464 15978 13492 16934
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13464 15638 13492 15914
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13268 14340 13320 14346
rect 13268 14282 13320 14288
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12442 12480 12582
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 11900 11898 11928 12378
rect 12544 12102 12572 12650
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11900 11626 11928 11834
rect 12912 11665 12940 12038
rect 13280 11898 13308 14282
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 12898 11656 12954 11665
rect 11888 11620 11940 11626
rect 12898 11591 12954 11600
rect 11888 11562 11940 11568
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 11888 11076 11940 11082
rect 11716 11036 11888 11064
rect 11888 11018 11940 11024
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11624 9382 11652 10066
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11716 8974 11744 9522
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11532 7410 11560 7754
rect 11716 7546 11744 8570
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11900 7206 11928 11018
rect 12636 10810 12664 11154
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 8906 12296 9318
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12268 8634 12296 8842
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12452 8362 12480 9046
rect 12636 8514 12664 10746
rect 12728 10606 12756 10950
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 10130 12756 10542
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12728 9926 12756 10066
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12728 9518 12756 9862
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 9110 12756 9454
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12728 8634 12756 9046
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12820 8634 12848 8978
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12636 8486 12756 8514
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 7954 12204 8230
rect 12452 8090 12480 8298
rect 12636 8294 12664 8366
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12176 7206 12204 7890
rect 12452 7274 12480 8026
rect 12440 7268 12492 7274
rect 12440 7210 12492 7216
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 6458 12204 7142
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 11152 6190 11204 6196
rect 11348 6208 11468 6236
rect 11164 5234 11192 6190
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11348 3534 11376 6208
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11440 5166 11468 5714
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11532 5030 11560 5646
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11532 2825 11560 4966
rect 12728 2961 12756 8486
rect 12820 6458 12848 8570
rect 12912 8090 12940 10474
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13004 8294 13032 8978
rect 13188 8498 13216 8978
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12912 7342 12940 8026
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12820 6186 12848 6394
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12912 5846 12940 7278
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13004 5914 13032 6734
rect 13188 6662 13216 7210
rect 13280 6866 13308 8774
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 13188 5642 13216 6598
rect 13280 6458 13308 6802
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13280 5846 13308 6394
rect 13464 5914 13492 14826
rect 13556 12850 13584 23462
rect 13648 19514 13676 27474
rect 14568 23866 14596 27526
rect 14646 27520 14702 27526
rect 16026 27532 16082 28000
rect 16026 27520 16028 27532
rect 16080 27520 16082 27532
rect 17406 27520 17462 28000
rect 18786 27520 18842 28000
rect 20166 27520 20222 28000
rect 21638 27520 21694 28000
rect 23018 27520 23074 28000
rect 24398 27554 24454 28000
rect 24136 27526 24454 27554
rect 16028 27474 16080 27480
rect 16040 27443 16068 27474
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 17420 23866 17448 27520
rect 18800 24410 18828 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 17604 23866 17632 24210
rect 14556 23860 14608 23866
rect 14556 23802 14608 23808
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 14568 23662 14596 23802
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16408 23322 16436 23598
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 15120 23089 15148 23258
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15106 23080 15162 23089
rect 15106 23015 15162 23024
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22438 15332 23122
rect 17604 22681 17632 23802
rect 20180 23798 20208 27520
rect 21652 23866 21680 27520
rect 23032 23866 23060 27520
rect 24032 24744 24084 24750
rect 24032 24686 24084 24692
rect 23480 24268 23532 24274
rect 23480 24210 23532 24216
rect 23492 23866 23520 24210
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 23020 23860 23072 23866
rect 23020 23802 23072 23808
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 17590 22672 17646 22681
rect 17590 22607 17646 22616
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13740 19310 13768 19722
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13740 16998 13768 17614
rect 13832 17610 13860 18770
rect 13924 17660 13952 22374
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 19260 21457 19288 23598
rect 19246 21448 19302 21457
rect 19246 21383 19302 21392
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 14016 19174 14044 19858
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14016 17785 14044 19110
rect 14002 17776 14058 17785
rect 14002 17711 14058 17720
rect 13924 17632 14136 17660
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13924 15910 13952 16594
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13832 15162 13860 15438
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13648 14618 13676 14894
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13832 13870 13860 14418
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13740 12986 13768 13330
rect 13924 13308 13952 15846
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 14016 14006 14044 14418
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 14004 13320 14056 13326
rect 13924 13280 14004 13308
rect 14004 13262 14056 13268
rect 14016 12986 14044 13262
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14108 12918 14136 17632
rect 14200 13814 14228 19654
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14372 19304 14424 19310
rect 14648 19304 14700 19310
rect 14372 19246 14424 19252
rect 14568 19264 14648 19292
rect 14384 18222 14412 19246
rect 14568 18834 14596 19264
rect 14648 19246 14700 19252
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14568 18630 14596 18770
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14476 18222 14504 18566
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 17882 14504 18158
rect 14568 18154 14596 18566
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14476 16658 14504 17818
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 15502 14320 16526
rect 14476 16250 14504 16594
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14568 15910 14596 18090
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14200 13786 14320 13814
rect 14292 13734 14320 13786
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14384 13462 14412 15438
rect 14568 14822 14596 15846
rect 14844 15026 14872 18702
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14936 15706 14964 15982
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14936 15434 14964 15642
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14292 12442 14320 12650
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 13912 12368 13964 12374
rect 13912 12310 13964 12316
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11694 13676 12038
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13648 10266 13676 11630
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13740 11286 13768 11562
rect 13832 11354 13860 12174
rect 13924 11762 13952 12310
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13740 10810 13768 11222
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13832 9722 13860 11086
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10198 14228 10406
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 14200 9586 14228 10134
rect 14476 9654 14504 13806
rect 14568 13802 14596 14758
rect 15304 14482 15332 19178
rect 15580 19174 15608 19858
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15580 18329 15608 19110
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15566 18320 15622 18329
rect 15566 18255 15622 18264
rect 15672 18222 15700 18566
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15396 17202 15424 17614
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15396 16794 15424 17138
rect 15488 17134 15516 18090
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15580 17814 15608 18022
rect 15568 17808 15620 17814
rect 15568 17750 15620 17756
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15488 16794 15516 17070
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15476 16652 15528 16658
rect 15580 16640 15608 17478
rect 15672 16726 15700 18158
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15528 16612 15608 16640
rect 15476 16594 15528 16600
rect 15488 15910 15516 16594
rect 15764 16114 15792 19450
rect 16224 19242 16252 19654
rect 16212 19236 16264 19242
rect 16212 19178 16264 19184
rect 16224 18873 16252 19178
rect 16316 18902 16344 20198
rect 19260 19990 19288 21383
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16948 19236 17000 19242
rect 16948 19178 17000 19184
rect 17040 19236 17092 19242
rect 17040 19178 17092 19184
rect 16304 18896 16356 18902
rect 16210 18864 16266 18873
rect 16304 18838 16356 18844
rect 16396 18896 16448 18902
rect 16396 18838 16448 18844
rect 16210 18799 16266 18808
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15856 16658 15884 18226
rect 16316 17882 16344 18838
rect 16408 18426 16436 18838
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16500 17338 16528 19178
rect 16960 18902 16988 19178
rect 16948 18896 17000 18902
rect 16948 18838 17000 18844
rect 17052 18290 17080 19178
rect 17512 19174 17540 19246
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17236 17746 17264 18022
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15580 15094 15608 15914
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14740 14000 14792 14006
rect 14738 13968 14740 13977
rect 14792 13968 14794 13977
rect 14738 13903 14794 13912
rect 14752 13870 14780 13903
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14556 13796 14608 13802
rect 14556 13738 14608 13744
rect 14568 13394 14596 13738
rect 14752 13530 14780 13806
rect 15304 13530 15332 14418
rect 15764 13814 15792 16050
rect 15856 15706 15884 16594
rect 16500 16114 16528 16730
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15948 14521 15976 15846
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16132 14890 16160 15642
rect 16120 14884 16172 14890
rect 16120 14826 16172 14832
rect 16132 14550 16160 14826
rect 16592 14822 16620 15914
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16684 14550 16712 15302
rect 16120 14544 16172 14550
rect 15934 14512 15990 14521
rect 16120 14486 16172 14492
rect 16672 14544 16724 14550
rect 16672 14486 16724 14492
rect 15934 14447 15990 14456
rect 16132 14074 16160 14486
rect 17052 14414 17080 16458
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17236 15162 17264 15438
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 15672 13786 15792 13814
rect 16500 13802 16528 14214
rect 16868 13938 16896 14214
rect 17052 14074 17080 14350
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16396 13796 16448 13802
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14568 12374 14596 12786
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14752 12102 14780 12650
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11286 14780 12038
rect 14844 11898 14872 12582
rect 15580 12374 15608 13126
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 15396 11830 15424 12038
rect 15580 11898 15608 12310
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10266 15332 11018
rect 15672 10810 15700 13786
rect 16396 13738 16448 13744
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16408 13530 16436 13738
rect 17420 13734 17448 14486
rect 17512 14006 17540 19110
rect 17880 18902 17908 19722
rect 18064 19514 18092 19858
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 18616 19310 18644 19858
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 18052 18896 18104 18902
rect 18052 18838 18104 18844
rect 17880 18426 17908 18838
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 17696 17066 17724 17818
rect 17972 17270 18000 18362
rect 18064 18086 18092 18838
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18064 17542 18092 18022
rect 18156 17746 18184 19110
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18432 18290 18460 18906
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18524 17882 18552 18090
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18144 17740 18196 17746
rect 18144 17682 18196 17688
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18156 17338 18184 17682
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 18800 17202 18828 19790
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19260 19310 19288 19722
rect 19444 19378 19472 19858
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19248 19304 19300 19310
rect 19444 19281 19472 19314
rect 19248 19246 19300 19252
rect 19430 19272 19486 19281
rect 18972 19236 19024 19242
rect 18972 19178 19024 19184
rect 18984 17882 19012 19178
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19076 18970 19104 19110
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 18788 17196 18840 17202
rect 18788 17138 18840 17144
rect 17684 17060 17736 17066
rect 17684 17002 17736 17008
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 17788 16794 17816 16934
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17604 15978 17632 16390
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17604 14414 17632 15914
rect 17788 15910 17816 16594
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17788 15473 17816 15846
rect 17868 15496 17920 15502
rect 17774 15464 17830 15473
rect 17868 15438 17920 15444
rect 17774 15399 17830 15408
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17696 14550 17724 14758
rect 17684 14544 17736 14550
rect 17684 14486 17736 14492
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17500 14000 17552 14006
rect 17500 13942 17552 13948
rect 17604 13938 17632 14350
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15948 12714 15976 13330
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 16040 12374 16068 12854
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16028 12368 16080 12374
rect 16028 12310 16080 12316
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 11762 15792 12174
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15764 11150 15792 11698
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15384 10736 15436 10742
rect 16224 10713 16252 12650
rect 16316 12442 16344 12786
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16868 11626 16896 12174
rect 16960 11830 16988 12242
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16960 11286 16988 11766
rect 17052 11762 17080 12174
rect 17144 11830 17172 12922
rect 17236 12646 17264 13262
rect 17788 12986 17816 15399
rect 17880 14278 17908 15438
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17788 12782 17816 12922
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17776 12640 17828 12646
rect 17880 12628 17908 13330
rect 17828 12600 17908 12628
rect 17776 12582 17828 12588
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17236 11694 17264 12582
rect 17788 12170 17816 12582
rect 17776 12164 17828 12170
rect 17776 12106 17828 12112
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16408 10713 16436 10950
rect 16960 10742 16988 11222
rect 16948 10736 17000 10742
rect 15384 10678 15436 10684
rect 16210 10704 16266 10713
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15396 10130 15424 10678
rect 16210 10639 16266 10648
rect 16394 10704 16450 10713
rect 16948 10678 17000 10684
rect 16394 10639 16450 10648
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15488 10130 15516 10542
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14292 8906 14320 9454
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13648 7410 13676 8230
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13280 5370 13308 5782
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13556 5370 13584 5714
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 12714 2952 12770 2961
rect 12714 2887 12770 2896
rect 11518 2816 11574 2825
rect 11518 2751 11574 2760
rect 10782 54 11100 82
rect 13648 82 13676 7346
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13832 5166 13860 7210
rect 14292 6866 14320 8842
rect 14384 8838 14412 9318
rect 14476 9178 14504 9454
rect 14752 9382 14780 9862
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15396 9722 15424 10066
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14384 8634 14412 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14384 8430 14412 8570
rect 15396 8566 15424 9658
rect 15488 9178 15516 10066
rect 15580 9518 15608 10406
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15856 9654 15884 9862
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15856 9518 15884 9590
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15844 9376 15896 9382
rect 15948 9364 15976 9454
rect 15896 9336 15976 9364
rect 15844 9318 15896 9324
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 15384 8560 15436 8566
rect 15384 8502 15436 8508
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7206 14596 8230
rect 14844 8090 14872 8502
rect 15672 8430 15700 8978
rect 15856 8634 15884 9318
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14844 7954 14872 8026
rect 14936 7954 14964 8366
rect 15672 8294 15700 8366
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 14844 7478 14872 7890
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14280 6860 14332 6866
rect 14332 6820 14412 6848
rect 14280 6802 14332 6808
rect 14384 6322 14412 6820
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 14016 5370 14044 6122
rect 14384 5914 14412 6258
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14568 5681 14596 7142
rect 14752 6934 14780 7278
rect 14844 7002 14872 7414
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14554 5672 14610 5681
rect 14554 5607 14610 5616
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 15304 5166 15332 8230
rect 15672 7954 15700 8230
rect 15476 7948 15528 7954
rect 15660 7948 15712 7954
rect 15528 7908 15608 7936
rect 15476 7890 15528 7896
rect 15476 7268 15528 7274
rect 15476 7210 15528 7216
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 7002 15424 7142
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15488 6866 15516 7210
rect 15580 7002 15608 7908
rect 15660 7890 15712 7896
rect 15672 7342 15700 7890
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15488 5914 15516 6802
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15580 5914 15608 6190
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15764 5778 15792 7822
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15764 5370 15792 5714
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15856 5302 15884 8570
rect 16040 7954 16068 9998
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16224 8838 16252 9522
rect 16868 9382 16896 10134
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16960 9586 16988 9998
rect 17236 9994 17264 10406
rect 17224 9988 17276 9994
rect 17224 9930 17276 9936
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16132 7818 16160 8434
rect 16224 8430 16252 8774
rect 16868 8498 16896 9318
rect 16960 9178 16988 9522
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 17236 9042 17264 9930
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16212 8424 16264 8430
rect 16488 8424 16540 8430
rect 16212 8366 16264 8372
rect 16316 8384 16488 8412
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 16132 7546 16160 7754
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16224 6934 16252 8366
rect 16316 8294 16344 8384
rect 16488 8366 16540 8372
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16684 7274 16712 7686
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16500 7002 16528 7210
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16592 5914 16620 6734
rect 16684 6458 16712 7210
rect 16868 6934 16896 8434
rect 17236 7750 17264 8978
rect 17512 8090 17540 11494
rect 17788 11218 17816 12106
rect 17972 11336 18000 16050
rect 18248 15706 18276 16390
rect 18616 16182 18644 16594
rect 19076 16454 19104 16934
rect 19260 16726 19288 19246
rect 19430 19207 19486 19216
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19444 17066 19472 17818
rect 19432 17060 19484 17066
rect 19432 17002 19484 17008
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 18604 16176 18656 16182
rect 18604 16118 18656 16124
rect 18696 15972 18748 15978
rect 18696 15914 18748 15920
rect 19248 15972 19300 15978
rect 19248 15914 19300 15920
rect 18708 15706 18736 15914
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 17880 11308 18000 11336
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17788 10810 17816 11154
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17880 10010 17908 11308
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17696 9982 17908 10010
rect 17972 9994 18000 11154
rect 17960 9988 18012 9994
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16868 6458 16896 6870
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 16684 5166 16712 6394
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 16592 4282 16620 4626
rect 16684 4622 16712 5102
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 13910 82 13966 480
rect 13648 54 13966 82
rect 16776 82 16804 5578
rect 16868 4826 16896 5646
rect 16960 5234 16988 5782
rect 17236 5574 17264 7686
rect 17328 7546 17356 7890
rect 17406 7848 17462 7857
rect 17406 7783 17462 7792
rect 17420 7750 17448 7783
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17512 5846 17540 7346
rect 17500 5840 17552 5846
rect 17696 5817 17724 9982
rect 17960 9930 18012 9936
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 9722 17908 9862
rect 17868 9716 17920 9722
rect 18064 9674 18092 15506
rect 18248 15026 18276 15642
rect 19260 15434 19288 15914
rect 19444 15706 19472 16526
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19444 15026 19472 15642
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18800 13814 18828 14554
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 18892 14074 18920 14418
rect 18880 14068 18932 14074
rect 18932 14028 19012 14056
rect 18880 14010 18932 14016
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18432 12306 18460 13262
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18432 11898 18460 12242
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18524 9722 18552 13806
rect 18800 13786 18920 13814
rect 18788 12368 18840 12374
rect 18788 12310 18840 12316
rect 18800 11558 18828 12310
rect 18892 11762 18920 13786
rect 18984 12170 19012 14028
rect 19260 13530 19288 14418
rect 19444 13938 19472 14826
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19248 13524 19300 13530
rect 19168 13484 19248 13512
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 19168 12102 19196 13484
rect 19248 13466 19300 13472
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19444 12918 19472 13398
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19444 12442 19472 12854
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 11286 18828 11494
rect 18788 11280 18840 11286
rect 18788 11222 18840 11228
rect 18800 11014 18828 11222
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18800 10470 18828 10950
rect 19076 10742 19104 11086
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18800 10198 18828 10406
rect 18788 10192 18840 10198
rect 18788 10134 18840 10140
rect 17868 9658 17920 9664
rect 17880 9382 17908 9658
rect 17972 9646 18092 9674
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17788 8634 17816 8978
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17880 7546 17908 7958
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17972 6769 18000 9646
rect 18800 9586 18828 10134
rect 18892 9926 18920 10542
rect 19168 9976 19196 12038
rect 19340 10532 19392 10538
rect 19340 10474 19392 10480
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19260 10130 19288 10406
rect 19352 10130 19380 10474
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19076 9948 19196 9976
rect 18880 9920 18932 9926
rect 18880 9862 18932 9868
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18064 8498 18092 8910
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18156 7993 18184 9386
rect 18142 7984 18198 7993
rect 18142 7919 18198 7928
rect 18616 7886 18644 9522
rect 18892 9518 18920 9862
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 7410 18276 7686
rect 18800 7410 18828 7890
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18236 7268 18288 7274
rect 18156 7228 18236 7256
rect 17958 6760 18014 6769
rect 17958 6695 18014 6704
rect 18156 6662 18184 7228
rect 18236 7210 18288 7216
rect 18328 6928 18380 6934
rect 18328 6870 18380 6876
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 6254 18184 6598
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18248 5914 18276 6734
rect 18340 6322 18368 6870
rect 18800 6730 18828 7346
rect 18788 6724 18840 6730
rect 18788 6666 18840 6672
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 17500 5782 17552 5788
rect 17682 5808 17738 5817
rect 17682 5743 17738 5752
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 17696 4690 17724 5743
rect 18892 5030 18920 9454
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18984 8022 19012 8230
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 19076 7546 19104 9948
rect 19260 9722 19288 10066
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 19248 9376 19300 9382
rect 19352 9364 19380 10066
rect 19300 9336 19380 9364
rect 19248 9318 19300 9324
rect 19260 9042 19288 9318
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19168 8634 19196 8978
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19168 8090 19196 8570
rect 19260 8566 19288 8978
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19260 7546 19288 8502
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19076 7342 19104 7482
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 19352 2009 19380 8366
rect 19536 8090 19564 23598
rect 20260 23588 20312 23594
rect 20260 23530 20312 23536
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 19904 18154 19932 18770
rect 19892 18148 19944 18154
rect 19892 18090 19944 18096
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19812 16114 19840 16594
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14618 20024 19654
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 20088 18970 20116 19246
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 20088 17338 20116 18022
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20088 16726 20116 17138
rect 20180 16726 20208 18566
rect 20076 16720 20128 16726
rect 20076 16662 20128 16668
rect 20168 16720 20220 16726
rect 20168 16662 20220 16668
rect 20180 16250 20208 16662
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20272 15570 20300 23530
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 23308 22778 23336 23122
rect 23296 22772 23348 22778
rect 23296 22714 23348 22720
rect 23308 22438 23336 22714
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 22468 19984 22520 19990
rect 22468 19926 22520 19932
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20444 18352 20496 18358
rect 20444 18294 20496 18300
rect 20352 18148 20404 18154
rect 20352 18090 20404 18096
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20272 15026 20300 15506
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19996 14006 20024 14554
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19708 13796 19760 13802
rect 19984 13796 20036 13802
rect 19760 13756 19984 13784
rect 19708 13738 19760 13744
rect 19984 13738 20036 13744
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19628 12986 19656 13194
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19996 11830 20024 13738
rect 20088 12986 20116 14826
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 20180 14006 20208 14486
rect 20168 14000 20220 14006
rect 20168 13942 20220 13948
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20272 13462 20300 13806
rect 20260 13456 20312 13462
rect 20260 13398 20312 13404
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20088 12646 20116 12922
rect 20364 12850 20392 18090
rect 20456 17202 20484 18294
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20548 17270 20576 18022
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20640 16658 20668 17546
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20548 14346 20576 15846
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20640 14618 20668 15098
rect 20732 14822 20760 19246
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20824 18358 20852 18702
rect 21100 18426 21128 18838
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21088 18420 21140 18426
rect 21088 18362 21140 18368
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20824 16794 20852 18294
rect 21180 18148 21232 18154
rect 21180 18090 21232 18096
rect 21192 17882 21220 18090
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20916 17270 20944 17478
rect 21100 17338 21128 17750
rect 21284 17678 21312 18702
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 21468 17678 21496 18226
rect 22376 17808 22428 17814
rect 22376 17750 22428 17756
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20916 16794 20944 17206
rect 21284 17202 21312 17614
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20916 16250 20944 16730
rect 21284 16590 21312 17138
rect 22388 17066 22416 17750
rect 22376 17060 22428 17066
rect 22376 17002 22428 17008
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20824 15706 20852 16050
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 21088 15632 21140 15638
rect 21088 15574 21140 15580
rect 21100 15162 21128 15574
rect 21376 15502 21404 16118
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20456 13530 20484 13874
rect 20732 13814 20760 14758
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 21100 14074 21128 14486
rect 21376 14414 21404 15438
rect 22296 14618 22324 15846
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21376 14006 21404 14350
rect 22296 14074 22324 14554
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 20732 13786 20852 13814
rect 20916 13802 20944 13942
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 11354 20024 11766
rect 20088 11762 20116 12582
rect 20272 12102 20300 12718
rect 20352 12708 20404 12714
rect 20352 12650 20404 12656
rect 20364 12306 20392 12650
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 20272 11354 20300 12038
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20364 11150 20392 12242
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20456 10674 20484 11494
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 9042 20024 9998
rect 20180 9586 20208 10474
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20180 9178 20208 9522
rect 20732 9450 20760 9998
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20732 9110 20760 9386
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19996 8634 20024 8978
rect 20824 8634 20852 13786
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20996 13456 21048 13462
rect 20996 13398 21048 13404
rect 21088 13456 21140 13462
rect 21088 13398 21140 13404
rect 21008 13297 21036 13398
rect 20994 13288 21050 13297
rect 20994 13223 21050 13232
rect 21008 12442 21036 13223
rect 21100 12986 21128 13398
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 21100 12374 21128 12922
rect 22020 12850 22048 13262
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21560 12442 21588 12582
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 21008 11558 21036 12106
rect 21100 11898 21128 12310
rect 21560 11898 21588 12378
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21560 11626 21588 11834
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 21008 11218 21036 11494
rect 21836 11286 21864 11630
rect 21824 11280 21876 11286
rect 21824 11222 21876 11228
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21008 10470 21036 11154
rect 21284 10538 21312 11154
rect 22192 10736 22244 10742
rect 22192 10678 22244 10684
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 21008 10130 21036 10406
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 21100 9722 21128 10406
rect 21180 10192 21232 10198
rect 21180 10134 21232 10140
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21192 9382 21220 10134
rect 21376 9926 21404 10610
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 21928 10266 21956 10474
rect 22204 10266 22232 10678
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21008 9110 21036 9318
rect 21376 9110 21404 9862
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 21364 9104 21416 9110
rect 21364 9046 21416 9052
rect 21008 8634 21036 9046
rect 21836 8634 21864 9862
rect 21928 9654 21956 10202
rect 22376 10192 22428 10198
rect 22376 10134 22428 10140
rect 22284 9988 22336 9994
rect 22284 9930 22336 9936
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 20536 8288 20588 8294
rect 20536 8230 20588 8236
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20548 8090 20576 8230
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 21008 8022 21036 8570
rect 21732 8356 21784 8362
rect 21836 8344 21864 8570
rect 21928 8498 21956 9590
rect 22296 9586 22324 9930
rect 22388 9654 22416 10134
rect 22376 9648 22428 9654
rect 22376 9590 22428 9596
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 22112 9178 22140 9386
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 21784 8316 21864 8344
rect 21732 8298 21784 8304
rect 20996 8016 21048 8022
rect 20996 7958 21048 7964
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 19522 7304 19578 7313
rect 20364 7274 20392 7822
rect 21008 7546 21036 7958
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 21836 7274 21864 7686
rect 21928 7410 21956 8434
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 19522 7239 19578 7248
rect 20352 7268 20404 7274
rect 19536 6866 19564 7239
rect 20352 7210 20404 7216
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20364 6934 20392 7210
rect 21836 7002 21864 7210
rect 22376 7200 22428 7206
rect 22480 7177 22508 19926
rect 23400 18970 23428 22510
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23112 18828 23164 18834
rect 23112 18770 23164 18776
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22572 16998 22600 17614
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22572 16794 22600 16934
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 22756 16726 22784 18362
rect 23124 18290 23152 18770
rect 23112 18284 23164 18290
rect 23112 18226 23164 18232
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23110 17640 23166 17649
rect 23110 17575 23166 17584
rect 23124 17338 23152 17575
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23124 17134 23152 17274
rect 23216 17202 23244 17750
rect 23492 17610 23520 23666
rect 23860 23089 23888 23802
rect 24044 23594 24072 24686
rect 24032 23588 24084 23594
rect 24032 23530 24084 23536
rect 24136 23322 24164 27526
rect 24398 27520 24454 27526
rect 25778 27520 25834 28000
rect 27158 27520 27214 28000
rect 25226 26888 25282 26897
rect 25226 26823 25282 26832
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24766 24984 24822 24993
rect 24766 24919 24822 24928
rect 24780 24886 24808 24919
rect 24768 24880 24820 24886
rect 24768 24822 24820 24828
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23730 24716 24210
rect 24766 24032 24822 24041
rect 24766 23967 24822 23976
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24216 23520 24268 23526
rect 24216 23462 24268 23468
rect 24124 23316 24176 23322
rect 24124 23258 24176 23264
rect 24124 23180 24176 23186
rect 24124 23122 24176 23128
rect 23846 23080 23902 23089
rect 23846 23015 23902 23024
rect 24136 22574 24164 23122
rect 24124 22568 24176 22574
rect 24124 22510 24176 22516
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 23572 18216 23624 18222
rect 23572 18158 23624 18164
rect 23480 17604 23532 17610
rect 23480 17546 23532 17552
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 23216 16726 23244 17138
rect 22744 16720 22796 16726
rect 22744 16662 22796 16668
rect 23204 16720 23256 16726
rect 23204 16662 23256 16668
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22572 16250 22600 16526
rect 22560 16244 22612 16250
rect 22560 16186 22612 16192
rect 22756 16182 22784 16662
rect 22744 16176 22796 16182
rect 22744 16118 22796 16124
rect 23112 15632 23164 15638
rect 23112 15574 23164 15580
rect 23124 15162 23152 15574
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 23492 15094 23520 15438
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22664 13870 22692 14214
rect 22848 14006 22876 14894
rect 22928 14544 22980 14550
rect 22928 14486 22980 14492
rect 22940 14346 22968 14486
rect 22928 14340 22980 14346
rect 22928 14282 22980 14288
rect 22940 14006 22968 14282
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22664 12102 22692 13126
rect 22940 12646 22968 13398
rect 23204 13252 23256 13258
rect 23308 13240 23336 14214
rect 23584 13818 23612 18158
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 23860 17066 23888 17206
rect 23756 17060 23808 17066
rect 23756 17002 23808 17008
rect 23848 17060 23900 17066
rect 23848 17002 23900 17008
rect 23768 16590 23796 17002
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23756 16584 23808 16590
rect 23756 16526 23808 16532
rect 23952 16250 23980 16594
rect 23940 16244 23992 16250
rect 23860 16204 23940 16232
rect 23860 15638 23888 16204
rect 23940 16186 23992 16192
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 23952 15706 23980 15846
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 23848 15632 23900 15638
rect 23848 15574 23900 15580
rect 23848 15088 23900 15094
rect 23848 15030 23900 15036
rect 23860 14550 23888 15030
rect 23952 15026 23980 15642
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23848 14544 23900 14550
rect 23900 14504 23980 14532
rect 23848 14486 23900 14492
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23860 13938 23888 14214
rect 23952 13938 23980 14504
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 23256 13212 23336 13240
rect 23400 13790 23612 13818
rect 24044 13814 24072 22374
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 24136 18698 24164 20334
rect 24124 18692 24176 18698
rect 24124 18634 24176 18640
rect 24124 17740 24176 17746
rect 24124 17682 24176 17688
rect 24136 16998 24164 17682
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 24136 14074 24164 16934
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 24228 13814 24256 23462
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24780 22778 24808 23967
rect 25240 23322 25268 26823
rect 25502 25800 25558 25809
rect 25502 25735 25558 25744
rect 25516 24410 25544 25735
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 25792 24138 25820 27520
rect 25780 24132 25832 24138
rect 25780 24074 25832 24080
rect 27172 23866 27200 27520
rect 27160 23860 27212 23866
rect 27160 23802 27212 23808
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24766 22672 24822 22681
rect 24766 22607 24822 22616
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24780 21690 24808 22607
rect 24858 21720 24914 21729
rect 24768 21684 24820 21690
rect 24858 21655 24914 21664
rect 24768 21626 24820 21632
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 16794 24716 21422
rect 24766 20632 24822 20641
rect 24872 20602 24900 21655
rect 24766 20567 24822 20576
rect 24860 20596 24912 20602
rect 24780 19514 24808 20567
rect 24860 20538 24912 20544
rect 24858 19544 24914 19553
rect 24768 19508 24820 19514
rect 24858 19479 24914 19488
rect 24768 19450 24820 19456
rect 24766 18592 24822 18601
rect 24766 18527 24822 18536
rect 24780 17882 24808 18527
rect 24872 18426 24900 19479
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 24858 16552 24914 16561
rect 24858 16487 24914 16496
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24584 16176 24636 16182
rect 24584 16118 24636 16124
rect 24596 15706 24624 16118
rect 24872 16114 24900 16487
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 25608 15910 25636 16594
rect 27620 16108 27672 16114
rect 27620 16050 27672 16056
rect 27632 16017 27660 16050
rect 27618 16008 27674 16017
rect 27618 15943 27674 15952
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 25596 15904 25648 15910
rect 25596 15846 25648 15852
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24492 14884 24544 14890
rect 24492 14826 24544 14832
rect 24504 14414 24532 14826
rect 24492 14408 24544 14414
rect 24688 14396 24716 15846
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24780 15026 24808 15506
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24860 14544 24912 14550
rect 24860 14486 24912 14492
rect 25410 14512 25466 14521
rect 24768 14408 24820 14414
rect 24688 14368 24768 14396
rect 24492 14350 24544 14356
rect 24768 14350 24820 14356
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24780 13938 24808 14350
rect 24872 14074 24900 14486
rect 25410 14447 25466 14456
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24964 14074 24992 14214
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 23204 13194 23256 13200
rect 23216 12850 23244 13194
rect 23204 12844 23256 12850
rect 23204 12786 23256 12792
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22940 12442 22968 12582
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 23204 12300 23256 12306
rect 23204 12242 23256 12248
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22664 11082 22692 12038
rect 23216 11286 23244 12242
rect 23400 11540 23428 13790
rect 23952 13786 24072 13814
rect 24136 13786 24256 13814
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23480 13456 23532 13462
rect 23480 13398 23532 13404
rect 23492 12986 23520 13398
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23768 12714 23796 13466
rect 23756 12708 23808 12714
rect 23756 12650 23808 12656
rect 23848 12708 23900 12714
rect 23848 12650 23900 12656
rect 23860 12442 23888 12650
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23860 11898 23888 12378
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23952 11830 23980 13786
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23572 11688 23624 11694
rect 23572 11630 23624 11636
rect 23308 11512 23428 11540
rect 23204 11280 23256 11286
rect 23204 11222 23256 11228
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 22652 11076 22704 11082
rect 22652 11018 22704 11024
rect 23124 10810 23152 11086
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 23216 10674 23244 11222
rect 23204 10668 23256 10674
rect 23204 10610 23256 10616
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 22940 9722 22968 10066
rect 22928 9716 22980 9722
rect 22928 9658 22980 9664
rect 23124 9382 23152 10066
rect 23308 9586 23336 11512
rect 23584 10810 23612 11630
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23584 10470 23612 10746
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23768 10266 23796 10474
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23768 9926 23796 10202
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 23400 9178 23428 9862
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 22664 8294 22692 8978
rect 22652 8288 22704 8294
rect 22652 8230 22704 8236
rect 22664 7449 22692 8230
rect 23676 7993 23704 9318
rect 23860 9042 23888 9590
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23860 8634 23888 8978
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23662 7984 23718 7993
rect 23662 7919 23718 7928
rect 22650 7440 22706 7449
rect 22650 7375 22706 7384
rect 22376 7142 22428 7148
rect 22466 7168 22522 7177
rect 21824 6996 21876 7002
rect 21824 6938 21876 6944
rect 20352 6928 20404 6934
rect 20352 6870 20404 6876
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19536 6458 19564 6802
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 22388 4826 22416 7142
rect 22466 7103 22522 7112
rect 23952 5137 23980 11766
rect 24032 11076 24084 11082
rect 24032 11018 24084 11024
rect 24044 10674 24072 11018
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 24032 10532 24084 10538
rect 24032 10474 24084 10480
rect 24044 10130 24072 10474
rect 24136 10266 24164 13786
rect 24872 13462 24900 14010
rect 25056 13530 25084 14350
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 24860 13456 24912 13462
rect 24860 13398 24912 13404
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24228 12986 24256 13262
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 25056 12374 25084 13466
rect 25044 12368 25096 12374
rect 24674 12336 24730 12345
rect 25044 12310 25096 12316
rect 24674 12271 24730 12280
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 24228 11898 24256 12174
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 24032 10124 24084 10130
rect 24032 10066 24084 10072
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 24136 9722 24164 9998
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 23938 5128 23994 5137
rect 23938 5063 23994 5072
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 21744 4282 21772 4626
rect 21732 4276 21784 4282
rect 21732 4218 21784 4224
rect 24228 4154 24256 11698
rect 24398 11656 24454 11665
rect 24398 11591 24454 11600
rect 24412 11354 24440 11591
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9722 24716 12271
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24780 10470 24808 11154
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 24780 9353 24808 10406
rect 24872 9722 24900 11834
rect 25056 11762 25084 12310
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 25148 11150 25176 11494
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 25424 10810 25452 14447
rect 25608 12073 25636 15846
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27632 14929 27660 14962
rect 27618 14920 27674 14929
rect 27618 14855 27674 14864
rect 25780 14816 25832 14822
rect 25780 14758 25832 14764
rect 25792 14521 25820 14758
rect 25778 14512 25834 14521
rect 25778 14447 25834 14456
rect 25780 13796 25832 13802
rect 25780 13738 25832 13744
rect 25594 12064 25650 12073
rect 25594 11999 25650 12008
rect 25792 11393 25820 13738
rect 25778 11384 25834 11393
rect 25778 11319 25834 11328
rect 25412 10804 25464 10810
rect 25412 10746 25464 10752
rect 25226 10704 25282 10713
rect 25226 10639 25282 10648
rect 25240 10266 25268 10639
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 25332 9654 25360 10066
rect 27618 9752 27674 9761
rect 27618 9687 27674 9696
rect 27632 9654 27660 9687
rect 25320 9648 25372 9654
rect 25320 9590 25372 9596
rect 27620 9648 27672 9654
rect 27620 9590 27672 9596
rect 24766 9344 24822 9353
rect 24766 9279 24822 9288
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 27712 8288 27764 8294
rect 27712 8230 27764 8236
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24136 4126 24256 4154
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 23294 3632 23350 3641
rect 23294 3567 23350 3576
rect 19430 2816 19486 2825
rect 19430 2751 19486 2760
rect 19338 2000 19394 2009
rect 19338 1935 19394 1944
rect 16946 82 17002 480
rect 19444 134 19472 2751
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 16776 54 17002 82
rect 19432 128 19484 134
rect 19432 70 19484 76
rect 20074 128 20130 480
rect 20074 76 20076 128
rect 20128 76 20130 128
rect 10782 0 10838 54
rect 13910 0 13966 54
rect 16946 0 17002 54
rect 20074 0 20130 76
rect 23202 82 23258 480
rect 23308 82 23336 3567
rect 24136 2650 24164 4126
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24124 2644 24176 2650
rect 24124 2586 24176 2592
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25148 2310 25176 2450
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 25148 1057 25176 2246
rect 25134 1048 25190 1057
rect 25134 983 25190 992
rect 23202 54 23336 82
rect 25976 82 26004 7482
rect 27618 4584 27674 4593
rect 27618 4519 27674 4528
rect 27632 4282 27660 4519
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27724 1465 27752 8230
rect 27710 1456 27766 1465
rect 27710 1391 27766 1400
rect 26330 82 26386 480
rect 25976 54 26386 82
rect 23202 0 23258 54
rect 26330 0 26386 54
<< via2 >>
rect 1306 27104 1362 27160
rect 110 20032 166 20088
rect 110 19080 166 19136
rect 1490 25744 1546 25800
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 1582 24792 1638 24848
rect 1582 23976 1638 24032
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 1490 22616 1546 22672
rect 1582 21664 1638 21720
rect 1214 15272 1270 15328
rect 1306 12280 1362 12336
rect 1214 10240 1270 10296
rect 110 9696 166 9752
rect 110 8744 166 8800
rect 110 7656 166 7712
rect 1950 17584 2006 17640
rect 1858 15408 1914 15464
rect 2042 11192 2098 11248
rect 2686 20576 2742 20632
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 3054 21392 3110 21448
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 3974 18536 4030 18592
rect 2686 13640 2742 13696
rect 3606 11192 3662 11248
rect 4066 8064 4122 8120
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5262 15408 5318 15464
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 9034 22616 9090 22672
rect 7378 19216 7434 19272
rect 6274 18264 6330 18320
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 7930 18808 7986 18864
rect 7838 17720 7894 17776
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 2318 7384 2374 7440
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 8298 13912 8354 13968
rect 8482 13232 8538 13288
rect 8298 8064 8354 8120
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 8942 7792 8998 7848
rect 8298 7248 8354 7304
rect 110 6840 166 6896
rect 110 5616 166 5672
rect 1766 5208 1822 5264
rect 110 3440 166 3496
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 9126 6296 9182 6352
rect 7562 5616 7618 5672
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5538 1400 5594 1456
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10138 10648 10194 10704
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 11334 11192 11390 11248
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 9862 5208 9918 5264
rect 9862 2624 9918 2680
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10782 3576 10838 3632
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10046 1264 10102 1320
rect 12898 11600 12954 11656
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 15106 23024 15162 23080
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 17590 22616 17646 22672
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 19246 21392 19302 21448
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14002 17720 14058 17776
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15566 18264 15622 18320
rect 16210 18808 16266 18864
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14738 13948 14740 13968
rect 14740 13948 14792 13968
rect 14792 13948 14794 13968
rect 14738 13912 14794 13948
rect 15934 14456 15990 14512
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 17774 15408 17830 15464
rect 16210 10648 16266 10704
rect 16394 10648 16450 10704
rect 12714 2896 12770 2952
rect 11518 2760 11574 2816
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14554 5616 14610 5672
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 19430 19216 19486 19272
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 17406 7792 17462 7848
rect 18142 7928 18198 7984
rect 17958 6704 18014 6760
rect 17682 5752 17738 5808
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 20994 13232 21050 13288
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19522 7248 19578 7304
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 23110 17584 23166 17640
rect 25226 26832 25282 26888
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 24928 24822 24984
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 23976 24822 24032
rect 23846 23024 23902 23080
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 25502 25744 25558 25800
rect 24766 22616 24822 22672
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24858 21664 24914 21720
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24766 20576 24822 20632
rect 24858 19488 24914 19544
rect 24766 18536 24822 18592
rect 24858 16496 24914 16552
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 27618 15952 27674 16008
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 25410 14456 25466 14512
rect 23662 7928 23718 7984
rect 22650 7384 22706 7440
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 22466 7112 22522 7168
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24674 12280 24730 12336
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 23938 5072 23994 5128
rect 24398 11600 24454 11656
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 27618 14864 27674 14920
rect 25778 14456 25834 14512
rect 25594 12008 25650 12064
rect 25778 11328 25834 11384
rect 25226 10648 25282 10704
rect 27618 9696 27674 9752
rect 24766 9288 24822 9344
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 23294 3576 23350 3632
rect 19430 2760 19486 2816
rect 19338 1944 19394 2000
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25134 992 25190 1048
rect 27618 4528 27674 4584
rect 27710 1400 27766 1456
<< metal3 >>
rect 0 27344 480 27464
rect 27520 27344 28000 27464
rect 62 27162 122 27344
rect 1301 27162 1367 27165
rect 62 27160 1367 27162
rect 62 27104 1306 27160
rect 1362 27104 1367 27160
rect 62 27102 1367 27104
rect 1301 27099 1367 27102
rect 25221 26890 25287 26893
rect 27662 26890 27722 27344
rect 25221 26888 27722 26890
rect 25221 26832 25226 26888
rect 25282 26832 27722 26888
rect 25221 26830 27722 26832
rect 25221 26827 25287 26830
rect 0 26256 480 26376
rect 27520 26256 28000 26376
rect 62 25802 122 26256
rect 1485 25802 1551 25805
rect 62 25800 1551 25802
rect 62 25744 1490 25800
rect 1546 25744 1551 25800
rect 62 25742 1551 25744
rect 1485 25739 1551 25742
rect 25497 25802 25563 25805
rect 27662 25802 27722 26256
rect 25497 25800 27722 25802
rect 25497 25744 25502 25800
rect 25558 25744 27722 25800
rect 25497 25742 27722 25744
rect 25497 25739 25563 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25304 480 25424
rect 27520 25304 28000 25424
rect 62 24850 122 25304
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 24761 24986 24827 24989
rect 27662 24986 27722 25304
rect 24761 24984 27722 24986
rect 24761 24928 24766 24984
rect 24822 24928 27722 24984
rect 24761 24926 27722 24928
rect 24761 24923 24827 24926
rect 1577 24850 1643 24853
rect 62 24848 1643 24850
rect 62 24792 1582 24848
rect 1638 24792 1643 24848
rect 62 24790 1643 24792
rect 1577 24787 1643 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24216 480 24336
rect 27520 24216 28000 24336
rect 62 24034 122 24216
rect 1577 24034 1643 24037
rect 62 24032 1643 24034
rect 62 23976 1582 24032
rect 1638 23976 1643 24032
rect 62 23974 1643 23976
rect 1577 23971 1643 23974
rect 24761 24034 24827 24037
rect 27662 24034 27722 24216
rect 24761 24032 27722 24034
rect 24761 23976 24766 24032
rect 24822 23976 27722 24032
rect 24761 23974 27722 23976
rect 24761 23971 24827 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23128 480 23248
rect 27520 23128 28000 23248
rect 62 22674 122 23128
rect 15101 23082 15167 23085
rect 23841 23082 23907 23085
rect 15101 23080 23907 23082
rect 15101 23024 15106 23080
rect 15162 23024 23846 23080
rect 23902 23024 23907 23080
rect 15101 23022 23907 23024
rect 15101 23019 15167 23022
rect 23841 23019 23907 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1485 22674 1551 22677
rect 62 22672 1551 22674
rect 62 22616 1490 22672
rect 1546 22616 1551 22672
rect 62 22614 1551 22616
rect 1485 22611 1551 22614
rect 9029 22674 9095 22677
rect 17585 22674 17651 22677
rect 9029 22672 17651 22674
rect 9029 22616 9034 22672
rect 9090 22616 17590 22672
rect 17646 22616 17651 22672
rect 9029 22614 17651 22616
rect 9029 22611 9095 22614
rect 17585 22611 17651 22614
rect 24761 22674 24827 22677
rect 27662 22674 27722 23128
rect 24761 22672 27722 22674
rect 24761 22616 24766 22672
rect 24822 22616 27722 22672
rect 24761 22614 27722 22616
rect 24761 22611 24827 22614
rect 10277 22336 10597 22337
rect 0 22176 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 27520 22176 28000 22296
rect 62 21722 122 22176
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 1577 21722 1643 21725
rect 62 21720 1643 21722
rect 62 21664 1582 21720
rect 1638 21664 1643 21720
rect 62 21662 1643 21664
rect 1577 21659 1643 21662
rect 24853 21722 24919 21725
rect 27662 21722 27722 22176
rect 24853 21720 27722 21722
rect 24853 21664 24858 21720
rect 24914 21664 27722 21720
rect 24853 21662 27722 21664
rect 24853 21659 24919 21662
rect 3049 21450 3115 21453
rect 19241 21450 19307 21453
rect 3049 21448 19307 21450
rect 3049 21392 3054 21448
rect 3110 21392 19246 21448
rect 19302 21392 19307 21448
rect 3049 21390 19307 21392
rect 3049 21387 3115 21390
rect 19241 21387 19307 21390
rect 10277 21248 10597 21249
rect 0 21088 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 27520 21088 28000 21208
rect 62 20634 122 21088
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 2681 20634 2747 20637
rect 62 20632 2747 20634
rect 62 20576 2686 20632
rect 2742 20576 2747 20632
rect 62 20574 2747 20576
rect 2681 20571 2747 20574
rect 24761 20634 24827 20637
rect 27662 20634 27722 21088
rect 24761 20632 27722 20634
rect 24761 20576 24766 20632
rect 24822 20576 27722 20632
rect 24761 20574 27722 20576
rect 24761 20571 24827 20574
rect 10277 20160 10597 20161
rect 0 20088 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 20032 110 20088
rect 166 20032 480 20088
rect 0 20000 480 20032
rect 27520 20000 28000 20120
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 24853 19546 24919 19549
rect 27662 19546 27722 20000
rect 24853 19544 27722 19546
rect 24853 19488 24858 19544
rect 24914 19488 27722 19544
rect 24853 19486 27722 19488
rect 24853 19483 24919 19486
rect 7373 19274 7439 19277
rect 19425 19274 19491 19277
rect 7373 19272 19491 19274
rect 7373 19216 7378 19272
rect 7434 19216 19430 19272
rect 19486 19216 19491 19272
rect 7373 19214 19491 19216
rect 7373 19211 7439 19214
rect 19425 19211 19491 19214
rect 0 19136 480 19168
rect 0 19080 110 19136
rect 166 19080 480 19136
rect 0 19048 480 19080
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19168
rect 19610 19007 19930 19008
rect 7925 18866 7991 18869
rect 16205 18866 16271 18869
rect 7925 18864 16271 18866
rect 7925 18808 7930 18864
rect 7986 18808 16210 18864
rect 16266 18808 16271 18864
rect 7925 18806 16271 18808
rect 7925 18803 7991 18806
rect 16205 18803 16271 18806
rect 3969 18594 4035 18597
rect 62 18592 4035 18594
rect 62 18536 3974 18592
rect 4030 18536 4035 18592
rect 62 18534 4035 18536
rect 62 18080 122 18534
rect 3969 18531 4035 18534
rect 24761 18594 24827 18597
rect 27662 18594 27722 19048
rect 24761 18592 27722 18594
rect 24761 18536 24766 18592
rect 24822 18536 27722 18592
rect 24761 18534 27722 18536
rect 24761 18531 24827 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 6269 18322 6335 18325
rect 15561 18322 15627 18325
rect 6269 18320 15627 18322
rect 6269 18264 6274 18320
rect 6330 18264 15566 18320
rect 15622 18264 15627 18320
rect 6269 18262 15627 18264
rect 6269 18259 6335 18262
rect 15561 18259 15627 18262
rect 0 17960 480 18080
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 18080
rect 19610 17919 19930 17920
rect 7833 17778 7899 17781
rect 13997 17778 14063 17781
rect 7833 17776 14063 17778
rect 7833 17720 7838 17776
rect 7894 17720 14002 17776
rect 14058 17720 14063 17776
rect 7833 17718 14063 17720
rect 7833 17715 7899 17718
rect 13997 17715 14063 17718
rect 1945 17642 2011 17645
rect 62 17640 2011 17642
rect 62 17584 1950 17640
rect 2006 17584 2011 17640
rect 62 17582 2011 17584
rect 62 17128 122 17582
rect 1945 17579 2011 17582
rect 23105 17642 23171 17645
rect 27662 17642 27722 17960
rect 23105 17640 27722 17642
rect 23105 17584 23110 17640
rect 23166 17584 27722 17640
rect 23105 17582 27722 17584
rect 23105 17579 23171 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 0 17008 480 17128
rect 27520 17008 28000 17128
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 24853 16554 24919 16557
rect 27662 16554 27722 17008
rect 24853 16552 27722 16554
rect 24853 16496 24858 16552
rect 24914 16496 27722 16552
rect 24853 16494 27722 16496
rect 24853 16491 24919 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 15920 480 16040
rect 27520 16008 28000 16040
rect 27520 15952 27618 16008
rect 27674 15952 28000 16008
rect 27520 15920 28000 15952
rect 62 15466 122 15920
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 1853 15466 1919 15469
rect 62 15464 1919 15466
rect 62 15408 1858 15464
rect 1914 15408 1919 15464
rect 62 15406 1919 15408
rect 1853 15403 1919 15406
rect 5257 15466 5323 15469
rect 17769 15466 17835 15469
rect 5257 15464 17835 15466
rect 5257 15408 5262 15464
rect 5318 15408 17774 15464
rect 17830 15408 17835 15464
rect 5257 15406 17835 15408
rect 5257 15403 5323 15406
rect 17769 15403 17835 15406
rect 1209 15330 1275 15333
rect 62 15328 1275 15330
rect 62 15272 1214 15328
rect 1270 15272 1275 15328
rect 62 15270 1275 15272
rect 62 14952 122 15270
rect 1209 15267 1275 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14832 480 14952
rect 27520 14920 28000 14952
rect 27520 14864 27618 14920
rect 27674 14864 28000 14920
rect 27520 14832 28000 14864
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 15929 14514 15995 14517
rect 25405 14514 25471 14517
rect 15929 14512 25471 14514
rect 15929 14456 15934 14512
rect 15990 14456 25410 14512
rect 25466 14456 25471 14512
rect 15929 14454 25471 14456
rect 15929 14451 15995 14454
rect 25405 14451 25471 14454
rect 25773 14514 25839 14517
rect 25773 14512 27722 14514
rect 25773 14456 25778 14512
rect 25834 14456 27722 14512
rect 25773 14454 27722 14456
rect 25773 14451 25839 14454
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 27662 14000 27722 14454
rect 0 13880 480 14000
rect 8293 13970 8359 13973
rect 14733 13970 14799 13973
rect 8293 13968 14799 13970
rect 8293 13912 8298 13968
rect 8354 13912 14738 13968
rect 14794 13912 14799 13968
rect 8293 13910 14799 13912
rect 8293 13907 8359 13910
rect 14733 13907 14799 13910
rect 27520 13880 28000 14000
rect 62 13698 122 13880
rect 2681 13698 2747 13701
rect 62 13696 2747 13698
rect 62 13640 2686 13696
rect 2742 13640 2747 13696
rect 62 13638 2747 13640
rect 2681 13635 2747 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 8477 13290 8543 13293
rect 20989 13290 21055 13293
rect 8477 13288 21055 13290
rect 8477 13232 8482 13288
rect 8538 13232 20994 13288
rect 21050 13232 21055 13288
rect 8477 13230 21055 13232
rect 8477 13227 8543 13230
rect 20989 13227 21055 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 0 12792 480 12912
rect 27520 12792 28000 12912
rect 62 12338 122 12792
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 1301 12338 1367 12341
rect 62 12336 1367 12338
rect 62 12280 1306 12336
rect 1362 12280 1367 12336
rect 62 12278 1367 12280
rect 1301 12275 1367 12278
rect 24669 12338 24735 12341
rect 27662 12338 27722 12792
rect 24669 12336 27722 12338
rect 24669 12280 24674 12336
rect 24730 12280 27722 12336
rect 24669 12278 27722 12280
rect 24669 12275 24735 12278
rect 25589 12066 25655 12069
rect 25589 12064 27722 12066
rect 25589 12008 25594 12064
rect 25650 12008 27722 12064
rect 25589 12006 27722 12008
rect 25589 12003 25655 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 27662 11824 27722 12006
rect 0 11704 480 11824
rect 27520 11704 28000 11824
rect 62 11250 122 11704
rect 12893 11658 12959 11661
rect 24393 11658 24459 11661
rect 12893 11656 24459 11658
rect 12893 11600 12898 11656
rect 12954 11600 24398 11656
rect 24454 11600 24459 11656
rect 12893 11598 24459 11600
rect 12893 11595 12959 11598
rect 24393 11595 24459 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 25773 11386 25839 11389
rect 25773 11384 27722 11386
rect 25773 11328 25778 11384
rect 25834 11328 27722 11384
rect 25773 11326 27722 11328
rect 25773 11323 25839 11326
rect 2037 11250 2103 11253
rect 62 11248 2103 11250
rect 62 11192 2042 11248
rect 2098 11192 2103 11248
rect 62 11190 2103 11192
rect 2037 11187 2103 11190
rect 3601 11250 3667 11253
rect 11329 11250 11395 11253
rect 3601 11248 11395 11250
rect 3601 11192 3606 11248
rect 3662 11192 11334 11248
rect 11390 11192 11395 11248
rect 3601 11190 11395 11192
rect 3601 11187 3667 11190
rect 11329 11187 11395 11190
rect 5610 10912 5930 10913
rect 0 10752 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 27662 10872 27722 11326
rect 24277 10847 24597 10848
rect 27520 10752 28000 10872
rect 62 10298 122 10752
rect 10133 10706 10199 10709
rect 16205 10706 16271 10709
rect 10133 10704 16271 10706
rect 10133 10648 10138 10704
rect 10194 10648 16210 10704
rect 16266 10648 16271 10704
rect 10133 10646 16271 10648
rect 10133 10643 10199 10646
rect 16205 10643 16271 10646
rect 16389 10706 16455 10709
rect 25221 10706 25287 10709
rect 16389 10704 25287 10706
rect 16389 10648 16394 10704
rect 16450 10648 25226 10704
rect 25282 10648 25287 10704
rect 16389 10646 25287 10648
rect 16389 10643 16455 10646
rect 25221 10643 25287 10646
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 1209 10298 1275 10301
rect 62 10296 1275 10298
rect 62 10240 1214 10296
rect 1270 10240 1275 10296
rect 62 10238 1275 10240
rect 1209 10235 1275 10238
rect 5610 9824 5930 9825
rect 0 9752 480 9784
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 0 9696 110 9752
rect 166 9696 480 9752
rect 0 9664 480 9696
rect 27520 9752 28000 9784
rect 27520 9696 27618 9752
rect 27674 9696 28000 9752
rect 27520 9664 28000 9696
rect 24761 9346 24827 9349
rect 24761 9344 27722 9346
rect 24761 9288 24766 9344
rect 24822 9288 27722 9344
rect 24761 9286 27722 9288
rect 24761 9283 24827 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 27662 8832 27722 9286
rect 0 8800 480 8832
rect 0 8744 110 8800
rect 166 8744 480 8800
rect 0 8712 480 8744
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8832
rect 24277 8671 24597 8672
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 4061 8122 4127 8125
rect 8293 8122 8359 8125
rect 4061 8120 8359 8122
rect 4061 8064 4066 8120
rect 4122 8064 8298 8120
rect 8354 8064 8359 8120
rect 4061 8062 8359 8064
rect 4061 8059 4127 8062
rect 8293 8059 8359 8062
rect 18137 7986 18203 7989
rect 23657 7986 23723 7989
rect 18137 7984 23723 7986
rect 18137 7928 18142 7984
rect 18198 7928 23662 7984
rect 23718 7928 23723 7984
rect 18137 7926 23723 7928
rect 18137 7923 18203 7926
rect 23657 7923 23723 7926
rect 8937 7850 9003 7853
rect 17401 7850 17467 7853
rect 8937 7848 17467 7850
rect 8937 7792 8942 7848
rect 8998 7792 17406 7848
rect 17462 7792 17467 7848
rect 8937 7790 17467 7792
rect 8937 7787 9003 7790
rect 17401 7787 17467 7790
rect 0 7712 480 7744
rect 0 7656 110 7712
rect 166 7656 480 7712
rect 0 7624 480 7656
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7744
rect 24277 7583 24597 7584
rect 2313 7442 2379 7445
rect 22645 7442 22711 7445
rect 2313 7440 22711 7442
rect 2313 7384 2318 7440
rect 2374 7384 22650 7440
rect 22706 7384 22711 7440
rect 2313 7382 22711 7384
rect 2313 7379 2379 7382
rect 22645 7379 22711 7382
rect 8293 7306 8359 7309
rect 19517 7306 19583 7309
rect 27662 7306 27722 7624
rect 8293 7304 27722 7306
rect 8293 7248 8298 7304
rect 8354 7248 19522 7304
rect 19578 7248 27722 7304
rect 8293 7246 27722 7248
rect 8293 7243 8359 7246
rect 19517 7243 19583 7246
rect 22461 7170 22527 7173
rect 22461 7168 27722 7170
rect 22461 7112 22466 7168
rect 22522 7112 27722 7168
rect 22461 7110 27722 7112
rect 22461 7107 22527 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 105 6898 171 6901
rect 105 6896 9690 6898
rect 105 6840 110 6896
rect 166 6840 9690 6896
rect 105 6838 9690 6840
rect 105 6835 171 6838
rect 9630 6762 9690 6838
rect 17953 6762 18019 6765
rect 9630 6760 18019 6762
rect 9630 6704 17958 6760
rect 18014 6704 18019 6760
rect 9630 6702 18019 6704
rect 17953 6699 18019 6702
rect 27662 6656 27722 7110
rect 0 6536 480 6656
rect 5610 6560 5930 6561
rect 62 5946 122 6536
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6656
rect 24277 6495 24597 6496
rect 9121 6354 9187 6357
rect 9121 6352 27722 6354
rect 9121 6296 9126 6352
rect 9182 6296 27722 6352
rect 9121 6294 27722 6296
rect 9121 6291 9187 6294
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 62 5886 9690 5946
rect 9630 5810 9690 5886
rect 17677 5810 17743 5813
rect 9630 5808 17743 5810
rect 9630 5752 17682 5808
rect 17738 5752 17743 5808
rect 9630 5750 17743 5752
rect 17677 5747 17743 5750
rect 27662 5704 27722 6294
rect 0 5672 480 5704
rect 0 5616 110 5672
rect 166 5616 480 5672
rect 0 5584 480 5616
rect 7557 5674 7623 5677
rect 14549 5674 14615 5677
rect 7557 5672 14615 5674
rect 7557 5616 7562 5672
rect 7618 5616 14554 5672
rect 14610 5616 14615 5672
rect 7557 5614 14615 5616
rect 7557 5611 7623 5614
rect 14549 5611 14615 5614
rect 27520 5584 28000 5704
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 1761 5266 1827 5269
rect 9857 5266 9923 5269
rect 1761 5264 9923 5266
rect 1761 5208 1766 5264
rect 1822 5208 9862 5264
rect 9918 5208 9923 5264
rect 1761 5206 9923 5208
rect 1761 5203 1827 5206
rect 9857 5203 9923 5206
rect 23933 5130 23999 5133
rect 62 5128 23999 5130
rect 62 5072 23938 5128
rect 23994 5072 23999 5128
rect 62 5070 23999 5072
rect 62 4616 122 5070
rect 23933 5067 23999 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 0 4496 480 4616
rect 27520 4584 28000 4616
rect 27520 4528 27618 4584
rect 27674 4528 28000 4584
rect 27520 4496 28000 4528
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 10777 3634 10843 3637
rect 23289 3634 23355 3637
rect 10777 3632 23355 3634
rect 10777 3576 10782 3632
rect 10838 3576 23294 3632
rect 23350 3576 23355 3632
rect 10777 3574 23355 3576
rect 10777 3571 10843 3574
rect 23289 3571 23355 3574
rect 0 3496 480 3528
rect 0 3440 110 3496
rect 166 3440 480 3496
rect 0 3408 480 3440
rect 27520 3408 28000 3528
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 12709 2954 12775 2957
rect 27662 2954 27722 3408
rect 12709 2952 27722 2954
rect 12709 2896 12714 2952
rect 12770 2896 27722 2952
rect 12709 2894 27722 2896
rect 12709 2891 12775 2894
rect 54 2756 60 2820
rect 124 2818 130 2820
rect 11513 2818 11579 2821
rect 19425 2818 19491 2821
rect 124 2758 9690 2818
rect 124 2756 130 2758
rect 9630 2682 9690 2758
rect 11513 2816 19491 2818
rect 11513 2760 11518 2816
rect 11574 2760 19430 2816
rect 19486 2760 19491 2816
rect 11513 2758 19491 2760
rect 11513 2755 11579 2758
rect 19425 2755 19491 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 9857 2682 9923 2685
rect 9630 2680 9923 2682
rect 9630 2624 9862 2680
rect 9918 2624 9923 2680
rect 9630 2622 9923 2624
rect 9857 2619 9923 2622
rect 0 2548 480 2576
rect 0 2484 60 2548
rect 124 2484 480 2548
rect 0 2456 480 2484
rect 27520 2456 28000 2576
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 19333 2002 19399 2005
rect 62 2000 19399 2002
rect 62 1944 19338 2000
rect 19394 1944 19399 2000
rect 62 1942 19399 1944
rect 62 1488 122 1942
rect 19333 1939 19399 1942
rect 27662 1730 27722 2456
rect 19290 1670 27722 1730
rect 19290 1594 19350 1670
rect 13770 1534 19350 1594
rect 0 1368 480 1488
rect 5533 1458 5599 1461
rect 13770 1458 13830 1534
rect 5533 1456 13830 1458
rect 5533 1400 5538 1456
rect 5594 1400 13830 1456
rect 5533 1398 13830 1400
rect 27520 1456 28000 1488
rect 27520 1400 27710 1456
rect 27766 1400 28000 1456
rect 5533 1395 5599 1398
rect 27520 1368 28000 1400
rect 10041 1322 10107 1325
rect 9630 1320 10107 1322
rect 9630 1264 10046 1320
rect 10102 1264 10107 1320
rect 9630 1262 10107 1264
rect 9630 1186 9690 1262
rect 10041 1259 10107 1262
rect 62 1126 9690 1186
rect 62 536 122 1126
rect 25129 1050 25195 1053
rect 25129 1048 27722 1050
rect 25129 992 25134 1048
rect 25190 992 27722 1048
rect 25129 990 27722 992
rect 25129 987 25195 990
rect 27662 536 27722 990
rect 0 416 480 536
rect 27520 416 28000 536
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 60 2756 124 2820
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 60 2484 124 2548
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 59 2820 125 2821
rect 59 2756 60 2820
rect 124 2756 125 2820
rect 59 2755 125 2756
rect 62 2549 122 2755
rect 59 2548 125 2549
rect 59 2484 60 2548
rect 124 2484 125 2548
rect 59 2483 125 2484
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_7
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_19
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_43
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_55
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_269 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_30 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_106
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_169
timestamp 1586364061
transform 1 0 16652 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_181
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_224
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_227
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_8  _072_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_101
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_137
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_162
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_170
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_174
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_198
timestamp 1586364061
transform 1 0 19320 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21804 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_223
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_240
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_252
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_264
timestamp 1586364061
transform 1 0 25392 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_272
timestamp 1586364061
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 774 592
use scs8hd_inv_8  _117_
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_97
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__C
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__C
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_133
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_137
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_141
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _092_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 314 592
use scs8hd_buf_1  _166_
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_146
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_157
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _146_
timestamp 1586364061
transform 1 0 16284 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_161
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_182
timestamp 1586364061
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_97
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_or2_4  _118_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 682 592
use scs8hd_fill_2  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_101
timestamp 1586364061
transform 1 0 10396 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_or3_4  _149_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use scs8hd_nand3_4  _073_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 1326 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_118
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_130
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_126
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_126
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_or2_4  _096_
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 682 592
use scs8hd_fill_2  FILLER_6_142
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_nor3_4  _162_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 1234 592
use scs8hd_fill_2  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_146
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_168
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_162
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_176
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_172
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_conb_1  _183_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_179
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_216
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_228
timestamp 1586364061
transform 1 0 22080 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__D
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_8  _066_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 774 592
use scs8hd_nor3_4  _161_
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_1  _089_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 14720 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__C
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__078__C
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_165
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_177
timestamp 1586364061
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17940 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_181
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_194
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_219
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_222
timestamp 1586364061
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_226
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_238
timestamp 1586364061
transform 1 0 23000 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_250
timestamp 1586364061
transform 1 0 24104 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_262
timestamp 1586364061
transform 1 0 25208 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_28
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__C
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_80
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_87
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _070_
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use scs8hd_or3_4  _165_
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_139
timestamp 1586364061
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use scs8hd_or3_4  _088_
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_161
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_165
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _171_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_214
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_229
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_233
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_17
timestamp 1586364061
transform 1 0 2668 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_29
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 590 592
use scs8hd_buf_1  _120_
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__127__D
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_74
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_77
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_or4_4  _119_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__D
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use scs8hd_or3_4  _150_
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__C
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_124
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__C
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 406 592
use scs8hd_or3_4  _078_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_150
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  _086_
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_174
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_10_226
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_238
timestamp 1586364061
transform 1 0 23000 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_250
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_262
timestamp 1586364061
transform 1 0 25208 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_22
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_11_50
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_65
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 314 592
use scs8hd_or4_4  _127_
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_or4_4  _135_
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_or2_4  _071_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_130
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 406 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_or3_4  _067_
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_195
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_203
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_249
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_261
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_273
timestamp 1586364061
transform 1 0 26220 0 1 8160
box -38 -48 406 592
use scs8hd_conb_1  _175_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_17
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _068_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_nor4_4  _164_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_101
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_121
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 406 592
use scs8hd_or2_4  _095_
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_128
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_136
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_146
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__067__C
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_167
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_171
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_174
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_185
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_189
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_209
timestamp 1586364061
transform 1 0 20332 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_226
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_230
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_237
timestamp 1586364061
transform 1 0 22908 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_248
timestamp 1586364061
transform 1 0 23920 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_260
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_272
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_6
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_10
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_17
timestamp 1586364061
transform 1 0 2668 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_17
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_21
timestamp 1586364061
transform 1 0 3036 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_21
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _173_
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_32
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_28
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_47
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_61
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_69
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_conb_1  _180_
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_73
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__C
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_100
timestamp 1586364061
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _163_
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 1602 592
use scs8hd_or3_4  _109_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 406 592
use scs8hd_nor3_4  _159_
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1234 592
use scs8hd_nor3_4  _160_
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__159__C
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_139
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_146
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _083_
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_152
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 866 592
use scs8hd_or3_4  _085_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_171
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_187
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_183
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_196
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_193
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_203
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_199
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_218
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_222
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_226
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_230
timestamp 1586364061
transform 1 0 22264 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_235
timestamp 1586364061
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_243
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_248
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 22632 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_254
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_252
timestamp 1586364061
transform 1 0 24288 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_265
timestamp 1586364061
transform 1 0 25484 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_264
timestamp 1586364061
transform 1 0 25392 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_273
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_8
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_21
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_25
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_28
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_45
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_49
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 130 592
use scs8hd_buf_1  _151_
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_56
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_67
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _148_
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_84
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_or2_4  _074_
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 314 592
use scs8hd_or3_4  _082_
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_148
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _099_
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_161
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_165
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_169
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 18952 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_180
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_190
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_203
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_207
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_213
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_227
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_265
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_53
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_99
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_109
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_116
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_177
timestamp 1586364061
transform 1 0 17388 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 590 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_228
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23000 0 -1 11424
box -38 -48 866 592
use scs8hd_fill_2  FILLER_16_236
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24104 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_252
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_258
timestamp 1586364061
transform 1 0 24840 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_270
timestamp 1586364061
transform 1 0 25944 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_18
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_30
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_45
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_49
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_55
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_72
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_87
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_128
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_151
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_164
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_168
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_189
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 20608 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 20424 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_204
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_215
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_262
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_273
timestamp 1586364061
transform 1 0 26220 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4140 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_52
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_8  _147_
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_133
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_8  _144_
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_180
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_3  FILLER_18_188
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_209
timestamp 1586364061
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_229
timestamp 1586364061
transform 1 0 22172 0 -1 12512
box -38 -48 406 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 22908 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22540 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_235
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_240
timestamp 1586364061
transform 1 0 23184 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_244
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_247
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_17
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_21
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_41
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_37
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_45
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_96
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_100
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_135
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_155
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _143_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_167
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_171
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_179
timestamp 1586364061
transform 1 0 17572 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_195
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_189
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_218
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_222
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_228
timestamp 1586364061
transform 1 0 22080 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_239
timestamp 1586364061
transform 1 0 23092 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_235
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22540 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use scs8hd_conb_1  _176_
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_19_265
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_17
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_21
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_38
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_79
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_96
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_100
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_137
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_141
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_178
timestamp 1586364061
transform 1 0 17480 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_187
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_182
timestamp 1586364061
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_195
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_191
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_205
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_209
timestamp 1586364061
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_222
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_226
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_265
timestamp 1586364061
transform 1 0 25484 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_17
timestamp 1586364061
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4140 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_21
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_48
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_65
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_69
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_112
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 590 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 13524 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_127
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_131
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_168
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_185
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_189
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_232
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_235
timestamp 1586364061
transform 1 0 22724 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_248
timestamp 1586364061
transform 1 0 23920 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_252
timestamp 1586364061
transform 1 0 24288 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_265
timestamp 1586364061
transform 1 0 25484 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_273
timestamp 1586364061
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_6
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_10
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_14
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_25
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_29
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_44
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_48
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_96
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_100
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12512 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_139
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 406 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_146
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_169
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_173
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_177
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_190
timestamp 1586364061
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_194
timestamp 1586364061
transform 1 0 18952 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_209
timestamp 1586364061
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_213
timestamp 1586364061
transform 1 0 20700 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_217
timestamp 1586364061
transform 1 0 21068 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_235
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_239
timestamp 1586364061
transform 1 0 23092 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_265
timestamp 1586364061
transform 1 0 25484 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_18
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_22
timestamp 1586364061
transform 1 0 3128 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_28
timestamp 1586364061
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_45
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_58
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_75
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_79
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_6  FILLER_24_85
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_123
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_127
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_137
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 15456 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_158
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_170
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_193
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_197
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_201
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_224
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22908 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_232
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_246
timestamp 1586364061
transform 1 0 23736 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_250
timestamp 1586364061
transform 1 0 24104 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_254
timestamp 1586364061
transform 1 0 24472 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_258
timestamp 1586364061
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_270
timestamp 1586364061
transform 1 0 25944 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_56
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_97
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_142
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_146
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_188
timestamp 1586364061
transform 1 0 18400 0 1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_198
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_202
timestamp 1586364061
transform 1 0 19688 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_205
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_209
timestamp 1586364061
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 22264 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_222
timestamp 1586364061
transform 1 0 21528 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_226
timestamp 1586364061
transform 1 0 21896 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22724 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23092 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_233
timestamp 1586364061
transform 1 0 22540 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_237
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_241
timestamp 1586364061
transform 1 0 23276 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_248
timestamp 1586364061
transform 1 0 23920 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_252
timestamp 1586364061
transform 1 0 24288 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_259
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_263
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_267
timestamp 1586364061
transform 1 0 25668 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_275
timestamp 1586364061
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_26
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_22
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_28
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_45
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_45
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_49
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_52
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_66
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_100
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 10212 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_112
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_127
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_138
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_134
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_135
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_145
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_152
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_167
timestamp 1586364061
transform 1 0 16468 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_178
timestamp 1586364061
transform 1 0 17480 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_174
timestamp 1586364061
transform 1 0 17112 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_187
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_182
timestamp 1586364061
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_182
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_191
timestamp 1586364061
transform 1 0 18676 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_194
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_212
timestamp 1586364061
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_225
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_229
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_247
timestamp 1586364061
transform 1 0 23828 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_241
timestamp 1586364061
transform 1 0 23276 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_252
timestamp 1586364061
transform 1 0 24288 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_254
timestamp 1586364061
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_270
timestamp 1586364061
transform 1 0 25944 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_18
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_22
timestamp 1586364061
transform 1 0 3128 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_28
timestamp 1586364061
transform 1 0 3680 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_45
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_53
timestamp 1586364061
transform 1 0 5980 0 -1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6072 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_65
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_121
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_138
timestamp 1586364061
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_142
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15364 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_146
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17296 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_170
timestamp 1586364061
transform 1 0 16744 0 -1 17952
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_187
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_191
timestamp 1586364061
transform 1 0 18676 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_228
timestamp 1586364061
transform 1 0 22080 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_241
timestamp 1586364061
transform 1 0 23276 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _201_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_253
timestamp 1586364061
transform 1 0 24380 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_259
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_9
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_26
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_43
timestamp 1586364061
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_76
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_91
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_108
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_115
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_119
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_138
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_151
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _177_
timestamp 1586364061
transform 1 0 20056 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_200
timestamp 1586364061
transform 1 0 19504 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_205
timestamp 1586364061
transform 1 0 19964 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_209
timestamp 1586364061
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_213
timestamp 1586364061
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_226
timestamp 1586364061
transform 1 0 21896 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_230
timestamp 1586364061
transform 1 0 22264 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23092 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_238
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_241
timestamp 1586364061
transform 1 0 23276 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_253
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_259
timestamp 1586364061
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_263
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_275
timestamp 1586364061
transform 1 0 26404 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_22
timestamp 1586364061
transform 1 0 3128 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_49
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_53
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6716 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_57
timestamp 1586364061
transform 1 0 6348 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_70
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_81
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_85
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_96
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_101
timestamp 1586364061
transform 1 0 10396 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_116
timestamp 1586364061
transform 1 0 11776 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_122
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use scs8hd_buf_1  _110_
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_158
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  FILLER_30_161
timestamp 1586364061
transform 1 0 15916 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_173
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_194
timestamp 1586364061
transform 1 0 18952 0 -1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_200
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_12  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_236
timestamp 1586364061
transform 1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_242
timestamp 1586364061
transform 1 0 23368 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_254
timestamp 1586364061
transform 1 0 24472 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_266
timestamp 1586364061
transform 1 0 25576 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_274
timestamp 1586364061
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_18
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_22
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_26
timestamp 1586364061
transform 1 0 3496 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_48
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_60
timestamp 1586364061
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_65
timestamp 1586364061
transform 1 0 7084 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_69
timestamp 1586364061
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_73
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_79
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 406 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_91
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_31_106
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 774 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_131
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_138
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_144
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_155
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_172
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_176
timestamp 1586364061
transform 1 0 17296 0 1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_222
timestamp 1586364061
transform 1 0 21528 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_234
timestamp 1586364061
transform 1 0 22632 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_242
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_259
timestamp 1586364061
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_263
timestamp 1586364061
transform 1 0 25300 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_275
timestamp 1586364061
transform 1 0 26404 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_32_35
timestamp 1586364061
transform 1 0 4324 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_39
timestamp 1586364061
transform 1 0 4692 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_46
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_58
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_62
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_66
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_77
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_32_89
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_96
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_107
timestamp 1586364061
transform 1 0 10948 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_119
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_32_157
timestamp 1586364061
transform 1 0 15548 0 -1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_165
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_177
timestamp 1586364061
transform 1 0 17388 0 -1 20128
box -38 -48 590 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_32_183
timestamp 1586364061
transform 1 0 17940 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_193
timestamp 1586364061
transform 1 0 18860 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_204
timestamp 1586364061
transform 1 0 19872 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_208
timestamp 1586364061
transform 1 0 20240 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_22
timestamp 1586364061
transform 1 0 3128 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_18
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_30
timestamp 1586364061
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_29
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_18
timestamp 1586364061
transform 1 0 2760 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_33
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_45
timestamp 1586364061
transform 1 0 5244 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_99
timestamp 1586364061
transform 1 0 10212 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_111
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_158
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_170
timestamp 1586364061
transform 1 0 16744 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_182
timestamp 1586364061
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 25116 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_259
timestamp 1586364061
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_263
timestamp 1586364061
transform 1 0 25300 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_275
timestamp 1586364061
transform 1 0 26404 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_conb_1  _174_
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 314 592
use scs8hd_buf_2  _188_
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_11
timestamp 1586364061
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_18
timestamp 1586364061
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_22
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_46
timestamp 1586364061
transform 1 0 5336 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_58
timestamp 1586364061
transform 1 0 6440 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_259
timestamp 1586364061
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_263
timestamp 1586364061
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_275
timestamp 1586364061
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_6
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_36_17
timestamp 1586364061
transform 1 0 2668 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_29
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_43
timestamp 1586364061
transform 1 0 5060 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_37_55
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_37_115
timestamp 1586364061
transform 1 0 11684 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_153
timestamp 1586364061
transform 1 0 15180 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_168
timestamp 1586364061
transform 1 0 16560 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_180
timestamp 1586364061
transform 1 0 17664 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 23276 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_243
timestamp 1586364061
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 25116 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_259
timestamp 1586364061
transform 1 0 24932 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_263
timestamp 1586364061
transform 1 0 25300 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_275
timestamp 1586364061
transform 1 0 26404 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_116
timestamp 1586364061
transform 1 0 11776 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_128
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_152
timestamp 1586364061
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_157
timestamp 1586364061
transform 1 0 15548 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_169
timestamp 1586364061
transform 1 0 16652 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_181
timestamp 1586364061
transform 1 0 17756 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_193
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_205
timestamp 1586364061
transform 1 0 19964 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 23276 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_245
timestamp 1586364061
transform 1 0 23644 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_253
timestamp 1586364061
transform 1 0 24380 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_buf_2  _186_
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_7
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_126
timestamp 1586364061
transform 1 0 12696 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_130
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_138
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_165
timestamp 1586364061
transform 1 0 16284 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_174
timestamp 1586364061
transform 1 0 17112 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_178
timestamp 1586364061
transform 1 0 17480 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_181
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 17572 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_195
timestamp 1586364061
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_190
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 18676 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_195
timestamp 1586364061
transform 1 0 19044 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_183
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 19780 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 20332 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_199
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_207
timestamp 1586364061
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_211
timestamp 1586364061
transform 1 0 20516 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_207
timestamp 1586364061
transform 1 0 20148 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_229
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 23460 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 23828 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_233
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_241
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_247
timestamp 1586364061
transform 1 0 23828 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_259
timestamp 1586364061
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_271
timestamp 1586364061
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_253
timestamp 1586364061
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_259
timestamp 1586364061
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_263
timestamp 1586364061
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_275
timestamp 1586364061
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 4526 0 4582 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 7654 0 7710 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 10782 0 10838 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 13910 0 13966 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 16946 0 17002 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 20074 0 20130 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 23202 0 23258 480 6 address[6]
port 6 nsew default input
rlabel metal3 s 0 416 480 536 6 chanx_left_in[0]
port 7 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[1]
port 8 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[2]
port 9 nsew default input
rlabel metal3 s 0 3408 480 3528 6 chanx_left_in[3]
port 10 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[4]
port 11 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[5]
port 12 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[6]
port 13 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[7]
port 14 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[8]
port 15 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[0]
port 16 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[1]
port 17 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[2]
port 18 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[3]
port 19 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[4]
port 20 nsew default tristate
rlabel metal3 s 0 24216 480 24336 6 chanx_left_out[5]
port 21 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[6]
port 22 nsew default tristate
rlabel metal3 s 0 26256 480 26376 6 chanx_left_out[7]
port 23 nsew default tristate
rlabel metal3 s 0 27344 480 27464 6 chanx_left_out[8]
port 24 nsew default tristate
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_in[0]
port 25 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 chanx_right_in[1]
port 26 nsew default input
rlabel metal3 s 27520 3408 28000 3528 6 chanx_right_in[2]
port 27 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 chanx_right_in[3]
port 28 nsew default input
rlabel metal3 s 27520 5584 28000 5704 6 chanx_right_in[4]
port 29 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_in[5]
port 30 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[6]
port 31 nsew default input
rlabel metal3 s 27520 8712 28000 8832 6 chanx_right_in[7]
port 32 nsew default input
rlabel metal3 s 27520 9664 28000 9784 6 chanx_right_in[8]
port 33 nsew default input
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[0]
port 34 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[1]
port 35 nsew default tristate
rlabel metal3 s 27520 21088 28000 21208 6 chanx_right_out[2]
port 36 nsew default tristate
rlabel metal3 s 27520 22176 28000 22296 6 chanx_right_out[3]
port 37 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[4]
port 38 nsew default tristate
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_out[5]
port 39 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[6]
port 40 nsew default tristate
rlabel metal3 s 27520 26256 28000 26376 6 chanx_right_out[7]
port 41 nsew default tristate
rlabel metal3 s 27520 27344 28000 27464 6 chanx_right_out[8]
port 42 nsew default tristate
rlabel metal2 s 662 27520 718 28000 6 chany_top_in[0]
port 43 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 chany_top_in[1]
port 44 nsew default input
rlabel metal2 s 3422 27520 3478 28000 6 chany_top_in[2]
port 45 nsew default input
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[3]
port 46 nsew default input
rlabel metal2 s 6182 27520 6238 28000 6 chany_top_in[4]
port 47 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 48 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[6]
port 49 nsew default input
rlabel metal2 s 10414 27520 10470 28000 6 chany_top_in[7]
port 50 nsew default input
rlabel metal2 s 11794 27520 11850 28000 6 chany_top_in[8]
port 51 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_out[0]
port 52 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[1]
port 53 nsew default tristate
rlabel metal2 s 18786 27520 18842 28000 6 chany_top_out[2]
port 54 nsew default tristate
rlabel metal2 s 20166 27520 20222 28000 6 chany_top_out[3]
port 55 nsew default tristate
rlabel metal2 s 21638 27520 21694 28000 6 chany_top_out[4]
port 56 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[5]
port 57 nsew default tristate
rlabel metal2 s 24398 27520 24454 28000 6 chany_top_out[6]
port 58 nsew default tristate
rlabel metal2 s 25778 27520 25834 28000 6 chany_top_out[7]
port 59 nsew default tristate
rlabel metal2 s 27158 27520 27214 28000 6 chany_top_out[8]
port 60 nsew default tristate
rlabel metal2 s 26330 0 26386 480 6 data_in
port 61 nsew default input
rlabel metal2 s 1490 0 1546 480 6 enable
port 62 nsew default input
rlabel metal3 s 0 15920 480 16040 6 left_bottom_grid_pin_11_
port 63 nsew default input
rlabel metal3 s 0 17008 480 17128 6 left_bottom_grid_pin_13_
port 64 nsew default input
rlabel metal3 s 0 17960 480 18080 6 left_bottom_grid_pin_15_
port 65 nsew default input
rlabel metal3 s 0 10752 480 10872 6 left_bottom_grid_pin_1_
port 66 nsew default input
rlabel metal3 s 0 11704 480 11824 6 left_bottom_grid_pin_3_
port 67 nsew default input
rlabel metal3 s 0 12792 480 12912 6 left_bottom_grid_pin_5_
port 68 nsew default input
rlabel metal3 s 0 13880 480 14000 6 left_bottom_grid_pin_7_
port 69 nsew default input
rlabel metal3 s 0 14832 480 14952 6 left_bottom_grid_pin_9_
port 70 nsew default input
rlabel metal3 s 0 9664 480 9784 6 left_top_grid_pin_10_
port 71 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 right_bottom_grid_pin_11_
port 72 nsew default input
rlabel metal3 s 27520 17008 28000 17128 6 right_bottom_grid_pin_13_
port 73 nsew default input
rlabel metal3 s 27520 17960 28000 18080 6 right_bottom_grid_pin_15_
port 74 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 right_bottom_grid_pin_1_
port 75 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 right_bottom_grid_pin_3_
port 76 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 right_bottom_grid_pin_5_
port 77 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 right_bottom_grid_pin_7_
port 78 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 right_bottom_grid_pin_9_
port 79 nsew default input
rlabel metal3 s 27520 416 28000 536 6 right_top_grid_pin_10_
port 80 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 top_left_grid_pin_13_
port 81 nsew default input
rlabel metal2 s 14646 27520 14702 28000 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
