magic
tech sky130A
magscale 1 2
timestamp 1609022596
<< locali >>
rect 3433 11747 3467 11849
rect 3341 11543 3375 11713
rect 11989 9911 12023 10217
rect 3801 7259 3835 7429
rect 15853 7395 15887 7497
rect 18981 7055 19015 7701
rect 10793 6103 10827 6205
rect 4077 5695 4111 5797
rect 6837 5559 6871 5661
<< viali >>
rect 1869 14025 1903 14059
rect 2605 14025 2639 14059
rect 3341 14025 3375 14059
rect 3617 14025 3651 14059
rect 3801 14025 3835 14059
rect 3985 14025 4019 14059
rect 6561 14025 6595 14059
rect 2973 13957 3007 13991
rect 6193 13957 6227 13991
rect 7021 13889 7055 13923
rect 1685 13821 1719 13855
rect 2053 13821 2087 13855
rect 2421 13821 2455 13855
rect 2789 13821 2823 13855
rect 3157 13821 3191 13855
rect 6009 13821 6043 13855
rect 6377 13821 6411 13855
rect 6837 13821 6871 13855
rect 13645 13821 13679 13855
rect 14473 13821 14507 13855
rect 15209 13821 15243 13855
rect 15577 13821 15611 13855
rect 2237 13685 2271 13719
rect 13829 13685 13863 13719
rect 14657 13685 14691 13719
rect 15393 13685 15427 13719
rect 15761 13685 15795 13719
rect 2513 13413 2547 13447
rect 2145 13209 2179 13243
rect 2237 12937 2271 12971
rect 2881 12801 2915 12835
rect 3157 12801 3191 12835
rect 2697 12733 2731 12767
rect 2329 12597 2363 12631
rect 2789 12597 2823 12631
rect 3525 12597 3559 12631
rect 2145 12393 2179 12427
rect 2758 12325 2792 12359
rect 2053 12257 2087 12291
rect 6092 12257 6126 12291
rect 2237 12189 2271 12223
rect 2513 12189 2547 12223
rect 5825 12189 5859 12223
rect 1685 12053 1719 12087
rect 3893 12053 3927 12087
rect 7205 12053 7239 12087
rect 2329 11849 2363 11883
rect 3433 11849 3467 11883
rect 4905 11849 4939 11883
rect 8861 11849 8895 11883
rect 2145 11713 2179 11747
rect 2881 11713 2915 11747
rect 3249 11713 3283 11747
rect 3341 11713 3375 11747
rect 3433 11713 3467 11747
rect 3525 11713 3559 11747
rect 8401 11713 8435 11747
rect 1869 11645 1903 11679
rect 2697 11645 2731 11679
rect 3792 11645 3826 11679
rect 4997 11645 5031 11679
rect 5253 11645 5287 11679
rect 7757 11645 7791 11679
rect 1501 11509 1535 11543
rect 1961 11509 1995 11543
rect 2789 11509 2823 11543
rect 3341 11509 3375 11543
rect 6377 11509 6411 11543
rect 1869 11305 1903 11339
rect 2697 11305 2731 11339
rect 3157 11305 3191 11339
rect 3525 11305 3559 11339
rect 5641 11305 5675 11339
rect 6193 11305 6227 11339
rect 1777 11237 1811 11271
rect 7104 11237 7138 11271
rect 2237 11169 2271 11203
rect 3065 11169 3099 11203
rect 6101 11169 6135 11203
rect 6653 11169 6687 11203
rect 10333 11169 10367 11203
rect 10600 11169 10634 11203
rect 12541 11169 12575 11203
rect 12808 11169 12842 11203
rect 2329 11101 2363 11135
rect 2513 11101 2547 11135
rect 3341 11101 3375 11135
rect 5365 11101 5399 11135
rect 6377 11101 6411 11135
rect 6837 11101 6871 11135
rect 13921 11033 13955 11067
rect 5733 10965 5767 10999
rect 8217 10965 8251 10999
rect 11713 10965 11747 10999
rect 1501 10761 1535 10795
rect 6377 10761 6411 10795
rect 10517 10761 10551 10795
rect 8769 10693 8803 10727
rect 1961 10625 1995 10659
rect 2145 10625 2179 10659
rect 2329 10625 2363 10659
rect 5273 10625 5307 10659
rect 5917 10625 5951 10659
rect 6101 10625 6135 10659
rect 11253 10625 11287 10659
rect 12173 10625 12207 10659
rect 12541 10625 12575 10659
rect 13093 10625 13127 10659
rect 13277 10625 13311 10659
rect 13553 10625 13587 10659
rect 16865 10625 16899 10659
rect 7389 10557 7423 10591
rect 7656 10557 7690 10591
rect 8861 10557 8895 10591
rect 9128 10557 9162 10591
rect 13737 10557 13771 10591
rect 18061 10557 18095 10591
rect 18429 10557 18463 10591
rect 2596 10489 2630 10523
rect 4997 10489 5031 10523
rect 11069 10489 11103 10523
rect 11989 10489 12023 10523
rect 14004 10489 14038 10523
rect 17785 10489 17819 10523
rect 1869 10421 1903 10455
rect 3709 10421 3743 10455
rect 4629 10421 4663 10455
rect 5089 10421 5123 10455
rect 5457 10421 5491 10455
rect 5825 10421 5859 10455
rect 10241 10421 10275 10455
rect 10609 10421 10643 10455
rect 10977 10421 11011 10455
rect 11529 10421 11563 10455
rect 11897 10421 11931 10455
rect 12633 10421 12667 10455
rect 13001 10421 13035 10455
rect 15117 10421 15151 10455
rect 16313 10421 16347 10455
rect 16681 10421 16715 10455
rect 16773 10421 16807 10455
rect 17509 10421 17543 10455
rect 18245 10421 18279 10455
rect 2421 10217 2455 10251
rect 5457 10217 5491 10251
rect 6653 10217 6687 10251
rect 6745 10217 6779 10251
rect 7481 10217 7515 10251
rect 10241 10217 10275 10251
rect 10609 10217 10643 10251
rect 11069 10217 11103 10251
rect 11621 10217 11655 10251
rect 11805 10217 11839 10251
rect 11989 10217 12023 10251
rect 15117 10217 15151 10251
rect 16681 10217 16715 10251
rect 16957 10217 16991 10251
rect 17417 10217 17451 10251
rect 18153 10217 18187 10251
rect 1501 10149 1535 10183
rect 10149 10149 10183 10183
rect 10977 10149 11011 10183
rect 2789 10081 2823 10115
rect 4997 10081 5031 10115
rect 5825 10081 5859 10115
rect 7573 10081 7607 10115
rect 7840 10081 7874 10115
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 5089 10013 5123 10047
rect 5273 10013 5307 10047
rect 5917 10013 5951 10047
rect 6101 10013 6135 10047
rect 6929 10013 6963 10047
rect 7113 10013 7147 10047
rect 10425 10013 10459 10047
rect 11253 10013 11287 10047
rect 6285 9945 6319 9979
rect 14004 10149 14038 10183
rect 18245 10149 18279 10183
rect 12541 10081 12575 10115
rect 13737 10081 13771 10115
rect 15568 10081 15602 10115
rect 16865 10081 16899 10115
rect 17325 10081 17359 10115
rect 12633 10013 12667 10047
rect 12817 10013 12851 10047
rect 15301 10013 15335 10047
rect 17509 10013 17543 10047
rect 18337 10013 18371 10047
rect 17785 9945 17819 9979
rect 4629 9877 4663 9911
rect 8953 9877 8987 9911
rect 9781 9877 9815 9911
rect 11437 9877 11471 9911
rect 11989 9877 12023 9911
rect 12173 9877 12207 9911
rect 13461 9877 13495 9911
rect 2881 9673 2915 9707
rect 3709 9673 3743 9707
rect 12725 9673 12759 9707
rect 13553 9673 13587 9707
rect 17785 9673 17819 9707
rect 2513 9605 2547 9639
rect 4537 9605 4571 9639
rect 5825 9605 5859 9639
rect 6837 9605 6871 9639
rect 14841 9605 14875 9639
rect 16497 9605 16531 9639
rect 18245 9605 18279 9639
rect 3433 9537 3467 9571
rect 4261 9537 4295 9571
rect 4997 9537 5031 9571
rect 5181 9537 5215 9571
rect 6377 9537 6411 9571
rect 7389 9537 7423 9571
rect 8585 9537 8619 9571
rect 10333 9537 10367 9571
rect 10977 9537 11011 9571
rect 11897 9537 11931 9571
rect 13369 9537 13403 9571
rect 14105 9537 14139 9571
rect 15393 9537 15427 9571
rect 16313 9537 16347 9571
rect 17049 9537 17083 9571
rect 1685 9469 1719 9503
rect 2053 9469 2087 9503
rect 2789 9469 2823 9503
rect 3341 9469 3375 9503
rect 4905 9469 4939 9503
rect 5549 9469 5583 9503
rect 6193 9469 6227 9503
rect 7205 9469 7239 9503
rect 7757 9469 7791 9503
rect 10057 9469 10091 9503
rect 11713 9469 11747 9503
rect 11805 9469 11839 9503
rect 14013 9469 14047 9503
rect 15209 9469 15243 9503
rect 16957 9469 16991 9503
rect 18061 9469 18095 9503
rect 18429 9469 18463 9503
rect 1593 9401 1627 9435
rect 7297 9401 7331 9435
rect 9597 9401 9631 9435
rect 13093 9401 13127 9435
rect 14473 9401 14507 9435
rect 16037 9401 16071 9435
rect 16865 9401 16899 9435
rect 17509 9401 17543 9435
rect 1869 9333 1903 9367
rect 2237 9333 2271 9367
rect 3249 9333 3283 9367
rect 4077 9333 4111 9367
rect 4169 9333 4203 9367
rect 5365 9333 5399 9367
rect 5733 9333 5767 9367
rect 6285 9333 6319 9367
rect 9689 9333 9723 9367
rect 10149 9333 10183 9367
rect 11345 9333 11379 9367
rect 12541 9333 12575 9367
rect 13185 9333 13219 9367
rect 13921 9333 13955 9367
rect 14657 9333 14691 9367
rect 15301 9333 15335 9367
rect 15669 9333 15703 9367
rect 16129 9333 16163 9367
rect 17693 9333 17727 9367
rect 3249 9129 3283 9163
rect 3617 9129 3651 9163
rect 5825 9129 5859 9163
rect 6193 9129 6227 9163
rect 12817 9129 12851 9163
rect 13461 9129 13495 9163
rect 16589 9129 16623 9163
rect 17601 9129 17635 9163
rect 18061 9129 18095 9163
rect 3801 9061 3835 9095
rect 5641 9061 5675 9095
rect 6285 9061 6319 9095
rect 10149 9061 10183 9095
rect 16313 9061 16347 9095
rect 17233 9061 17267 9095
rect 17969 9061 18003 9095
rect 2136 8993 2170 9027
rect 4353 8993 4387 9027
rect 6745 8993 6779 9027
rect 7472 8993 7506 9027
rect 9137 8993 9171 9027
rect 10057 8993 10091 9027
rect 10609 8993 10643 9027
rect 10793 8993 10827 9027
rect 11244 8993 11278 9027
rect 12725 8993 12759 9027
rect 13369 8993 13403 9027
rect 13829 8993 13863 9027
rect 16129 8993 16163 9027
rect 17141 8993 17175 9027
rect 18429 8993 18463 9027
rect 1869 8925 1903 8959
rect 4537 8925 4571 8959
rect 4997 8925 5031 8959
rect 6377 8925 6411 8959
rect 6837 8925 6871 8959
rect 7205 8925 7239 8959
rect 9229 8925 9263 8959
rect 9413 8925 9447 8959
rect 10333 8925 10367 8959
rect 10977 8925 11011 8959
rect 13553 8925 13587 8959
rect 16037 8925 16071 8959
rect 17325 8925 17359 8959
rect 18153 8925 18187 8959
rect 13001 8857 13035 8891
rect 8585 8789 8619 8823
rect 8769 8789 8803 8823
rect 9689 8789 9723 8823
rect 12357 8789 12391 8823
rect 12541 8789 12575 8823
rect 16773 8789 16807 8823
rect 2881 8585 2915 8619
rect 3065 8585 3099 8619
rect 5365 8585 5399 8619
rect 13921 8585 13955 8619
rect 15945 8585 15979 8619
rect 3341 8517 3375 8551
rect 6377 8517 6411 8551
rect 13001 8517 13035 8551
rect 17785 8517 17819 8551
rect 18245 8517 18279 8551
rect 1501 8449 1535 8483
rect 6101 8449 6135 8483
rect 8217 8449 8251 8483
rect 10793 8449 10827 8483
rect 13553 8449 13587 8483
rect 14565 8449 14599 8483
rect 16497 8449 16531 8483
rect 16681 8449 16715 8483
rect 17325 8449 17359 8483
rect 3525 8381 3559 8415
rect 6561 8381 6595 8415
rect 7941 8381 7975 8415
rect 8401 8381 8435 8415
rect 10609 8381 10643 8415
rect 11161 8381 11195 8415
rect 13369 8381 13403 8415
rect 17141 8381 17175 8415
rect 17601 8381 17635 8415
rect 18061 8381 18095 8415
rect 18429 8381 18463 8415
rect 1768 8313 1802 8347
rect 3792 8313 3826 8347
rect 6009 8313 6043 8347
rect 8033 8313 8067 8347
rect 10149 8313 10183 8347
rect 12909 8313 12943 8347
rect 13461 8313 13495 8347
rect 14832 8313 14866 8347
rect 4905 8245 4939 8279
rect 5549 8245 5583 8279
rect 5917 8245 5951 8279
rect 6837 8245 6871 8279
rect 7573 8245 7607 8279
rect 10241 8245 10275 8279
rect 10701 8245 10735 8279
rect 16773 8245 16807 8279
rect 17233 8245 17267 8279
rect 2697 8041 2731 8075
rect 3065 8041 3099 8075
rect 3433 8041 3467 8075
rect 4537 8041 4571 8075
rect 4905 8041 4939 8075
rect 5365 8041 5399 8075
rect 7297 8041 7331 8075
rect 7849 8041 7883 8075
rect 8309 8041 8343 8075
rect 8677 8041 8711 8075
rect 8769 8041 8803 8075
rect 11621 8041 11655 8075
rect 12633 8041 12667 8075
rect 13829 8041 13863 8075
rect 16681 8041 16715 8075
rect 6000 7973 6034 8007
rect 7941 7973 7975 8007
rect 10486 7973 10520 8007
rect 12541 7973 12575 8007
rect 13369 7973 13403 8007
rect 17233 7973 17267 8007
rect 1685 7905 1719 7939
rect 2605 7905 2639 7939
rect 3525 7905 3559 7939
rect 4445 7905 4479 7939
rect 5273 7905 5307 7939
rect 5733 7905 5767 7939
rect 11897 7905 11931 7939
rect 12081 7905 12115 7939
rect 13461 7905 13495 7939
rect 15557 7905 15591 7939
rect 17141 7905 17175 7939
rect 17877 7905 17911 7939
rect 18245 7905 18279 7939
rect 2881 7837 2915 7871
rect 3709 7837 3743 7871
rect 4721 7837 4755 7871
rect 5457 7837 5491 7871
rect 8125 7837 8159 7871
rect 8861 7837 8895 7871
rect 10057 7837 10091 7871
rect 10241 7837 10275 7871
rect 12725 7837 12759 7871
rect 13553 7837 13587 7871
rect 15301 7837 15335 7871
rect 17325 7837 17359 7871
rect 16773 7769 16807 7803
rect 18061 7769 18095 7803
rect 1869 7701 1903 7735
rect 2053 7701 2087 7735
rect 2237 7701 2271 7735
rect 4077 7701 4111 7735
rect 7113 7701 7147 7735
rect 7481 7701 7515 7735
rect 11713 7701 11747 7735
rect 12173 7701 12207 7735
rect 13001 7701 13035 7735
rect 17601 7701 17635 7735
rect 18429 7701 18463 7735
rect 18981 7701 19015 7735
rect 2973 7497 3007 7531
rect 3893 7497 3927 7531
rect 5549 7497 5583 7531
rect 6469 7497 6503 7531
rect 9873 7497 9907 7531
rect 15209 7497 15243 7531
rect 15853 7497 15887 7531
rect 15945 7497 15979 7531
rect 16497 7497 16531 7531
rect 3801 7429 3835 7463
rect 6837 7429 6871 7463
rect 2421 7361 2455 7395
rect 2605 7361 2639 7395
rect 3617 7361 3651 7395
rect 1501 7293 1535 7327
rect 1593 7293 1627 7327
rect 2329 7293 2363 7327
rect 16313 7429 16347 7463
rect 18429 7429 18463 7463
rect 4537 7361 4571 7395
rect 5365 7361 5399 7395
rect 6101 7361 6135 7395
rect 6653 7361 6687 7395
rect 7389 7361 7423 7395
rect 8217 7361 8251 7395
rect 12081 7361 12115 7395
rect 12909 7361 12943 7395
rect 13001 7361 13035 7395
rect 15853 7361 15887 7395
rect 16957 7361 16991 7395
rect 17141 7361 17175 7395
rect 6009 7293 6043 7327
rect 7297 7293 7331 7327
rect 8493 7293 8527 7327
rect 8760 7293 8794 7327
rect 9965 7293 9999 7327
rect 10221 7293 10255 7327
rect 11897 7293 11931 7327
rect 13829 7293 13863 7327
rect 16129 7293 16163 7327
rect 17601 7293 17635 7327
rect 18061 7293 18095 7327
rect 3433 7225 3467 7259
rect 3801 7225 3835 7259
rect 4261 7225 4295 7259
rect 5089 7225 5123 7259
rect 11989 7225 12023 7259
rect 12817 7225 12851 7259
rect 14096 7225 14130 7259
rect 16865 7225 16899 7259
rect 17325 7225 17359 7259
rect 1777 7157 1811 7191
rect 1961 7157 1995 7191
rect 2789 7157 2823 7191
rect 3341 7157 3375 7191
rect 4353 7157 4387 7191
rect 4721 7157 4755 7191
rect 5181 7157 5215 7191
rect 5917 7157 5951 7191
rect 7205 7157 7239 7191
rect 7665 7157 7699 7191
rect 8033 7157 8067 7191
rect 8125 7157 8159 7191
rect 11345 7157 11379 7191
rect 11529 7157 11563 7191
rect 12449 7157 12483 7191
rect 13277 7157 13311 7191
rect 13645 7157 13679 7191
rect 17785 7157 17819 7191
rect 18245 7157 18279 7191
rect 18981 7021 19015 7055
rect 3341 6953 3375 6987
rect 4169 6953 4203 6987
rect 5641 6953 5675 6987
rect 5825 6953 5859 6987
rect 8125 6953 8159 6987
rect 13369 6953 13403 6987
rect 13461 6953 13495 6987
rect 13921 6953 13955 6987
rect 17969 6953 18003 6987
rect 18429 6953 18463 6987
rect 7021 6885 7055 6919
rect 14749 6885 14783 6919
rect 17233 6885 17267 6919
rect 1685 6817 1719 6851
rect 2053 6817 2087 6851
rect 2421 6817 2455 6851
rect 2789 6817 2823 6851
rect 3801 6817 3835 6851
rect 4528 6817 4562 6851
rect 6285 6817 6319 6851
rect 8033 6817 8067 6851
rect 8493 6817 8527 6851
rect 10784 6817 10818 6851
rect 12541 6817 12575 6851
rect 15301 6817 15335 6851
rect 15568 6817 15602 6851
rect 17141 6817 17175 6851
rect 4261 6749 4295 6783
rect 6377 6749 6411 6783
rect 6469 6749 6503 6783
rect 6745 6749 6779 6783
rect 8585 6749 8619 6783
rect 8769 6749 8803 6783
rect 8953 6749 8987 6783
rect 10517 6749 10551 6783
rect 11989 6749 12023 6783
rect 12633 6749 12667 6783
rect 12725 6749 12759 6783
rect 13553 6749 13587 6783
rect 14841 6749 14875 6783
rect 15025 6749 15059 6783
rect 17325 6749 17359 6783
rect 18061 6749 18095 6783
rect 18153 6749 18187 6783
rect 1593 6681 1627 6715
rect 2237 6681 2271 6715
rect 2605 6681 2639 6715
rect 2973 6681 3007 6715
rect 5917 6681 5951 6715
rect 14381 6681 14415 6715
rect 16681 6681 16715 6715
rect 16773 6681 16807 6715
rect 1869 6613 1903 6647
rect 3249 6613 3283 6647
rect 9229 6613 9263 6647
rect 11897 6613 11931 6647
rect 12173 6613 12207 6647
rect 13001 6613 13035 6647
rect 17601 6613 17635 6647
rect 1593 6409 1627 6443
rect 6653 6409 6687 6443
rect 8125 6409 8159 6443
rect 16865 6409 16899 6443
rect 17785 6409 17819 6443
rect 10149 6341 10183 6375
rect 15301 6341 15335 6375
rect 6285 6273 6319 6307
rect 6837 6273 6871 6307
rect 8769 6273 8803 6307
rect 9781 6273 9815 6307
rect 12909 6273 12943 6307
rect 13001 6273 13035 6307
rect 13369 6273 13403 6307
rect 13921 6273 13955 6307
rect 16589 6273 16623 6307
rect 17417 6273 17451 6307
rect 1685 6205 1719 6239
rect 2145 6205 2179 6239
rect 3617 6205 3651 6239
rect 8493 6205 8527 6239
rect 9505 6205 9539 6239
rect 10333 6205 10367 6239
rect 10793 6205 10827 6239
rect 10885 6205 10919 6239
rect 11152 6205 11186 6239
rect 12817 6205 12851 6239
rect 17325 6205 17359 6239
rect 18061 6205 18095 6239
rect 18429 6205 18463 6239
rect 2412 6137 2446 6171
rect 3862 6137 3896 6171
rect 5641 6137 5675 6171
rect 6193 6137 6227 6171
rect 8585 6137 8619 6171
rect 9045 6137 9079 6171
rect 14166 6137 14200 6171
rect 17233 6137 17267 6171
rect 1869 6069 1903 6103
rect 3525 6069 3559 6103
rect 4997 6069 5031 6103
rect 5733 6069 5767 6103
rect 6101 6069 6135 6103
rect 10793 6069 10827 6103
rect 12265 6069 12299 6103
rect 12449 6069 12483 6103
rect 15853 6069 15887 6103
rect 16037 6069 16071 6103
rect 16405 6069 16439 6103
rect 16497 6069 16531 6103
rect 18245 6069 18279 6103
rect 2605 5865 2639 5899
rect 3525 5865 3559 5899
rect 4169 5865 4203 5899
rect 4997 5865 5031 5899
rect 5365 5865 5399 5899
rect 5457 5865 5491 5899
rect 5825 5865 5859 5899
rect 7849 5865 7883 5899
rect 11069 5865 11103 5899
rect 11805 5865 11839 5899
rect 14197 5865 14231 5899
rect 15669 5865 15703 5899
rect 15853 5865 15887 5899
rect 16221 5865 16255 5899
rect 16681 5865 16715 5899
rect 17509 5865 17543 5899
rect 4077 5797 4111 5831
rect 4537 5797 4571 5831
rect 11713 5797 11747 5831
rect 1685 5729 1719 5763
rect 2053 5729 2087 5763
rect 3065 5729 3099 5763
rect 6009 5729 6043 5763
rect 7021 5729 7055 5763
rect 7389 5729 7423 5763
rect 9689 5729 9723 5763
rect 9956 5729 9990 5763
rect 13073 5729 13107 5763
rect 16313 5729 16347 5763
rect 17049 5729 17083 5763
rect 17693 5729 17727 5763
rect 17877 5729 17911 5763
rect 2513 5661 2547 5695
rect 3617 5661 3651 5695
rect 3801 5661 3835 5695
rect 4077 5661 4111 5695
rect 4629 5661 4663 5695
rect 4721 5661 4755 5695
rect 5549 5661 5583 5695
rect 6837 5661 6871 5695
rect 7757 5661 7791 5695
rect 11897 5661 11931 5695
rect 12817 5661 12851 5695
rect 16497 5661 16531 5695
rect 17141 5661 17175 5695
rect 17233 5661 17267 5695
rect 2881 5593 2915 5627
rect 18061 5593 18095 5627
rect 1869 5525 1903 5559
rect 2237 5525 2271 5559
rect 3157 5525 3191 5559
rect 6837 5525 6871 5559
rect 11345 5525 11379 5559
rect 18245 5525 18279 5559
rect 18429 5525 18463 5559
rect 4077 5321 4111 5355
rect 16221 5321 16255 5355
rect 16681 5321 16715 5355
rect 2605 5253 2639 5287
rect 6653 5253 6687 5287
rect 12449 5253 12483 5287
rect 18429 5253 18463 5287
rect 3709 5185 3743 5219
rect 3893 5185 3927 5219
rect 4721 5185 4755 5219
rect 5273 5185 5307 5219
rect 11253 5185 11287 5219
rect 12265 5185 12299 5219
rect 14289 5185 14323 5219
rect 16313 5185 16347 5219
rect 16589 5185 16623 5219
rect 17233 5185 17267 5219
rect 1593 5117 1627 5151
rect 2145 5117 2179 5151
rect 2697 5117 2731 5151
rect 3617 5117 3651 5151
rect 6837 5117 6871 5151
rect 7104 5117 7138 5151
rect 9229 5117 9263 5151
rect 17601 5117 17635 5151
rect 18061 5117 18095 5151
rect 1869 5049 1903 5083
rect 2973 5049 3007 5083
rect 4445 5049 4479 5083
rect 5518 5049 5552 5083
rect 9496 5049 9530 5083
rect 11345 5049 11379 5083
rect 13277 5049 13311 5083
rect 13369 5049 13403 5083
rect 17049 5049 17083 5083
rect 2329 4981 2363 5015
rect 3249 4981 3283 5015
rect 4537 4981 4571 5015
rect 8217 4981 8251 5015
rect 10609 4981 10643 5015
rect 14381 4981 14415 5015
rect 17141 4981 17175 5015
rect 17785 4981 17819 5015
rect 18245 4981 18279 5015
rect 2237 4777 2271 4811
rect 4537 4777 4571 4811
rect 4905 4777 4939 4811
rect 5365 4777 5399 4811
rect 5825 4777 5859 4811
rect 6193 4777 6227 4811
rect 9781 4777 9815 4811
rect 12081 4777 12115 4811
rect 13507 4777 13541 4811
rect 16589 4777 16623 4811
rect 16957 4777 16991 4811
rect 10508 4709 10542 4743
rect 12265 4709 12299 4743
rect 12366 4709 12400 4743
rect 15485 4709 15519 4743
rect 16405 4709 16439 4743
rect 17049 4709 17083 4743
rect 1685 4641 1719 4675
rect 4445 4641 4479 4675
rect 4997 4641 5031 4675
rect 5733 4641 5767 4675
rect 6561 4641 6595 4675
rect 8300 4641 8334 4675
rect 13404 4641 13438 4675
rect 14232 4641 14266 4675
rect 17417 4641 17451 4675
rect 17877 4641 17911 4675
rect 18245 4641 18279 4675
rect 5181 4573 5215 4607
rect 6009 4573 6043 4607
rect 8033 4573 8067 4607
rect 10241 4573 10275 4607
rect 13277 4573 13311 4607
rect 15393 4573 15427 4607
rect 17233 4573 17267 4607
rect 9413 4505 9447 4539
rect 17601 4505 17635 4539
rect 1869 4437 1903 4471
rect 2145 4437 2179 4471
rect 6377 4437 6411 4471
rect 11621 4437 11655 4471
rect 14335 4437 14369 4471
rect 15025 4437 15059 4471
rect 18061 4437 18095 4471
rect 18429 4437 18463 4471
rect 5365 4233 5399 4267
rect 6469 4233 6503 4267
rect 8493 4233 8527 4267
rect 2697 4165 2731 4199
rect 8585 4165 8619 4199
rect 9413 4165 9447 4199
rect 11989 4165 12023 4199
rect 1869 4097 1903 4131
rect 5917 4097 5951 4131
rect 6101 4097 6135 4131
rect 10977 4097 11011 4131
rect 12909 4097 12943 4131
rect 13369 4097 13403 4131
rect 14197 4097 14231 4131
rect 14841 4097 14875 4131
rect 16589 4097 16623 4131
rect 17233 4097 17267 4131
rect 1593 4029 1627 4063
rect 2145 4029 2179 4063
rect 2513 4029 2547 4063
rect 2973 4029 3007 4063
rect 3985 4029 4019 4063
rect 7113 4029 7147 4063
rect 8953 4029 8987 4063
rect 9781 4029 9815 4063
rect 10333 4029 10367 4063
rect 10701 4029 10735 4063
rect 11161 4029 11195 4063
rect 11529 4029 11563 4063
rect 12576 4029 12610 4063
rect 18061 4029 18095 4063
rect 18429 4029 18463 4063
rect 3065 3961 3099 3995
rect 4252 3961 4286 3995
rect 6285 3961 6319 3995
rect 7380 3961 7414 3995
rect 9321 3961 9355 3995
rect 11897 3961 11931 3995
rect 13001 3961 13035 3995
rect 14289 3961 14323 3995
rect 15393 3961 15427 3995
rect 15485 3961 15519 3995
rect 16405 3961 16439 3995
rect 16681 3961 16715 3995
rect 2329 3893 2363 3927
rect 5457 3893 5491 3927
rect 5825 3893 5859 3927
rect 6929 3893 6963 3927
rect 9873 3893 9907 3927
rect 12173 3893 12207 3927
rect 12679 3893 12713 3927
rect 17785 3893 17819 3927
rect 18245 3893 18279 3927
rect 2145 3689 2179 3723
rect 8033 3689 8067 3723
rect 9321 3689 9355 3723
rect 12081 3689 12115 3723
rect 12909 3689 12943 3723
rect 15853 3689 15887 3723
rect 16865 3689 16899 3723
rect 2329 3621 2363 3655
rect 5448 3621 5482 3655
rect 10692 3621 10726 3655
rect 1685 3553 1719 3587
rect 5181 3553 5215 3587
rect 6920 3553 6954 3587
rect 8493 3553 8527 3587
rect 8953 3553 8987 3587
rect 9873 3553 9907 3587
rect 10241 3553 10275 3587
rect 11897 3553 11931 3587
rect 12300 3553 12334 3587
rect 12608 3553 12642 3587
rect 13921 3553 13955 3587
rect 15025 3553 15059 3587
rect 15336 3553 15370 3587
rect 15439 3553 15473 3587
rect 15644 3553 15678 3587
rect 16313 3553 16347 3587
rect 16681 3553 16715 3587
rect 16957 3553 16991 3587
rect 17325 3553 17359 3587
rect 17877 3553 17911 3587
rect 18245 3553 18279 3587
rect 6653 3485 6687 3519
rect 8125 3485 8159 3519
rect 8861 3485 8895 3519
rect 10425 3485 10459 3519
rect 14841 3485 14875 3519
rect 1869 3417 1903 3451
rect 6561 3417 6595 3451
rect 9689 3417 9723 3451
rect 11805 3417 11839 3451
rect 14013 3417 14047 3451
rect 16037 3417 16071 3451
rect 17509 3417 17543 3451
rect 9137 3349 9171 3383
rect 10057 3349 10091 3383
rect 12403 3349 12437 3383
rect 12679 3349 12713 3383
rect 13645 3349 13679 3383
rect 15715 3349 15749 3383
rect 17141 3349 17175 3383
rect 17693 3349 17727 3383
rect 18061 3349 18095 3383
rect 18429 3349 18463 3383
rect 2973 3145 3007 3179
rect 8033 3145 8067 3179
rect 8125 3145 8159 3179
rect 2237 3077 2271 3111
rect 2605 3077 2639 3111
rect 2881 3077 2915 3111
rect 7021 3077 7055 3111
rect 7113 3077 7147 3111
rect 8493 3077 8527 3111
rect 15761 3077 15795 3111
rect 17417 3077 17451 3111
rect 8769 3009 8803 3043
rect 9597 3009 9631 3043
rect 11161 3009 11195 3043
rect 12173 3009 12207 3043
rect 16037 3009 16071 3043
rect 1685 2941 1719 2975
rect 2053 2941 2087 2975
rect 2421 2941 2455 2975
rect 7481 2941 7515 2975
rect 12449 2941 12483 2975
rect 15117 2941 15151 2975
rect 15577 2941 15611 2975
rect 17233 2941 17267 2975
rect 17601 2941 17635 2975
rect 18061 2941 18095 2975
rect 18429 2941 18463 2975
rect 7849 2873 7883 2907
rect 8861 2873 8895 2907
rect 9965 2873 9999 2907
rect 10057 2873 10091 2907
rect 10977 2873 11011 2907
rect 11253 2873 11287 2907
rect 12725 2873 12759 2907
rect 12817 2873 12851 2907
rect 13737 2873 13771 2907
rect 14013 2873 14047 2907
rect 14105 2873 14139 2907
rect 15025 2873 15059 2907
rect 16129 2873 16163 2907
rect 17049 2873 17083 2907
rect 1869 2805 1903 2839
rect 15301 2805 15335 2839
rect 17785 2805 17819 2839
rect 18245 2805 18279 2839
rect 3249 2601 3283 2635
rect 8309 2601 8343 2635
rect 8999 2601 9033 2635
rect 15163 2601 15197 2635
rect 5641 2533 5675 2567
rect 11345 2533 11379 2567
rect 12265 2533 12299 2567
rect 12817 2533 12851 2567
rect 14013 2533 14047 2567
rect 15669 2533 15703 2567
rect 18337 2533 18371 2567
rect 1593 2465 1627 2499
rect 2145 2465 2179 2499
rect 2789 2465 2823 2499
rect 3341 2465 3375 2499
rect 4077 2465 4111 2499
rect 5365 2465 5399 2499
rect 6469 2465 6503 2499
rect 6929 2465 6963 2499
rect 7297 2465 7331 2499
rect 7757 2465 7791 2499
rect 8125 2465 8159 2499
rect 8493 2465 8527 2499
rect 8896 2465 8930 2499
rect 9229 2465 9263 2499
rect 9965 2465 9999 2499
rect 10701 2465 10735 2499
rect 15060 2465 15094 2499
rect 16681 2465 16715 2499
rect 17049 2465 17083 2499
rect 17417 2465 17451 2499
rect 17785 2465 17819 2499
rect 1777 2397 1811 2431
rect 2329 2397 2363 2431
rect 3525 2397 3559 2431
rect 4261 2397 4295 2431
rect 7665 2397 7699 2431
rect 9781 2397 9815 2431
rect 10333 2397 10367 2431
rect 11253 2397 11287 2431
rect 12357 2397 12391 2431
rect 12725 2397 12759 2431
rect 13001 2397 13035 2431
rect 13921 2397 13955 2431
rect 14197 2397 14231 2431
rect 15577 2397 15611 2431
rect 15853 2397 15887 2431
rect 7941 2329 7975 2363
rect 8677 2329 8711 2363
rect 2973 2261 3007 2295
rect 6653 2261 6687 2295
rect 9413 2261 9447 2295
rect 10149 2261 10183 2295
rect 10793 2261 10827 2295
rect 16865 2261 16899 2295
rect 17233 2261 17267 2295
rect 17601 2261 17635 2295
rect 17969 2261 18003 2295
<< metal1 >>
rect 3326 15240 3332 15292
rect 3384 15280 3390 15292
rect 6178 15280 6184 15292
rect 3384 15252 6184 15280
rect 3384 15240 3390 15252
rect 6178 15240 6184 15252
rect 6236 15240 6242 15292
rect 3234 15172 3240 15224
rect 3292 15212 3298 15224
rect 6546 15212 6552 15224
rect 3292 15184 6552 15212
rect 3292 15172 3298 15184
rect 6546 15172 6552 15184
rect 6604 15172 6610 15224
rect 10962 15172 10968 15224
rect 11020 15212 11026 15224
rect 15838 15212 15844 15224
rect 11020 15184 15844 15212
rect 11020 15172 11026 15184
rect 15838 15172 15844 15184
rect 15896 15172 15902 15224
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 4062 14424 4068 14476
rect 4120 14464 4126 14476
rect 8478 14464 8484 14476
rect 4120 14436 8484 14464
rect 4120 14424 4126 14436
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 3326 14356 3332 14408
rect 3384 14396 3390 14408
rect 11790 14396 11796 14408
rect 3384 14368 11796 14396
rect 3384 14356 3390 14368
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 3786 14288 3792 14340
rect 3844 14328 3850 14340
rect 14182 14328 14188 14340
rect 3844 14300 14188 14328
rect 3844 14288 3850 14300
rect 14182 14288 14188 14300
rect 14240 14288 14246 14340
rect 14274 14288 14280 14340
rect 14332 14328 14338 14340
rect 19610 14328 19616 14340
rect 14332 14300 19616 14328
rect 14332 14288 14338 14300
rect 19610 14288 19616 14300
rect 19668 14288 19674 14340
rect 2406 14220 2412 14272
rect 2464 14260 2470 14272
rect 3602 14260 3608 14272
rect 2464 14232 3608 14260
rect 2464 14220 2470 14232
rect 3602 14220 3608 14232
rect 3660 14260 3666 14272
rect 12434 14260 12440 14272
rect 3660 14232 12440 14260
rect 3660 14220 3666 14232
rect 12434 14220 12440 14232
rect 12492 14260 12498 14272
rect 18322 14260 18328 14272
rect 12492 14232 18328 14260
rect 12492 14220 12498 14232
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 290 14016 296 14068
rect 348 14056 354 14068
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 348 14028 1869 14056
rect 348 14016 354 14028
rect 1857 14025 1869 14028
rect 1903 14025 1915 14059
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 1857 14019 1915 14025
rect 2148 14028 2605 14056
rect 1578 13948 1584 14000
rect 1636 13988 1642 14000
rect 2148 13988 2176 14028
rect 2593 14025 2605 14028
rect 2639 14025 2651 14059
rect 2593 14019 2651 14025
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 3329 14059 3387 14065
rect 3329 14056 3341 14059
rect 2924 14028 3341 14056
rect 2924 14016 2930 14028
rect 3329 14025 3341 14028
rect 3375 14025 3387 14059
rect 3602 14056 3608 14068
rect 3563 14028 3608 14056
rect 3329 14019 3387 14025
rect 3602 14016 3608 14028
rect 3660 14016 3666 14068
rect 3786 14056 3792 14068
rect 3747 14028 3792 14056
rect 3786 14016 3792 14028
rect 3844 14016 3850 14068
rect 3973 14059 4031 14065
rect 3973 14025 3985 14059
rect 4019 14056 4031 14059
rect 6549 14059 6607 14065
rect 4019 14028 6500 14056
rect 4019 14025 4031 14028
rect 3973 14019 4031 14025
rect 1636 13960 2176 13988
rect 1636 13948 1642 13960
rect 2222 13948 2228 14000
rect 2280 13988 2286 14000
rect 2961 13991 3019 13997
rect 2961 13988 2973 13991
rect 2280 13960 2973 13988
rect 2280 13948 2286 13960
rect 2961 13957 2973 13960
rect 3007 13957 3019 13991
rect 2961 13951 3019 13957
rect 934 13880 940 13932
rect 992 13920 998 13932
rect 3804 13920 3832 14016
rect 992 13892 2176 13920
rect 992 13880 998 13892
rect 1670 13852 1676 13864
rect 1631 13824 1676 13852
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 2038 13852 2044 13864
rect 1999 13824 2044 13852
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2148 13852 2176 13892
rect 2792 13892 3832 13920
rect 2406 13852 2412 13864
rect 2148 13824 2268 13852
rect 2367 13824 2412 13852
rect 2240 13725 2268 13824
rect 2406 13812 2412 13824
rect 2464 13812 2470 13864
rect 2792 13861 2820 13892
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13852 3203 13855
rect 3988 13852 4016 14019
rect 5994 13948 6000 14000
rect 6052 13988 6058 14000
rect 6181 13991 6239 13997
rect 6181 13988 6193 13991
rect 6052 13960 6193 13988
rect 6052 13948 6058 13960
rect 6181 13957 6193 13960
rect 6227 13957 6239 13991
rect 6472 13988 6500 14028
rect 6549 14025 6561 14059
rect 6595 14056 6607 14059
rect 6730 14056 6736 14068
rect 6595 14028 6736 14056
rect 6595 14025 6607 14028
rect 6549 14019 6607 14025
rect 6730 14016 6736 14028
rect 6788 14016 6794 14068
rect 6472 13960 7144 13988
rect 6181 13951 6239 13957
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 6104 13892 7021 13920
rect 6104 13864 6132 13892
rect 7009 13889 7021 13892
rect 7055 13889 7067 13923
rect 7116 13920 7144 13960
rect 10870 13948 10876 14000
rect 10928 13988 10934 14000
rect 15746 13988 15752 14000
rect 10928 13960 15752 13988
rect 10928 13948 10934 13960
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 13262 13920 13268 13932
rect 7116 13892 13268 13920
rect 7009 13883 7067 13889
rect 13262 13880 13268 13892
rect 13320 13920 13326 13932
rect 14274 13920 14280 13932
rect 13320 13892 14280 13920
rect 13320 13880 13326 13892
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 15654 13920 15660 13932
rect 15212 13892 15660 13920
rect 3191 13824 4016 13852
rect 5997 13855 6055 13861
rect 3191 13821 3203 13824
rect 3145 13815 3203 13821
rect 5997 13821 6009 13855
rect 6043 13852 6055 13855
rect 6086 13852 6092 13864
rect 6043 13824 6092 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 6270 13812 6276 13864
rect 6328 13852 6334 13864
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 6328 13824 6377 13852
rect 6328 13812 6334 13824
rect 6365 13821 6377 13824
rect 6411 13852 6423 13855
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6411 13824 6837 13852
rect 6411 13821 6423 13824
rect 6365 13815 6423 13821
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 13633 13855 13691 13861
rect 13633 13821 13645 13855
rect 13679 13852 13691 13855
rect 14366 13852 14372 13864
rect 13679 13824 14372 13852
rect 13679 13821 13691 13824
rect 13633 13815 13691 13821
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 15102 13852 15108 13864
rect 14507 13824 15108 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 15212 13861 15240 13892
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13821 15255 13855
rect 15562 13852 15568 13864
rect 15475 13824 15568 13852
rect 15197 13815 15255 13821
rect 15562 13812 15568 13824
rect 15620 13852 15626 13864
rect 16390 13852 16396 13864
rect 15620 13824 16396 13852
rect 15620 13812 15626 13824
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 4246 13744 4252 13796
rect 4304 13784 4310 13796
rect 4304 13756 14688 13784
rect 4304 13744 4310 13756
rect 2225 13719 2283 13725
rect 2225 13685 2237 13719
rect 2271 13685 2283 13719
rect 2225 13679 2283 13685
rect 8662 13676 8668 13728
rect 8720 13716 8726 13728
rect 10686 13716 10692 13728
rect 8720 13688 10692 13716
rect 8720 13676 8726 13688
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 13814 13716 13820 13728
rect 13775 13688 13820 13716
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 14660 13725 14688 13756
rect 14645 13719 14703 13725
rect 14645 13685 14657 13719
rect 14691 13685 14703 13719
rect 15378 13716 15384 13728
rect 15339 13688 15384 13716
rect 14645 13679 14703 13685
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 15470 13676 15476 13728
rect 15528 13716 15534 13728
rect 15749 13719 15807 13725
rect 15749 13716 15761 13719
rect 15528 13688 15761 13716
rect 15528 13676 15534 13688
rect 15749 13685 15761 13688
rect 15795 13685 15807 13719
rect 15749 13679 15807 13685
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 3326 13472 3332 13524
rect 3384 13512 3390 13524
rect 4430 13512 4436 13524
rect 3384 13484 4436 13512
rect 3384 13472 3390 13484
rect 4430 13472 4436 13484
rect 4488 13472 4494 13524
rect 9306 13472 9312 13524
rect 9364 13512 9370 13524
rect 11146 13512 11152 13524
rect 9364 13484 11152 13512
rect 9364 13472 9370 13484
rect 11146 13472 11152 13484
rect 11204 13472 11210 13524
rect 15378 13512 15384 13524
rect 11256 13484 15384 13512
rect 2038 13404 2044 13456
rect 2096 13444 2102 13456
rect 2501 13447 2559 13453
rect 2501 13444 2513 13447
rect 2096 13416 2513 13444
rect 2096 13404 2102 13416
rect 2501 13413 2513 13416
rect 2547 13444 2559 13447
rect 2547 13416 4752 13444
rect 2547 13413 2559 13416
rect 2501 13407 2559 13413
rect 4724 13376 4752 13416
rect 4798 13404 4804 13456
rect 4856 13444 4862 13456
rect 11256 13444 11284 13484
rect 15378 13472 15384 13484
rect 15436 13472 15442 13524
rect 4856 13416 11284 13444
rect 4856 13404 4862 13416
rect 13170 13404 13176 13456
rect 13228 13444 13234 13456
rect 14366 13444 14372 13456
rect 13228 13416 14372 13444
rect 13228 13404 13234 13416
rect 14366 13404 14372 13416
rect 14424 13404 14430 13456
rect 12250 13376 12256 13388
rect 4724 13348 12256 13376
rect 12250 13336 12256 13348
rect 12308 13376 12314 13388
rect 12308 13348 12480 13376
rect 12308 13336 12314 13348
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 12066 13308 12072 13320
rect 11296 13280 12072 13308
rect 11296 13268 11302 13280
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12452 13308 12480 13348
rect 12526 13336 12532 13388
rect 12584 13376 12590 13388
rect 14734 13376 14740 13388
rect 12584 13348 14740 13376
rect 12584 13336 12590 13348
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 17678 13376 17684 13388
rect 14844 13348 17684 13376
rect 14844 13308 14872 13348
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 12452 13280 14872 13308
rect 15654 13268 15660 13320
rect 15712 13308 15718 13320
rect 16390 13308 16396 13320
rect 15712 13280 16396 13308
rect 15712 13268 15718 13280
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 1670 13200 1676 13252
rect 1728 13240 1734 13252
rect 2133 13243 2191 13249
rect 2133 13240 2145 13243
rect 1728 13212 2145 13240
rect 1728 13200 1734 13212
rect 2133 13209 2145 13212
rect 2179 13240 2191 13243
rect 9398 13240 9404 13252
rect 2179 13212 9404 13240
rect 2179 13209 2191 13212
rect 2133 13203 2191 13209
rect 9398 13200 9404 13212
rect 9456 13240 9462 13252
rect 17034 13240 17040 13252
rect 9456 13212 17040 13240
rect 9456 13200 9462 13212
rect 17034 13200 17040 13212
rect 17092 13200 17098 13252
rect 10594 13132 10600 13184
rect 10652 13172 10658 13184
rect 14090 13172 14096 13184
rect 10652 13144 14096 13172
rect 10652 13132 10658 13144
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 14182 13132 14188 13184
rect 14240 13172 14246 13184
rect 18966 13172 18972 13184
rect 14240 13144 18972 13172
rect 14240 13132 14246 13144
rect 18966 13132 18972 13144
rect 19024 13132 19030 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 2774 12968 2780 12980
rect 2271 12940 2780 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 2774 12928 2780 12940
rect 2832 12968 2838 12980
rect 2832 12940 3004 12968
rect 2832 12928 2838 12940
rect 2498 12792 2504 12844
rect 2556 12832 2562 12844
rect 2869 12835 2927 12841
rect 2869 12832 2881 12835
rect 2556 12804 2881 12832
rect 2556 12792 2562 12804
rect 2869 12801 2881 12804
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12764 2743 12767
rect 2976 12764 3004 12940
rect 10226 12928 10232 12980
rect 10284 12968 10290 12980
rect 13446 12968 13452 12980
rect 10284 12940 13452 12968
rect 10284 12928 10290 12940
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 5442 12860 5448 12912
rect 5500 12900 5506 12912
rect 15470 12900 15476 12912
rect 5500 12872 15476 12900
rect 5500 12860 5506 12872
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 3142 12832 3148 12844
rect 3103 12804 3148 12832
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3510 12792 3516 12844
rect 3568 12832 3574 12844
rect 13814 12832 13820 12844
rect 3568 12804 13820 12832
rect 3568 12792 3574 12804
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 10778 12764 10784 12776
rect 2731 12736 10784 12764
rect 2731 12733 2743 12736
rect 2685 12727 2743 12733
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 11882 12764 11888 12776
rect 11296 12736 11888 12764
rect 11296 12724 11302 12736
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 2314 12628 2320 12640
rect 2275 12600 2320 12628
rect 2314 12588 2320 12600
rect 2372 12588 2378 12640
rect 2406 12588 2412 12640
rect 2464 12628 2470 12640
rect 2777 12631 2835 12637
rect 2777 12628 2789 12631
rect 2464 12600 2789 12628
rect 2464 12588 2470 12600
rect 2777 12597 2789 12600
rect 2823 12628 2835 12631
rect 3513 12631 3571 12637
rect 3513 12628 3525 12631
rect 2823 12600 3525 12628
rect 2823 12597 2835 12600
rect 2777 12591 2835 12597
rect 3513 12597 3525 12600
rect 3559 12628 3571 12631
rect 10870 12628 10876 12640
rect 3559 12600 10876 12628
rect 3559 12597 3571 12600
rect 3513 12591 3571 12597
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 2133 12427 2191 12433
rect 2133 12393 2145 12427
rect 2179 12424 2191 12427
rect 2314 12424 2320 12436
rect 2179 12396 2320 12424
rect 2179 12393 2191 12396
rect 2133 12387 2191 12393
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 7742 12424 7748 12436
rect 2424 12396 7748 12424
rect 2222 12316 2228 12368
rect 2280 12356 2286 12368
rect 2424 12356 2452 12396
rect 7742 12384 7748 12396
rect 7800 12424 7806 12436
rect 8018 12424 8024 12436
rect 7800 12396 8024 12424
rect 7800 12384 7806 12396
rect 8018 12384 8024 12396
rect 8076 12384 8082 12436
rect 13906 12384 13912 12436
rect 13964 12424 13970 12436
rect 14550 12424 14556 12436
rect 13964 12396 14556 12424
rect 13964 12384 13970 12396
rect 14550 12384 14556 12396
rect 14608 12384 14614 12436
rect 2280 12328 2452 12356
rect 2280 12316 2286 12328
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 2746 12359 2804 12365
rect 2746 12356 2758 12359
rect 2556 12328 2758 12356
rect 2556 12316 2562 12328
rect 2746 12325 2758 12328
rect 2792 12325 2804 12359
rect 2746 12319 2804 12325
rect 3234 12316 3240 12368
rect 3292 12356 3298 12368
rect 10962 12356 10968 12368
rect 3292 12328 10968 12356
rect 3292 12316 3298 12328
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12288 2099 12291
rect 2314 12288 2320 12300
rect 2087 12260 2320 12288
rect 2087 12257 2099 12260
rect 2041 12251 2099 12257
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 2590 12288 2596 12300
rect 2516 12260 2596 12288
rect 2516 12229 2544 12260
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 6080 12291 6138 12297
rect 6080 12257 6092 12291
rect 6126 12288 6138 12291
rect 6362 12288 6368 12300
rect 6126 12260 6368 12288
rect 6126 12257 6138 12260
rect 6080 12251 6138 12257
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12189 2559 12223
rect 2501 12183 2559 12189
rect 1673 12087 1731 12093
rect 1673 12053 1685 12087
rect 1719 12084 1731 12087
rect 1854 12084 1860 12096
rect 1719 12056 1860 12084
rect 1719 12053 1731 12056
rect 1673 12047 1731 12053
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 2240 12084 2268 12183
rect 4982 12180 4988 12232
rect 5040 12220 5046 12232
rect 5813 12223 5871 12229
rect 5813 12220 5825 12223
rect 5040 12192 5825 12220
rect 5040 12180 5046 12192
rect 5813 12189 5825 12192
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 3510 12112 3516 12164
rect 3568 12152 3574 12164
rect 16574 12152 16580 12164
rect 3568 12124 4016 12152
rect 3568 12112 3574 12124
rect 3786 12084 3792 12096
rect 2240 12056 3792 12084
rect 3786 12044 3792 12056
rect 3844 12084 3850 12096
rect 3881 12087 3939 12093
rect 3881 12084 3893 12087
rect 3844 12056 3893 12084
rect 3844 12044 3850 12056
rect 3881 12053 3893 12056
rect 3927 12053 3939 12087
rect 3988 12084 4016 12124
rect 6748 12124 16580 12152
rect 6748 12084 6776 12124
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 3988 12056 6776 12084
rect 7193 12087 7251 12093
rect 3881 12047 3939 12053
rect 7193 12053 7205 12087
rect 7239 12084 7251 12087
rect 7282 12084 7288 12096
rect 7239 12056 7288 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 2314 11880 2320 11892
rect 2275 11852 2320 11880
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 2682 11840 2688 11892
rect 2740 11880 2746 11892
rect 3421 11883 3479 11889
rect 3421 11880 3433 11883
rect 2740 11852 3433 11880
rect 2740 11840 2746 11852
rect 3421 11849 3433 11852
rect 3467 11849 3479 11883
rect 4893 11883 4951 11889
rect 4893 11880 4905 11883
rect 3421 11843 3479 11849
rect 3528 11852 4905 11880
rect 3528 11812 3556 11852
rect 4893 11849 4905 11852
rect 4939 11849 4951 11883
rect 4893 11843 4951 11849
rect 2148 11784 3556 11812
rect 2148 11753 2176 11784
rect 2133 11747 2191 11753
rect 2133 11713 2145 11747
rect 2179 11713 2191 11747
rect 2133 11707 2191 11713
rect 2498 11704 2504 11756
rect 2556 11744 2562 11756
rect 2869 11747 2927 11753
rect 2869 11744 2881 11747
rect 2556 11716 2881 11744
rect 2556 11704 2562 11716
rect 2869 11713 2881 11716
rect 2915 11713 2927 11747
rect 3234 11744 3240 11756
rect 3195 11716 3240 11744
rect 2869 11707 2927 11713
rect 3234 11704 3240 11716
rect 3292 11744 3298 11756
rect 3329 11747 3387 11753
rect 3329 11744 3341 11747
rect 3292 11716 3341 11744
rect 3292 11704 3298 11716
rect 3329 11713 3341 11716
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11744 3479 11747
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 3467 11716 3525 11744
rect 3467 11713 3479 11716
rect 3421 11707 3479 11713
rect 3513 11713 3525 11716
rect 3559 11713 3571 11747
rect 4908 11744 4936 11843
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 7800 11852 8861 11880
rect 7800 11840 7806 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 15562 11840 15568 11892
rect 15620 11880 15626 11892
rect 16206 11880 16212 11892
rect 15620 11852 16212 11880
rect 15620 11840 15626 11852
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 8386 11744 8392 11756
rect 4908 11716 5120 11744
rect 8347 11716 8392 11744
rect 3513 11707 3571 11713
rect 1854 11676 1860 11688
rect 1815 11648 1860 11676
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 3142 11676 3148 11688
rect 2731 11648 3148 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 3234 11568 3240 11620
rect 3292 11608 3298 11620
rect 3528 11608 3556 11707
rect 3786 11685 3792 11688
rect 3780 11676 3792 11685
rect 3747 11648 3792 11676
rect 3780 11639 3792 11648
rect 3786 11636 3792 11639
rect 3844 11636 3850 11688
rect 4982 11676 4988 11688
rect 4724 11648 4988 11676
rect 4724 11608 4752 11648
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 5092 11676 5120 11716
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 5241 11679 5299 11685
rect 5241 11676 5253 11679
rect 5092 11648 5253 11676
rect 5241 11645 5253 11648
rect 5287 11645 5299 11679
rect 7742 11676 7748 11688
rect 7703 11648 7748 11676
rect 5241 11639 5299 11645
rect 7742 11636 7748 11648
rect 7800 11636 7806 11688
rect 14642 11676 14648 11688
rect 7852 11648 14648 11676
rect 7852 11608 7880 11648
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 3292 11580 3464 11608
rect 3528 11580 4752 11608
rect 4816 11580 7880 11608
rect 3292 11568 3298 11580
rect 1489 11543 1547 11549
rect 1489 11509 1501 11543
rect 1535 11540 1547 11543
rect 1670 11540 1676 11552
rect 1535 11512 1676 11540
rect 1535 11509 1547 11512
rect 1489 11503 1547 11509
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 1949 11543 2007 11549
rect 1949 11540 1961 11543
rect 1912 11512 1961 11540
rect 1912 11500 1918 11512
rect 1949 11509 1961 11512
rect 1995 11509 2007 11543
rect 1949 11503 2007 11509
rect 2590 11500 2596 11552
rect 2648 11540 2654 11552
rect 2777 11543 2835 11549
rect 2777 11540 2789 11543
rect 2648 11512 2789 11540
rect 2648 11500 2654 11512
rect 2777 11509 2789 11512
rect 2823 11540 2835 11543
rect 3329 11543 3387 11549
rect 3329 11540 3341 11543
rect 2823 11512 3341 11540
rect 2823 11509 2835 11512
rect 2777 11503 2835 11509
rect 3329 11509 3341 11512
rect 3375 11509 3387 11543
rect 3436 11540 3464 11580
rect 4816 11540 4844 11580
rect 6362 11540 6368 11552
rect 3436 11512 4844 11540
rect 6323 11512 6368 11540
rect 3329 11503 3387 11509
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 2685 11339 2743 11345
rect 2685 11336 2697 11339
rect 2004 11308 2697 11336
rect 2004 11296 2010 11308
rect 2685 11305 2697 11308
rect 2731 11305 2743 11339
rect 3145 11339 3203 11345
rect 3145 11336 3157 11339
rect 2685 11299 2743 11305
rect 2884 11308 3157 11336
rect 1578 11228 1584 11280
rect 1636 11268 1642 11280
rect 1765 11271 1823 11277
rect 1765 11268 1777 11271
rect 1636 11240 1777 11268
rect 1636 11228 1642 11240
rect 1765 11237 1777 11240
rect 1811 11268 1823 11271
rect 2884 11268 2912 11308
rect 3145 11305 3157 11308
rect 3191 11336 3203 11339
rect 3234 11336 3240 11348
rect 3191 11308 3240 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 3510 11336 3516 11348
rect 3471 11308 3516 11336
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 3694 11296 3700 11348
rect 3752 11336 3758 11348
rect 5629 11339 5687 11345
rect 5629 11336 5641 11339
rect 3752 11308 5641 11336
rect 3752 11296 3758 11308
rect 5629 11305 5641 11308
rect 5675 11336 5687 11339
rect 6181 11339 6239 11345
rect 6181 11336 6193 11339
rect 5675 11308 6193 11336
rect 5675 11305 5687 11308
rect 5629 11299 5687 11305
rect 6181 11305 6193 11308
rect 6227 11336 6239 11339
rect 17310 11336 17316 11348
rect 6227 11308 17316 11336
rect 6227 11305 6239 11308
rect 6181 11299 6239 11305
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 3786 11268 3792 11280
rect 1811 11240 2912 11268
rect 2976 11240 3792 11268
rect 1811 11237 1823 11240
rect 1765 11231 1823 11237
rect 2222 11200 2228 11212
rect 2183 11172 2228 11200
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11132 2559 11135
rect 2976 11132 3004 11240
rect 3786 11228 3792 11240
rect 3844 11228 3850 11280
rect 4982 11228 4988 11280
rect 5040 11268 5046 11280
rect 6822 11268 6828 11280
rect 5040 11240 6828 11268
rect 5040 11228 5046 11240
rect 6822 11228 6828 11240
rect 6880 11228 6886 11280
rect 7092 11271 7150 11277
rect 7092 11237 7104 11271
rect 7138 11268 7150 11271
rect 7282 11268 7288 11280
rect 7138 11240 7288 11268
rect 7138 11237 7150 11240
rect 7092 11231 7150 11237
rect 7282 11228 7288 11240
rect 7340 11228 7346 11280
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11200 3111 11203
rect 3510 11200 3516 11212
rect 3099 11172 3516 11200
rect 3099 11169 3111 11172
rect 3053 11163 3111 11169
rect 2547 11104 3004 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 3068 11064 3096 11163
rect 3510 11160 3516 11172
rect 3568 11160 3574 11212
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11200 6147 11203
rect 6638 11200 6644 11212
rect 6135 11172 6644 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 10410 11200 10416 11212
rect 10367 11172 10416 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 10588 11203 10646 11209
rect 10588 11169 10600 11203
rect 10634 11200 10646 11203
rect 11330 11200 11336 11212
rect 10634 11172 11336 11200
rect 10634 11169 10646 11172
rect 10588 11163 10646 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11200 12587 11203
rect 12618 11200 12624 11212
rect 12575 11172 12624 11200
rect 12575 11169 12587 11172
rect 12529 11163 12587 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 12796 11203 12854 11209
rect 12796 11169 12808 11203
rect 12842 11200 12854 11203
rect 13262 11200 13268 11212
rect 12842 11172 13268 11200
rect 12842 11169 12854 11172
rect 12796 11163 12854 11169
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 3329 11135 3387 11141
rect 3329 11132 3341 11135
rect 3252 11104 3341 11132
rect 3252 11076 3280 11104
rect 3329 11101 3341 11104
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 5353 11135 5411 11141
rect 5353 11132 5365 11135
rect 4396 11104 5365 11132
rect 4396 11092 4402 11104
rect 5353 11101 5365 11104
rect 5399 11132 5411 11135
rect 5902 11132 5908 11144
rect 5399 11104 5908 11132
rect 5399 11101 5411 11104
rect 5353 11095 5411 11101
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 6362 11132 6368 11144
rect 6323 11104 6368 11132
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 6822 11132 6828 11144
rect 6783 11104 6828 11132
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 11624 11104 12572 11132
rect 2832 11036 3096 11064
rect 2832 11024 2838 11036
rect 3234 11024 3240 11076
rect 3292 11024 3298 11076
rect 3418 11024 3424 11076
rect 3476 11064 3482 11076
rect 6086 11064 6092 11076
rect 3476 11036 6092 11064
rect 3476 11024 3482 11036
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 5718 10996 5724 11008
rect 5679 10968 5724 10996
rect 5718 10956 5724 10968
rect 5776 10956 5782 11008
rect 8202 10996 8208 11008
rect 8163 10968 8208 10996
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 11624 10996 11652 11104
rect 8352 10968 11652 10996
rect 11701 10999 11759 11005
rect 8352 10956 8358 10968
rect 11701 10965 11713 10999
rect 11747 10996 11759 10999
rect 11882 10996 11888 11008
rect 11747 10968 11888 10996
rect 11747 10965 11759 10968
rect 11701 10959 11759 10965
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 12544 10996 12572 11104
rect 13538 11092 13544 11144
rect 13596 11132 13602 11144
rect 15194 11132 15200 11144
rect 13596 11104 15200 11132
rect 13596 11092 13602 11104
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 13630 11024 13636 11076
rect 13688 11064 13694 11076
rect 13909 11067 13967 11073
rect 13909 11064 13921 11067
rect 13688 11036 13921 11064
rect 13688 11024 13694 11036
rect 13909 11033 13921 11036
rect 13955 11033 13967 11067
rect 13909 11027 13967 11033
rect 16114 11024 16120 11076
rect 16172 11064 16178 11076
rect 17770 11064 17776 11076
rect 16172 11036 17776 11064
rect 16172 11024 16178 11036
rect 17770 11024 17776 11036
rect 17828 11024 17834 11076
rect 16298 10996 16304 11008
rect 12544 10968 16304 10996
rect 16298 10956 16304 10968
rect 16356 10956 16362 11008
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 1489 10795 1547 10801
rect 1489 10761 1501 10795
rect 1535 10792 1547 10795
rect 2222 10792 2228 10804
rect 1535 10764 2228 10792
rect 1535 10761 1547 10764
rect 1489 10755 1547 10761
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 2682 10792 2688 10804
rect 2332 10764 2688 10792
rect 1762 10684 1768 10736
rect 1820 10724 1826 10736
rect 2332 10724 2360 10764
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 3786 10792 3792 10804
rect 3108 10764 3792 10792
rect 3108 10752 3114 10764
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 6178 10752 6184 10804
rect 6236 10792 6242 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 6236 10764 6377 10792
rect 6236 10752 6242 10764
rect 6365 10761 6377 10764
rect 6411 10792 6423 10795
rect 6638 10792 6644 10804
rect 6411 10764 6644 10792
rect 6411 10761 6423 10764
rect 6365 10755 6423 10761
rect 6638 10752 6644 10764
rect 6696 10792 6702 10804
rect 10505 10795 10563 10801
rect 6696 10764 10456 10792
rect 6696 10752 6702 10764
rect 8754 10724 8760 10736
rect 1820 10696 2360 10724
rect 8715 10696 8760 10724
rect 1820 10684 1826 10696
rect 1946 10656 1952 10668
rect 1907 10628 1952 10656
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 2332 10665 2360 10696
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10625 2191 10659
rect 2133 10619 2191 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 5258 10656 5264 10668
rect 5171 10628 5264 10656
rect 2317 10619 2375 10625
rect 1854 10452 1860 10464
rect 1815 10424 1860 10452
rect 1854 10412 1860 10424
rect 1912 10412 1918 10464
rect 2148 10452 2176 10619
rect 5258 10616 5264 10628
rect 5316 10656 5322 10668
rect 5316 10628 5672 10656
rect 5316 10616 5322 10628
rect 2584 10523 2642 10529
rect 2584 10489 2596 10523
rect 2630 10520 2642 10523
rect 3234 10520 3240 10532
rect 2630 10492 3240 10520
rect 2630 10489 2642 10492
rect 2584 10483 2642 10489
rect 3234 10480 3240 10492
rect 3292 10480 3298 10532
rect 4062 10480 4068 10532
rect 4120 10520 4126 10532
rect 4890 10520 4896 10532
rect 4120 10492 4896 10520
rect 4120 10480 4126 10492
rect 4890 10480 4896 10492
rect 4948 10480 4954 10532
rect 4985 10523 5043 10529
rect 4985 10489 4997 10523
rect 5031 10520 5043 10523
rect 5644 10520 5672 10628
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 5905 10659 5963 10665
rect 5905 10656 5917 10659
rect 5776 10628 5917 10656
rect 5776 10616 5782 10628
rect 5905 10625 5917 10628
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 6089 10659 6147 10665
rect 6089 10625 6101 10659
rect 6135 10656 6147 10659
rect 6178 10656 6184 10668
rect 6135 10628 6184 10656
rect 6135 10625 6147 10628
rect 6089 10619 6147 10625
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 10428 10656 10456 10764
rect 10505 10761 10517 10795
rect 10551 10792 10563 10795
rect 10778 10792 10784 10804
rect 10551 10764 10784 10792
rect 10551 10761 10563 10764
rect 10505 10755 10563 10761
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 18046 10792 18052 10804
rect 10980 10764 18052 10792
rect 10980 10656 11008 10764
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 13630 10724 13636 10736
rect 12176 10696 13636 10724
rect 10428 10628 11008 10656
rect 11241 10659 11299 10665
rect 11241 10625 11253 10659
rect 11287 10656 11299 10659
rect 11330 10656 11336 10668
rect 11287 10628 11336 10656
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 11330 10616 11336 10628
rect 11388 10656 11394 10668
rect 12176 10665 12204 10696
rect 13630 10684 13636 10696
rect 13688 10684 13694 10736
rect 12161 10659 12219 10665
rect 12161 10656 12173 10659
rect 11388 10628 12173 10656
rect 11388 10616 11394 10628
rect 12161 10625 12173 10628
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 12710 10656 12716 10668
rect 12575 10628 12716 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 12710 10616 12716 10628
rect 12768 10656 12774 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 12768 10628 13093 10656
rect 12768 10616 12774 10628
rect 13081 10625 13093 10628
rect 13127 10625 13139 10659
rect 13262 10656 13268 10668
rect 13223 10628 13268 10656
rect 13081 10619 13139 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 13538 10656 13544 10668
rect 13499 10628 13544 10656
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 16632 10628 16865 10656
rect 16632 10616 16638 10628
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7374 10588 7380 10600
rect 6880 10560 7380 10588
rect 6880 10548 6886 10560
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 7644 10591 7702 10597
rect 7644 10557 7656 10591
rect 7690 10588 7702 10591
rect 8202 10588 8208 10600
rect 7690 10560 8208 10588
rect 7690 10557 7702 10560
rect 7644 10551 7702 10557
rect 7659 10520 7687 10551
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 9116 10591 9174 10597
rect 9116 10557 9128 10591
rect 9162 10588 9174 10591
rect 11882 10588 11888 10600
rect 9162 10560 11888 10588
rect 9162 10557 9174 10560
rect 9116 10551 9174 10557
rect 5031 10492 5488 10520
rect 5644 10492 7687 10520
rect 8864 10520 8892 10551
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 13725 10591 13783 10597
rect 13725 10588 13737 10591
rect 12676 10560 13737 10588
rect 12676 10548 12682 10560
rect 13725 10557 13737 10560
rect 13771 10588 13783 10591
rect 13814 10588 13820 10600
rect 13771 10560 13820 10588
rect 13771 10557 13783 10560
rect 13725 10551 13783 10557
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 14976 10560 18061 10588
rect 14976 10548 14982 10560
rect 18049 10557 18061 10560
rect 18095 10588 18107 10591
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 18095 10560 18429 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18417 10557 18429 10560
rect 18463 10557 18475 10591
rect 18417 10551 18475 10557
rect 10410 10520 10416 10532
rect 8864 10492 10416 10520
rect 5031 10489 5043 10492
rect 4985 10483 5043 10489
rect 2498 10452 2504 10464
rect 2148 10424 2504 10452
rect 2498 10412 2504 10424
rect 2556 10452 2562 10464
rect 3050 10452 3056 10464
rect 2556 10424 3056 10452
rect 2556 10412 2562 10424
rect 3050 10412 3056 10424
rect 3108 10452 3114 10464
rect 3697 10455 3755 10461
rect 3697 10452 3709 10455
rect 3108 10424 3709 10452
rect 3108 10412 3114 10424
rect 3697 10421 3709 10424
rect 3743 10421 3755 10455
rect 3697 10415 3755 10421
rect 4617 10455 4675 10461
rect 4617 10421 4629 10455
rect 4663 10452 4675 10455
rect 4798 10452 4804 10464
rect 4663 10424 4804 10452
rect 4663 10421 4675 10424
rect 4617 10415 4675 10421
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5074 10452 5080 10464
rect 5035 10424 5080 10452
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5460 10461 5488 10492
rect 10410 10480 10416 10492
rect 10468 10480 10474 10532
rect 11054 10520 11060 10532
rect 10967 10492 11060 10520
rect 11054 10480 11060 10492
rect 11112 10520 11118 10532
rect 11698 10520 11704 10532
rect 11112 10492 11704 10520
rect 11112 10480 11118 10492
rect 11698 10480 11704 10492
rect 11756 10480 11762 10532
rect 11977 10523 12035 10529
rect 11977 10489 11989 10523
rect 12023 10520 12035 10523
rect 12023 10492 12664 10520
rect 12023 10489 12035 10492
rect 11977 10483 12035 10489
rect 5445 10455 5503 10461
rect 5445 10421 5457 10455
rect 5491 10421 5503 10455
rect 5445 10415 5503 10421
rect 5813 10455 5871 10461
rect 5813 10421 5825 10455
rect 5859 10452 5871 10455
rect 5902 10452 5908 10464
rect 5859 10424 5908 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 10134 10452 10140 10464
rect 7524 10424 10140 10452
rect 7524 10412 7530 10424
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 10229 10455 10287 10461
rect 10229 10421 10241 10455
rect 10275 10452 10287 10455
rect 10318 10452 10324 10464
rect 10275 10424 10324 10452
rect 10275 10421 10287 10424
rect 10229 10415 10287 10421
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 10597 10455 10655 10461
rect 10597 10452 10609 10455
rect 10560 10424 10609 10452
rect 10560 10412 10566 10424
rect 10597 10421 10609 10424
rect 10643 10421 10655 10455
rect 10962 10452 10968 10464
rect 10923 10424 10968 10452
rect 10597 10415 10655 10421
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 11885 10455 11943 10461
rect 11885 10421 11897 10455
rect 11931 10452 11943 10455
rect 12158 10452 12164 10464
rect 11931 10424 12164 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 12636 10461 12664 10492
rect 13262 10480 13268 10532
rect 13320 10520 13326 10532
rect 13992 10523 14050 10529
rect 13320 10492 13768 10520
rect 13320 10480 13326 10492
rect 13740 10464 13768 10492
rect 13992 10489 14004 10523
rect 14038 10520 14050 10523
rect 15010 10520 15016 10532
rect 14038 10492 15016 10520
rect 14038 10489 14050 10492
rect 13992 10483 14050 10489
rect 15010 10480 15016 10492
rect 15068 10480 15074 10532
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 17770 10520 17776 10532
rect 15620 10492 17776 10520
rect 15620 10480 15626 10492
rect 17770 10480 17776 10492
rect 17828 10480 17834 10532
rect 12621 10455 12679 10461
rect 12621 10421 12633 10455
rect 12667 10421 12679 10455
rect 12621 10415 12679 10421
rect 12989 10455 13047 10461
rect 12989 10421 13001 10455
rect 13035 10452 13047 10455
rect 13354 10452 13360 10464
rect 13035 10424 13360 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 13354 10412 13360 10424
rect 13412 10452 13418 10464
rect 13538 10452 13544 10464
rect 13412 10424 13544 10452
rect 13412 10412 13418 10424
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 15105 10455 15163 10461
rect 15105 10452 15117 10455
rect 13780 10424 15117 10452
rect 13780 10412 13786 10424
rect 15105 10421 15117 10424
rect 15151 10421 15163 10455
rect 16298 10452 16304 10464
rect 16259 10424 16304 10452
rect 15105 10415 15163 10421
rect 16298 10412 16304 10424
rect 16356 10412 16362 10464
rect 16666 10452 16672 10464
rect 16627 10424 16672 10452
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 16761 10455 16819 10461
rect 16761 10421 16773 10455
rect 16807 10452 16819 10455
rect 16942 10452 16948 10464
rect 16807 10424 16948 10452
rect 16807 10421 16819 10424
rect 16761 10415 16819 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 17494 10452 17500 10464
rect 17455 10424 17500 10452
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 18233 10455 18291 10461
rect 18233 10421 18245 10455
rect 18279 10452 18291 10455
rect 18322 10452 18328 10464
rect 18279 10424 18328 10452
rect 18279 10421 18291 10424
rect 18233 10415 18291 10421
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 2314 10208 2320 10260
rect 2372 10248 2378 10260
rect 2409 10251 2467 10257
rect 2409 10248 2421 10251
rect 2372 10220 2421 10248
rect 2372 10208 2378 10220
rect 2409 10217 2421 10220
rect 2455 10217 2467 10251
rect 2409 10211 2467 10217
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4120 10220 5028 10248
rect 4120 10208 4126 10220
rect 1489 10183 1547 10189
rect 1489 10149 1501 10183
rect 1535 10180 1547 10183
rect 1854 10180 1860 10192
rect 1535 10152 1860 10180
rect 1535 10149 1547 10152
rect 1489 10143 1547 10149
rect 1854 10140 1860 10152
rect 1912 10180 1918 10192
rect 2866 10180 2872 10192
rect 1912 10152 2872 10180
rect 1912 10140 1918 10152
rect 2866 10140 2872 10152
rect 2924 10180 2930 10192
rect 5000 10180 5028 10220
rect 5074 10208 5080 10260
rect 5132 10248 5138 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 5132 10220 5457 10248
rect 5132 10208 5138 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 6270 10248 6276 10260
rect 5776 10220 6276 10248
rect 5776 10208 5782 10220
rect 6270 10208 6276 10220
rect 6328 10208 6334 10260
rect 6638 10248 6644 10260
rect 6599 10220 6644 10248
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 6733 10251 6791 10257
rect 6733 10217 6745 10251
rect 6779 10248 6791 10251
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 6779 10220 7481 10248
rect 6779 10217 6791 10220
rect 6733 10211 6791 10217
rect 5534 10180 5540 10192
rect 2924 10152 4936 10180
rect 5000 10152 5540 10180
rect 2924 10140 2930 10152
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 3694 10112 3700 10124
rect 2823 10084 3700 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3050 10044 3056 10056
rect 3011 10016 3056 10044
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 4338 9908 4344 9920
rect 3568 9880 4344 9908
rect 3568 9868 3574 9880
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 4614 9908 4620 9920
rect 4575 9880 4620 9908
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 4908 9908 4936 10152
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 5902 10140 5908 10192
rect 5960 10140 5966 10192
rect 4985 10115 5043 10121
rect 4985 10081 4997 10115
rect 5031 10112 5043 10115
rect 5626 10112 5632 10124
rect 5031 10084 5632 10112
rect 5031 10081 5043 10084
rect 4985 10075 5043 10081
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 5810 10112 5816 10124
rect 5771 10084 5816 10112
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 5920 10112 5948 10140
rect 6270 10112 6276 10124
rect 5920 10084 6276 10112
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6840 10112 6868 10220
rect 7469 10217 7481 10220
rect 7515 10248 7527 10251
rect 8294 10248 8300 10260
rect 7515 10220 8300 10248
rect 7515 10217 7527 10220
rect 7469 10211 7527 10217
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 10229 10251 10287 10257
rect 10229 10217 10241 10251
rect 10275 10248 10287 10251
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 10275 10220 10609 10248
rect 10275 10217 10287 10220
rect 10229 10211 10287 10217
rect 10597 10217 10609 10220
rect 10643 10217 10655 10251
rect 10597 10211 10655 10217
rect 10870 10208 10876 10260
rect 10928 10248 10934 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 10928 10220 11069 10248
rect 10928 10208 10934 10220
rect 11057 10217 11069 10220
rect 11103 10248 11115 10251
rect 11609 10251 11667 10257
rect 11609 10248 11621 10251
rect 11103 10220 11621 10248
rect 11103 10217 11115 10220
rect 11057 10211 11115 10217
rect 11609 10217 11621 10220
rect 11655 10217 11667 10251
rect 11609 10211 11667 10217
rect 11698 10208 11704 10260
rect 11756 10248 11762 10260
rect 11793 10251 11851 10257
rect 11793 10248 11805 10251
rect 11756 10220 11805 10248
rect 11756 10208 11762 10220
rect 11793 10217 11805 10220
rect 11839 10217 11851 10251
rect 11793 10211 11851 10217
rect 11977 10251 12035 10257
rect 11977 10217 11989 10251
rect 12023 10248 12035 10251
rect 12158 10248 12164 10260
rect 12023 10220 12164 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 12158 10208 12164 10220
rect 12216 10248 12222 10260
rect 14918 10248 14924 10260
rect 12216 10220 14924 10248
rect 12216 10208 12222 10220
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 15010 10208 15016 10260
rect 15068 10248 15074 10260
rect 15105 10251 15163 10257
rect 15105 10248 15117 10251
rect 15068 10220 15117 10248
rect 15068 10208 15074 10220
rect 15105 10217 15117 10220
rect 15151 10217 15163 10251
rect 15105 10211 15163 10217
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 16632 10220 16681 10248
rect 16632 10208 16638 10220
rect 16669 10217 16681 10220
rect 16715 10217 16727 10251
rect 16942 10248 16948 10260
rect 16903 10220 16948 10248
rect 16669 10211 16727 10217
rect 16942 10208 16948 10220
rect 17000 10208 17006 10260
rect 17402 10248 17408 10260
rect 17363 10220 17408 10248
rect 17402 10208 17408 10220
rect 17460 10208 17466 10260
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 17552 10220 18153 10248
rect 17552 10208 17558 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 18141 10211 18199 10217
rect 10137 10183 10195 10189
rect 10137 10149 10149 10183
rect 10183 10180 10195 10183
rect 10502 10180 10508 10192
rect 10183 10152 10508 10180
rect 10183 10149 10195 10152
rect 10137 10143 10195 10149
rect 10502 10140 10508 10152
rect 10560 10140 10566 10192
rect 10778 10140 10784 10192
rect 10836 10180 10842 10192
rect 10965 10183 11023 10189
rect 10965 10180 10977 10183
rect 10836 10152 10977 10180
rect 10836 10140 10842 10152
rect 10965 10149 10977 10152
rect 11011 10180 11023 10183
rect 13992 10183 14050 10189
rect 11011 10152 13952 10180
rect 11011 10149 11023 10152
rect 10965 10143 11023 10149
rect 7282 10112 7288 10124
rect 6512 10084 6868 10112
rect 6932 10084 7288 10112
rect 6512 10072 6518 10084
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5258 10044 5264 10056
rect 5219 10016 5264 10044
rect 5077 10007 5135 10013
rect 5092 9976 5120 10007
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5902 10044 5908 10056
rect 5863 10016 5908 10044
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10044 6147 10047
rect 6178 10044 6184 10056
rect 6135 10016 6184 10044
rect 6135 10013 6147 10016
rect 6089 10007 6147 10013
rect 6178 10004 6184 10016
rect 6236 10044 6242 10056
rect 6932 10053 6960 10084
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7374 10072 7380 10124
rect 7432 10112 7438 10124
rect 7834 10121 7840 10124
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 7432 10084 7573 10112
rect 7432 10072 7438 10084
rect 7561 10081 7573 10084
rect 7607 10081 7619 10115
rect 7828 10112 7840 10121
rect 7795 10084 7840 10112
rect 7561 10075 7619 10081
rect 7828 10075 7840 10084
rect 7892 10112 7898 10124
rect 8754 10112 8760 10124
rect 7892 10084 8760 10112
rect 7834 10072 7840 10075
rect 7892 10072 7898 10084
rect 8754 10072 8760 10084
rect 8812 10072 8818 10124
rect 11882 10112 11888 10124
rect 11072 10084 11888 10112
rect 6917 10047 6975 10053
rect 6917 10044 6929 10047
rect 6236 10016 6929 10044
rect 6236 10004 6242 10016
rect 6917 10013 6929 10016
rect 6963 10013 6975 10047
rect 7098 10044 7104 10056
rect 7059 10016 7104 10044
rect 6917 10007 6975 10013
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10044 10471 10047
rect 11072 10044 11100 10084
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 12529 10115 12587 10121
rect 12529 10081 12541 10115
rect 12575 10112 12587 10115
rect 13262 10112 13268 10124
rect 12575 10084 13268 10112
rect 12575 10081 12587 10084
rect 12529 10075 12587 10081
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 13814 10112 13820 10124
rect 13771 10084 13820 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 13924 10112 13952 10152
rect 13992 10149 14004 10183
rect 14038 10180 14050 10183
rect 16206 10180 16212 10192
rect 14038 10152 16212 10180
rect 14038 10149 14050 10152
rect 13992 10143 14050 10149
rect 16206 10140 16212 10152
rect 16264 10140 16270 10192
rect 17770 10140 17776 10192
rect 17828 10180 17834 10192
rect 18233 10183 18291 10189
rect 18233 10180 18245 10183
rect 17828 10152 18245 10180
rect 17828 10140 17834 10152
rect 18233 10149 18245 10152
rect 18279 10149 18291 10183
rect 18233 10143 18291 10149
rect 15556 10115 15614 10121
rect 13924 10084 14872 10112
rect 10459 10016 11100 10044
rect 11241 10047 11299 10053
rect 10459 10013 10471 10016
rect 10413 10007 10471 10013
rect 11241 10013 11253 10047
rect 11287 10044 11299 10047
rect 11330 10044 11336 10056
rect 11287 10016 11336 10044
rect 11287 10013 11299 10016
rect 11241 10007 11299 10013
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 12618 10044 12624 10056
rect 12579 10016 12624 10044
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10044 12863 10047
rect 13630 10044 13636 10056
rect 12851 10016 13636 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 6273 9979 6331 9985
rect 6273 9976 6285 9979
rect 5092 9948 6285 9976
rect 6273 9945 6285 9948
rect 6319 9945 6331 9979
rect 14844 9976 14872 10084
rect 15556 10081 15568 10115
rect 15602 10112 15614 10115
rect 16574 10112 16580 10124
rect 15602 10084 16580 10112
rect 15602 10081 15614 10084
rect 15556 10075 15614 10081
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 16850 10112 16856 10124
rect 16811 10084 16856 10112
rect 16850 10072 16856 10084
rect 16908 10112 16914 10124
rect 17313 10115 17371 10121
rect 17313 10112 17325 10115
rect 16908 10084 17325 10112
rect 16908 10072 16914 10084
rect 17313 10081 17325 10084
rect 17359 10112 17371 10115
rect 17954 10112 17960 10124
rect 17359 10084 17960 10112
rect 17359 10081 17371 10084
rect 17313 10075 17371 10081
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 14918 10004 14924 10056
rect 14976 10044 14982 10056
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 14976 10016 15301 10044
rect 14976 10004 14982 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 16592 10044 16620 10072
rect 17497 10047 17555 10053
rect 17497 10044 17509 10047
rect 16592 10016 17509 10044
rect 15289 10007 15347 10013
rect 17497 10013 17509 10016
rect 17543 10044 17555 10047
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 17543 10016 18337 10044
rect 17543 10013 17555 10016
rect 17497 10007 17555 10013
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 6273 9939 6331 9945
rect 7300 9948 7604 9976
rect 7300 9908 7328 9948
rect 4908 9880 7328 9908
rect 7576 9908 7604 9948
rect 8496 9948 9904 9976
rect 14844 9948 15332 9976
rect 8496 9908 8524 9948
rect 7576 9880 8524 9908
rect 8941 9911 8999 9917
rect 8941 9877 8953 9911
rect 8987 9908 8999 9911
rect 9398 9908 9404 9920
rect 8987 9880 9404 9908
rect 8987 9877 8999 9880
rect 8941 9871 8999 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 9766 9908 9772 9920
rect 9727 9880 9772 9908
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 9876 9908 9904 9948
rect 11425 9911 11483 9917
rect 11425 9908 11437 9911
rect 9876 9880 11437 9908
rect 11425 9877 11437 9880
rect 11471 9908 11483 9911
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11471 9880 11989 9908
rect 11471 9877 11483 9880
rect 11425 9871 11483 9877
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 12158 9908 12164 9920
rect 12119 9880 12164 9908
rect 11977 9871 12035 9877
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 13449 9911 13507 9917
rect 13449 9877 13461 9911
rect 13495 9908 13507 9911
rect 13538 9908 13544 9920
rect 13495 9880 13544 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 15304 9908 15332 9948
rect 16666 9936 16672 9988
rect 16724 9976 16730 9988
rect 17773 9979 17831 9985
rect 17773 9976 17785 9979
rect 16724 9948 17785 9976
rect 16724 9936 16730 9948
rect 17773 9945 17785 9948
rect 17819 9945 17831 9979
rect 17773 9939 17831 9945
rect 16850 9908 16856 9920
rect 15304 9880 16856 9908
rect 16850 9868 16856 9880
rect 16908 9868 16914 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 2866 9704 2872 9716
rect 2827 9676 2872 9704
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 3694 9704 3700 9716
rect 3655 9676 3700 9704
rect 3694 9664 3700 9676
rect 3752 9664 3758 9716
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 12434 9704 12440 9716
rect 3844 9676 12440 9704
rect 3844 9664 3850 9676
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 12713 9707 12771 9713
rect 12713 9704 12725 9707
rect 12676 9676 12725 9704
rect 12676 9664 12682 9676
rect 12713 9673 12725 9676
rect 12759 9673 12771 9707
rect 12713 9667 12771 9673
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 13541 9707 13599 9713
rect 13541 9704 13553 9707
rect 13320 9676 13553 9704
rect 13320 9664 13326 9676
rect 13541 9673 13553 9676
rect 13587 9673 13599 9707
rect 13541 9667 13599 9673
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 15194 9704 15200 9716
rect 13872 9676 15200 9704
rect 13872 9664 13878 9676
rect 15194 9664 15200 9676
rect 15252 9664 15258 9716
rect 16040 9676 16712 9704
rect 2501 9639 2559 9645
rect 2501 9605 2513 9639
rect 2547 9636 2559 9639
rect 2590 9636 2596 9648
rect 2547 9608 2596 9636
rect 2547 9605 2559 9608
rect 2501 9599 2559 9605
rect 2516 9568 2544 9599
rect 2590 9596 2596 9608
rect 2648 9596 2654 9648
rect 3510 9596 3516 9648
rect 3568 9636 3574 9648
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 3568 9608 4537 9636
rect 3568 9596 3574 9608
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 5442 9636 5448 9648
rect 4525 9599 4583 9605
rect 4724 9608 5448 9636
rect 4724 9580 4752 9608
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 5684 9608 5764 9636
rect 5684 9596 5690 9608
rect 1688 9540 2544 9568
rect 1688 9509 1716 9540
rect 3234 9528 3240 9580
rect 3292 9568 3298 9580
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 3292 9540 3433 9568
rect 3292 9528 3298 9540
rect 3421 9537 3433 9540
rect 3467 9568 3479 9571
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 3467 9540 4261 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4706 9568 4712 9580
rect 4249 9531 4307 9537
rect 4540 9540 4712 9568
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9469 1731 9503
rect 1673 9463 1731 9469
rect 2041 9503 2099 9509
rect 2041 9469 2053 9503
rect 2087 9469 2099 9503
rect 2041 9463 2099 9469
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 2056 9432 2084 9463
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 2832 9472 3341 9500
rect 2832 9460 2838 9472
rect 3329 9469 3341 9472
rect 3375 9500 3387 9503
rect 4540 9500 4568 9540
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4856 9540 4997 9568
rect 4856 9528 4862 9540
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5350 9568 5356 9580
rect 5215 9540 5356 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 5736 9568 5764 9608
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 5868 9608 5913 9636
rect 6012 9608 6837 9636
rect 5868 9596 5874 9608
rect 6012 9568 6040 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 6825 9599 6883 9605
rect 7024 9608 13216 9636
rect 5736 9540 6040 9568
rect 6362 9528 6368 9580
rect 6420 9568 6426 9580
rect 6420 9540 6465 9568
rect 6420 9528 6426 9540
rect 6638 9528 6644 9580
rect 6696 9568 6702 9580
rect 7024 9568 7052 9608
rect 6696 9540 7052 9568
rect 6696 9528 6702 9540
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7340 9540 7389 9568
rect 7340 9528 7346 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8573 9571 8631 9577
rect 8573 9568 8585 9571
rect 7892 9540 8585 9568
rect 7892 9528 7898 9540
rect 8573 9537 8585 9540
rect 8619 9568 8631 9571
rect 9214 9568 9220 9580
rect 8619 9540 9220 9568
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 9214 9528 9220 9540
rect 9272 9568 9278 9580
rect 10318 9568 10324 9580
rect 9272 9540 10180 9568
rect 10279 9540 10324 9568
rect 9272 9528 9278 9540
rect 3375 9472 4568 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 4672 9472 4905 9500
rect 4672 9460 4678 9472
rect 4893 9469 4905 9472
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 5132 9472 5549 9500
rect 5132 9460 5138 9472
rect 5537 9469 5549 9472
rect 5583 9469 5595 9503
rect 5537 9463 5595 9469
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 6656 9500 6684 9528
rect 6227 9472 6684 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 7098 9460 7104 9512
rect 7156 9500 7162 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 7156 9472 7205 9500
rect 7156 9460 7162 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7193 9463 7251 9469
rect 7300 9472 7757 9500
rect 7300 9441 7328 9472
rect 7745 9469 7757 9472
rect 7791 9500 7803 9503
rect 8018 9500 8024 9512
rect 7791 9472 8024 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 9858 9460 9864 9512
rect 9916 9500 9922 9512
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9916 9472 10057 9500
rect 9916 9460 9922 9472
rect 10045 9469 10057 9472
rect 10091 9469 10103 9503
rect 10152 9500 10180 9540
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10962 9568 10968 9580
rect 10923 9540 10968 9568
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11606 9568 11612 9580
rect 11072 9540 11612 9568
rect 11072 9500 11100 9540
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 11882 9568 11888 9580
rect 11843 9540 11888 9568
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 13188 9568 13216 9608
rect 13630 9596 13636 9648
rect 13688 9636 13694 9648
rect 13688 9608 14412 9636
rect 13688 9596 13694 9608
rect 13262 9568 13268 9580
rect 13188 9540 13268 9568
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 13357 9571 13415 9577
rect 13357 9537 13369 9571
rect 13403 9568 13415 9571
rect 13722 9568 13728 9580
rect 13403 9540 13728 9568
rect 13403 9537 13415 9540
rect 13357 9531 13415 9537
rect 13722 9528 13728 9540
rect 13780 9568 13786 9580
rect 14093 9571 14151 9577
rect 14093 9568 14105 9571
rect 13780 9540 14105 9568
rect 13780 9528 13786 9540
rect 14093 9537 14105 9540
rect 14139 9537 14151 9571
rect 14384 9568 14412 9608
rect 14458 9596 14464 9648
rect 14516 9636 14522 9648
rect 14829 9639 14887 9645
rect 14829 9636 14841 9639
rect 14516 9608 14841 9636
rect 14516 9596 14522 9608
rect 14829 9605 14841 9608
rect 14875 9605 14887 9639
rect 16040 9636 16068 9676
rect 14829 9599 14887 9605
rect 14936 9608 16068 9636
rect 14936 9568 14964 9608
rect 16206 9596 16212 9648
rect 16264 9596 16270 9648
rect 16485 9639 16543 9645
rect 16485 9636 16497 9639
rect 16408 9608 16497 9636
rect 14384 9540 14964 9568
rect 14093 9531 14151 9537
rect 15010 9528 15016 9580
rect 15068 9568 15074 9580
rect 15381 9571 15439 9577
rect 15381 9568 15393 9571
rect 15068 9540 15393 9568
rect 15068 9528 15074 9540
rect 15381 9537 15393 9540
rect 15427 9537 15439 9571
rect 16224 9568 16252 9596
rect 16301 9571 16359 9577
rect 16301 9568 16313 9571
rect 16224 9540 16313 9568
rect 15381 9531 15439 9537
rect 16301 9537 16313 9540
rect 16347 9537 16359 9571
rect 16301 9531 16359 9537
rect 10152 9472 11100 9500
rect 10045 9463 10103 9469
rect 11514 9460 11520 9512
rect 11572 9500 11578 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11572 9472 11713 9500
rect 11572 9460 11578 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 11793 9503 11851 9509
rect 11793 9469 11805 9503
rect 11839 9500 11851 9503
rect 12158 9500 12164 9512
rect 11839 9472 12164 9500
rect 11839 9469 11851 9472
rect 11793 9463 11851 9469
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 13998 9500 14004 9512
rect 13596 9472 14004 9500
rect 13596 9460 13602 9472
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 16206 9500 16212 9512
rect 15243 9472 16212 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 7285 9435 7343 9441
rect 7285 9432 7297 9435
rect 1627 9404 7297 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 7285 9401 7297 9404
rect 7331 9401 7343 9435
rect 9585 9435 9643 9441
rect 9585 9432 9597 9435
rect 7285 9395 7343 9401
rect 7852 9404 9597 9432
rect 1854 9364 1860 9376
rect 1815 9336 1860 9364
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 2222 9364 2228 9376
rect 2183 9336 2228 9364
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 3237 9367 3295 9373
rect 3237 9333 3249 9367
rect 3283 9364 3295 9367
rect 3418 9364 3424 9376
rect 3283 9336 3424 9364
rect 3283 9333 3295 9336
rect 3237 9327 3295 9333
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 4065 9367 4123 9373
rect 4065 9364 4077 9367
rect 4028 9336 4077 9364
rect 4028 9324 4034 9336
rect 4065 9333 4077 9336
rect 4111 9333 4123 9367
rect 4065 9327 4123 9333
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 5258 9364 5264 9376
rect 4212 9336 5264 9364
rect 4212 9324 4218 9336
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5353 9367 5411 9373
rect 5353 9333 5365 9367
rect 5399 9364 5411 9367
rect 5534 9364 5540 9376
rect 5399 9336 5540 9364
rect 5399 9333 5411 9336
rect 5353 9327 5411 9333
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 5721 9367 5779 9373
rect 5721 9364 5733 9367
rect 5684 9336 5733 9364
rect 5684 9324 5690 9336
rect 5721 9333 5733 9336
rect 5767 9364 5779 9367
rect 6273 9367 6331 9373
rect 6273 9364 6285 9367
rect 5767 9336 6285 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 6273 9333 6285 9336
rect 6319 9364 6331 9367
rect 6454 9364 6460 9376
rect 6319 9336 6460 9364
rect 6319 9333 6331 9336
rect 6273 9327 6331 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 7852 9364 7880 9404
rect 9585 9401 9597 9404
rect 9631 9432 9643 9435
rect 10226 9432 10232 9444
rect 9631 9404 10232 9432
rect 9631 9401 9643 9404
rect 9585 9395 9643 9401
rect 10226 9392 10232 9404
rect 10284 9432 10290 9444
rect 13078 9432 13084 9444
rect 10284 9404 11468 9432
rect 13039 9404 13084 9432
rect 10284 9392 10290 9404
rect 9674 9364 9680 9376
rect 6788 9336 7880 9364
rect 9635 9336 9680 9364
rect 6788 9324 6794 9336
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10137 9367 10195 9373
rect 10137 9333 10149 9367
rect 10183 9364 10195 9367
rect 11333 9367 11391 9373
rect 11333 9364 11345 9367
rect 10183 9336 11345 9364
rect 10183 9333 10195 9336
rect 10137 9327 10195 9333
rect 11333 9333 11345 9336
rect 11379 9333 11391 9367
rect 11440 9364 11468 9404
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 14461 9435 14519 9441
rect 14461 9401 14473 9435
rect 14507 9432 14519 9435
rect 15010 9432 15016 9444
rect 14507 9404 15016 9432
rect 14507 9401 14519 9404
rect 14461 9395 14519 9401
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 16025 9435 16083 9441
rect 16025 9401 16037 9435
rect 16071 9432 16083 9435
rect 16408 9432 16436 9608
rect 16485 9605 16497 9608
rect 16531 9605 16543 9639
rect 16684 9636 16712 9676
rect 17402 9664 17408 9716
rect 17460 9704 17466 9716
rect 17773 9707 17831 9713
rect 17773 9704 17785 9707
rect 17460 9676 17785 9704
rect 17460 9664 17466 9676
rect 17773 9673 17785 9676
rect 17819 9673 17831 9707
rect 17773 9667 17831 9673
rect 16942 9636 16948 9648
rect 16684 9608 16948 9636
rect 16485 9599 16543 9605
rect 16942 9596 16948 9608
rect 17000 9596 17006 9648
rect 17678 9596 17684 9648
rect 17736 9636 17742 9648
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 17736 9608 18245 9636
rect 17736 9596 17742 9608
rect 18233 9605 18245 9608
rect 18279 9605 18291 9639
rect 18233 9599 18291 9605
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16632 9540 17049 9568
rect 16632 9528 16638 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 16945 9503 17003 9509
rect 16945 9469 16957 9503
rect 16991 9500 17003 9503
rect 17586 9500 17592 9512
rect 16991 9472 17592 9500
rect 16991 9469 17003 9472
rect 16945 9463 17003 9469
rect 17586 9460 17592 9472
rect 17644 9460 17650 9512
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 18046 9460 18052 9472
rect 18104 9500 18110 9512
rect 18417 9503 18475 9509
rect 18417 9500 18429 9503
rect 18104 9472 18429 9500
rect 18104 9460 18110 9472
rect 18417 9469 18429 9472
rect 18463 9469 18475 9503
rect 18417 9463 18475 9469
rect 16071 9404 16436 9432
rect 16071 9401 16083 9404
rect 16025 9395 16083 9401
rect 16482 9392 16488 9444
rect 16540 9432 16546 9444
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 16540 9404 16865 9432
rect 16540 9392 16546 9404
rect 16853 9401 16865 9404
rect 16899 9432 16911 9435
rect 17402 9432 17408 9444
rect 16899 9404 17408 9432
rect 16899 9401 16911 9404
rect 16853 9395 16911 9401
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 17494 9392 17500 9444
rect 17552 9432 17558 9444
rect 17862 9432 17868 9444
rect 17552 9404 17868 9432
rect 17552 9392 17558 9404
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 12529 9367 12587 9373
rect 12529 9364 12541 9367
rect 11440 9336 12541 9364
rect 11333 9327 11391 9333
rect 12529 9333 12541 9336
rect 12575 9364 12587 9367
rect 13173 9367 13231 9373
rect 13173 9364 13185 9367
rect 12575 9336 13185 9364
rect 12575 9333 12587 9336
rect 12529 9327 12587 9333
rect 13173 9333 13185 9336
rect 13219 9364 13231 9367
rect 13630 9364 13636 9376
rect 13219 9336 13636 9364
rect 13219 9333 13231 9336
rect 13173 9327 13231 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 13909 9367 13967 9373
rect 13909 9364 13921 9367
rect 13780 9336 13921 9364
rect 13780 9324 13786 9336
rect 13909 9333 13921 9336
rect 13955 9364 13967 9367
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 13955 9336 14657 9364
rect 13955 9333 13967 9336
rect 13909 9327 13967 9333
rect 14645 9333 14657 9336
rect 14691 9364 14703 9367
rect 15194 9364 15200 9376
rect 14691 9336 15200 9364
rect 14691 9333 14703 9336
rect 14645 9327 14703 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 15289 9367 15347 9373
rect 15289 9333 15301 9367
rect 15335 9364 15347 9367
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 15335 9336 15669 9364
rect 15335 9333 15347 9336
rect 15289 9327 15347 9333
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 15657 9327 15715 9333
rect 16117 9367 16175 9373
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 16574 9364 16580 9376
rect 16163 9336 16580 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 17681 9367 17739 9373
rect 17681 9364 17693 9367
rect 17276 9336 17693 9364
rect 17276 9324 17282 9336
rect 17681 9333 17693 9336
rect 17727 9364 17739 9367
rect 17770 9364 17776 9376
rect 17727 9336 17776 9364
rect 17727 9333 17739 9336
rect 17681 9327 17739 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 3234 9160 3240 9172
rect 3195 9132 3240 9160
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3602 9160 3608 9172
rect 3515 9132 3608 9160
rect 3602 9120 3608 9132
rect 3660 9160 3666 9172
rect 4154 9160 4160 9172
rect 3660 9132 4160 9160
rect 3660 9120 3666 9132
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 5166 9160 5172 9172
rect 4264 9132 5172 9160
rect 3418 9052 3424 9104
rect 3476 9092 3482 9104
rect 3789 9095 3847 9101
rect 3789 9092 3801 9095
rect 3476 9064 3801 9092
rect 3476 9052 3482 9064
rect 3789 9061 3801 9064
rect 3835 9092 3847 9095
rect 4264 9092 4292 9132
rect 5166 9120 5172 9132
rect 5224 9160 5230 9172
rect 5442 9160 5448 9172
rect 5224 9132 5448 9160
rect 5224 9120 5230 9132
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 5813 9163 5871 9169
rect 5813 9129 5825 9163
rect 5859 9160 5871 9163
rect 5902 9160 5908 9172
rect 5859 9132 5908 9160
rect 5859 9129 5871 9132
rect 5813 9123 5871 9129
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 6181 9163 6239 9169
rect 6181 9129 6193 9163
rect 6227 9160 6239 9163
rect 6227 9132 6592 9160
rect 6227 9129 6239 9132
rect 6181 9123 6239 9129
rect 3835 9064 4292 9092
rect 3835 9061 3847 9064
rect 3789 9055 3847 9061
rect 5350 9052 5356 9104
rect 5408 9092 5414 9104
rect 5629 9095 5687 9101
rect 5629 9092 5641 9095
rect 5408 9064 5641 9092
rect 5408 9052 5414 9064
rect 5629 9061 5641 9064
rect 5675 9092 5687 9095
rect 6273 9095 6331 9101
rect 6273 9092 6285 9095
rect 5675 9064 6285 9092
rect 5675 9061 5687 9064
rect 5629 9055 5687 9061
rect 6273 9061 6285 9064
rect 6319 9061 6331 9095
rect 6273 9055 6331 9061
rect 6362 9052 6368 9104
rect 6420 9052 6426 9104
rect 6564 9092 6592 9132
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 12805 9163 12863 9169
rect 12805 9160 12817 9163
rect 6788 9132 12817 9160
rect 6788 9120 6794 9132
rect 12805 9129 12817 9132
rect 12851 9160 12863 9163
rect 13449 9163 13507 9169
rect 13449 9160 13461 9163
rect 12851 9132 13461 9160
rect 12851 9129 12863 9132
rect 12805 9123 12863 9129
rect 13449 9129 13461 9132
rect 13495 9160 13507 9163
rect 16577 9163 16635 9169
rect 16577 9160 16589 9163
rect 13495 9132 16589 9160
rect 13495 9129 13507 9132
rect 13449 9123 13507 9129
rect 16577 9129 16589 9132
rect 16623 9129 16635 9163
rect 17586 9160 17592 9172
rect 17547 9132 17592 9160
rect 16577 9123 16635 9129
rect 6564 9064 6776 9092
rect 2124 9027 2182 9033
rect 2124 8993 2136 9027
rect 2170 9024 2182 9027
rect 2682 9024 2688 9036
rect 2170 8996 2688 9024
rect 2170 8993 2182 8996
rect 2124 8987 2182 8993
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 9024 4399 9027
rect 5810 9024 5816 9036
rect 4387 8996 5816 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1762 8956 1768 8968
rect 1544 8928 1768 8956
rect 1544 8916 1550 8928
rect 1762 8916 1768 8928
rect 1820 8956 1826 8968
rect 1857 8959 1915 8965
rect 1857 8956 1869 8959
rect 1820 8928 1869 8956
rect 1820 8916 1826 8928
rect 1857 8925 1869 8928
rect 1903 8925 1915 8959
rect 1857 8919 1915 8925
rect 4246 8916 4252 8968
rect 4304 8956 4310 8968
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 4304 8928 4537 8956
rect 4304 8916 4310 8928
rect 4525 8925 4537 8928
rect 4571 8925 4583 8959
rect 4982 8956 4988 8968
rect 4943 8928 4988 8956
rect 4525 8919 4583 8925
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 5074 8916 5080 8968
rect 5132 8956 5138 8968
rect 6270 8956 6276 8968
rect 5132 8928 6276 8956
rect 5132 8916 5138 8928
rect 6270 8916 6276 8928
rect 6328 8916 6334 8968
rect 6380 8965 6408 9052
rect 6748 9036 6776 9064
rect 7006 9052 7012 9104
rect 7064 9092 7070 9104
rect 9674 9092 9680 9104
rect 7064 9064 9680 9092
rect 7064 9052 7070 9064
rect 9674 9052 9680 9064
rect 9732 9052 9738 9104
rect 10134 9092 10140 9104
rect 10095 9064 10140 9092
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 16301 9095 16359 9101
rect 16301 9092 16313 9095
rect 10284 9064 16313 9092
rect 10284 9052 10290 9064
rect 16301 9061 16313 9064
rect 16347 9092 16359 9095
rect 16482 9092 16488 9104
rect 16347 9064 16488 9092
rect 16347 9061 16359 9064
rect 16301 9055 16359 9061
rect 16482 9052 16488 9064
rect 16540 9052 16546 9104
rect 16592 9092 16620 9123
rect 17586 9120 17592 9132
rect 17644 9120 17650 9172
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 17920 9132 18061 9160
rect 17920 9120 17926 9132
rect 18049 9129 18061 9132
rect 18095 9160 18107 9163
rect 18690 9160 18696 9172
rect 18095 9132 18696 9160
rect 18095 9129 18107 9132
rect 18049 9123 18107 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 17221 9095 17279 9101
rect 17221 9092 17233 9095
rect 16592 9064 17233 9092
rect 17221 9061 17233 9064
rect 17267 9092 17279 9095
rect 17494 9092 17500 9104
rect 17267 9064 17500 9092
rect 17267 9061 17279 9064
rect 17221 9055 17279 9061
rect 17494 9052 17500 9064
rect 17552 9052 17558 9104
rect 17957 9095 18015 9101
rect 17957 9092 17969 9095
rect 17604 9064 17969 9092
rect 6730 9024 6736 9036
rect 6691 8996 6736 9024
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 7460 9027 7518 9033
rect 7460 8993 7472 9027
rect 7506 9024 7518 9027
rect 8938 9024 8944 9036
rect 7506 8996 8944 9024
rect 7506 8993 7518 8996
rect 7460 8987 7518 8993
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 9122 9024 9128 9036
rect 9035 8996 9128 9024
rect 9122 8984 9128 8996
rect 9180 9024 9186 9036
rect 9950 9024 9956 9036
rect 9180 8996 9956 9024
rect 9180 8984 9186 8996
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10594 9024 10600 9036
rect 10091 8996 10600 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6696 8928 6837 8956
rect 6696 8916 6702 8928
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8925 7251 8959
rect 9214 8956 9220 8968
rect 9175 8928 9220 8956
rect 7193 8919 7251 8925
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 7208 8888 7236 8919
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9398 8956 9404 8968
rect 9359 8928 9404 8956
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 10060 8956 10088 8987
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 10778 9024 10784 9036
rect 10739 8996 10784 9024
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 11232 9027 11290 9033
rect 11232 8993 11244 9027
rect 11278 9024 11290 9027
rect 11606 9024 11612 9036
rect 11278 8996 11612 9024
rect 11278 8993 11290 8996
rect 11232 8987 11290 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 12713 9027 12771 9033
rect 12713 9024 12725 9027
rect 11756 8996 12725 9024
rect 11756 8984 11762 8996
rect 12713 8993 12725 8996
rect 12759 8993 12771 9027
rect 12713 8987 12771 8993
rect 13262 8984 13268 9036
rect 13320 9024 13326 9036
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 13320 8996 13369 9024
rect 13320 8984 13326 8996
rect 13357 8993 13369 8996
rect 13403 9024 13415 9027
rect 13817 9027 13875 9033
rect 13817 9024 13829 9027
rect 13403 8996 13829 9024
rect 13403 8993 13415 8996
rect 13357 8987 13415 8993
rect 13817 8993 13829 8996
rect 13863 9024 13875 9027
rect 16117 9027 16175 9033
rect 16117 9024 16129 9027
rect 13863 8996 16129 9024
rect 13863 8993 13875 8996
rect 13817 8987 13875 8993
rect 16117 8993 16129 8996
rect 16163 9024 16175 9027
rect 17126 9024 17132 9036
rect 16163 8996 17132 9024
rect 16163 8993 16175 8996
rect 16117 8987 16175 8993
rect 17126 8984 17132 8996
rect 17184 8984 17190 9036
rect 17604 9024 17632 9064
rect 17957 9061 17969 9064
rect 18003 9092 18015 9095
rect 18138 9092 18144 9104
rect 18003 9064 18144 9092
rect 18003 9061 18015 9064
rect 17957 9055 18015 9061
rect 18138 9052 18144 9064
rect 18196 9052 18202 9104
rect 18417 9027 18475 9033
rect 18417 9024 18429 9027
rect 17236 8996 17632 9024
rect 17788 8996 18429 9024
rect 9548 8928 10088 8956
rect 10321 8959 10379 8965
rect 9548 8916 9554 8928
rect 10321 8925 10333 8959
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 5592 8860 7236 8888
rect 8128 8860 8892 8888
rect 5592 8848 5598 8860
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 8128 8820 8156 8860
rect 8570 8820 8576 8832
rect 5960 8792 8156 8820
rect 8531 8792 8576 8820
rect 5960 8780 5966 8792
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 8754 8820 8760 8832
rect 8715 8792 8760 8820
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 8864 8820 8892 8860
rect 8938 8848 8944 8900
rect 8996 8888 9002 8900
rect 9416 8888 9444 8916
rect 10226 8888 10232 8900
rect 8996 8860 9444 8888
rect 9508 8860 10232 8888
rect 8996 8848 9002 8860
rect 9508 8820 9536 8860
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 9674 8820 9680 8832
rect 8864 8792 9536 8820
rect 9635 8792 9680 8820
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10336 8820 10364 8919
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 10980 8888 11008 8919
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 13596 8928 13641 8956
rect 13596 8916 13602 8928
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 15194 8956 15200 8968
rect 14056 8928 15200 8956
rect 14056 8916 14062 8928
rect 15194 8916 15200 8928
rect 15252 8916 15258 8968
rect 16025 8959 16083 8965
rect 16025 8925 16037 8959
rect 16071 8956 16083 8959
rect 17236 8956 17264 8996
rect 16071 8928 17264 8956
rect 16071 8925 16083 8928
rect 16025 8919 16083 8925
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17368 8928 17413 8956
rect 17368 8916 17374 8928
rect 17494 8916 17500 8968
rect 17552 8956 17558 8968
rect 17788 8956 17816 8996
rect 18417 8993 18429 8996
rect 18463 8993 18475 9027
rect 18417 8987 18475 8993
rect 17552 8928 17816 8956
rect 18141 8959 18199 8965
rect 17552 8916 17558 8928
rect 18141 8925 18153 8959
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 10468 8860 11008 8888
rect 10468 8848 10474 8860
rect 10778 8820 10784 8832
rect 9824 8792 10784 8820
rect 9824 8780 9830 8792
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 10980 8820 11008 8860
rect 11900 8860 12572 8888
rect 11900 8820 11928 8860
rect 10980 8792 11928 8820
rect 12345 8823 12403 8829
rect 12345 8789 12357 8823
rect 12391 8820 12403 8823
rect 12434 8820 12440 8832
rect 12391 8792 12440 8820
rect 12391 8789 12403 8792
rect 12345 8783 12403 8789
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 12544 8829 12572 8860
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 12989 8891 13047 8897
rect 12989 8888 13001 8891
rect 12768 8860 13001 8888
rect 12768 8848 12774 8860
rect 12989 8857 13001 8860
rect 13035 8857 13047 8891
rect 12989 8851 13047 8857
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 17328 8888 17356 8916
rect 18156 8888 18184 8919
rect 16540 8860 16896 8888
rect 17328 8860 18184 8888
rect 16540 8848 16546 8860
rect 12529 8823 12587 8829
rect 12529 8789 12541 8823
rect 12575 8820 12587 8823
rect 13906 8820 13912 8832
rect 12575 8792 13912 8820
rect 12575 8789 12587 8792
rect 12529 8783 12587 8789
rect 13906 8780 13912 8792
rect 13964 8820 13970 8832
rect 14918 8820 14924 8832
rect 13964 8792 14924 8820
rect 13964 8780 13970 8792
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 16298 8780 16304 8832
rect 16356 8820 16362 8832
rect 16761 8823 16819 8829
rect 16761 8820 16773 8823
rect 16356 8792 16773 8820
rect 16356 8780 16362 8792
rect 16761 8789 16773 8792
rect 16807 8789 16819 8823
rect 16868 8820 16896 8860
rect 17954 8820 17960 8832
rect 16868 8792 17960 8820
rect 16761 8783 16819 8789
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 2869 8619 2927 8625
rect 2869 8616 2881 8619
rect 2740 8588 2881 8616
rect 2740 8576 2746 8588
rect 2869 8585 2881 8588
rect 2915 8585 2927 8619
rect 2869 8579 2927 8585
rect 3053 8619 3111 8625
rect 3053 8585 3065 8619
rect 3099 8616 3111 8619
rect 3418 8616 3424 8628
rect 3099 8588 3424 8616
rect 3099 8585 3111 8588
rect 3053 8579 3111 8585
rect 3418 8576 3424 8588
rect 3476 8616 3482 8628
rect 3786 8616 3792 8628
rect 3476 8588 3792 8616
rect 3476 8576 3482 8588
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 5350 8616 5356 8628
rect 5311 8588 5356 8616
rect 5350 8576 5356 8588
rect 5408 8616 5414 8628
rect 11054 8616 11060 8628
rect 5408 8588 11060 8616
rect 5408 8576 5414 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 13354 8616 13360 8628
rect 11572 8588 13360 8616
rect 11572 8576 11578 8588
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 13909 8619 13967 8625
rect 13909 8585 13921 8619
rect 13955 8616 13967 8619
rect 15933 8619 15991 8625
rect 13955 8588 15516 8616
rect 13955 8585 13967 8588
rect 13909 8579 13967 8585
rect 3326 8548 3332 8560
rect 3287 8520 3332 8548
rect 3326 8508 3332 8520
rect 3384 8508 3390 8560
rect 4614 8508 4620 8560
rect 4672 8548 4678 8560
rect 5902 8548 5908 8560
rect 4672 8520 5908 8548
rect 4672 8508 4678 8520
rect 5902 8508 5908 8520
rect 5960 8508 5966 8560
rect 6362 8548 6368 8560
rect 6323 8520 6368 8548
rect 6362 8508 6368 8520
rect 6420 8508 6426 8560
rect 8754 8548 8760 8560
rect 7852 8520 8760 8548
rect 1486 8480 1492 8492
rect 1447 8452 1492 8480
rect 1486 8440 1492 8452
rect 1544 8440 1550 8492
rect 6086 8480 6092 8492
rect 6047 8452 6092 8480
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 7374 8440 7380 8492
rect 7432 8480 7438 8492
rect 7650 8480 7656 8492
rect 7432 8452 7656 8480
rect 7432 8440 7438 8452
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 1504 8412 1532 8440
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 1504 8384 3525 8412
rect 3513 8381 3525 8384
rect 3559 8412 3571 8415
rect 5626 8412 5632 8424
rect 3559 8384 5632 8412
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 6549 8415 6607 8421
rect 6549 8381 6561 8415
rect 6595 8412 6607 8415
rect 7742 8412 7748 8424
rect 6595 8384 7748 8412
rect 6595 8381 6607 8384
rect 6549 8375 6607 8381
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 7852 8412 7880 8520
rect 8754 8508 8760 8520
rect 8812 8508 8818 8560
rect 8846 8508 8852 8560
rect 8904 8548 8910 8560
rect 9674 8548 9680 8560
rect 8904 8520 9680 8548
rect 8904 8508 8910 8520
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 12618 8508 12624 8560
rect 12676 8548 12682 8560
rect 12989 8551 13047 8557
rect 12989 8548 13001 8551
rect 12676 8520 13001 8548
rect 12676 8508 12682 8520
rect 12989 8517 13001 8520
rect 13035 8517 13047 8551
rect 13814 8548 13820 8560
rect 12989 8511 13047 8517
rect 13407 8520 13820 8548
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8480 8263 8483
rect 8570 8480 8576 8492
rect 8251 8452 8576 8480
rect 8251 8449 8263 8452
rect 8205 8443 8263 8449
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 9766 8480 9772 8492
rect 9456 8452 9772 8480
rect 9456 8440 9462 8452
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10410 8480 10416 8492
rect 10100 8452 10416 8480
rect 10100 8440 10106 8452
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10778 8480 10784 8492
rect 10739 8452 10784 8480
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 13407 8480 13435 8520
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 13538 8480 13544 8492
rect 11164 8452 13435 8480
rect 13499 8452 13544 8480
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7852 8384 7941 8412
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 8386 8412 8392 8424
rect 8347 8384 8392 8412
rect 7929 8375 7987 8381
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 10226 8412 10232 8424
rect 8720 8384 10232 8412
rect 8720 8372 8726 8384
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8412 10655 8415
rect 10870 8412 10876 8424
rect 10643 8384 10876 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 10870 8372 10876 8384
rect 10928 8412 10934 8424
rect 11164 8421 11192 8452
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 11149 8415 11207 8421
rect 11149 8412 11161 8415
rect 10928 8384 11161 8412
rect 10928 8372 10934 8384
rect 11149 8381 11161 8384
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 11330 8372 11336 8424
rect 11388 8412 11394 8424
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 11388 8384 13369 8412
rect 11388 8372 11394 8384
rect 13357 8381 13369 8384
rect 13403 8412 13415 8415
rect 13924 8412 13952 8579
rect 15488 8548 15516 8588
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16666 8616 16672 8628
rect 15979 8588 16672 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16666 8576 16672 8588
rect 16724 8616 16730 8628
rect 17218 8616 17224 8628
rect 16724 8588 17224 8616
rect 16724 8576 16730 8588
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 17126 8548 17132 8560
rect 15488 8520 17132 8548
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 17773 8551 17831 8557
rect 17773 8517 17785 8551
rect 17819 8517 17831 8551
rect 17773 8511 17831 8517
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 14056 8452 14565 8480
rect 14056 8440 14062 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 16482 8480 16488 8492
rect 16443 8452 16488 8480
rect 14553 8443 14611 8449
rect 16482 8440 16488 8452
rect 16540 8440 16546 8492
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8480 16727 8483
rect 16758 8480 16764 8492
rect 16715 8452 16764 8480
rect 16715 8449 16727 8452
rect 16669 8443 16727 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 17310 8480 17316 8492
rect 16868 8452 17316 8480
rect 16500 8412 16528 8440
rect 13403 8384 13952 8412
rect 14752 8384 16528 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 1756 8347 1814 8353
rect 1756 8313 1768 8347
rect 1802 8344 1814 8347
rect 2498 8344 2504 8356
rect 1802 8316 2504 8344
rect 1802 8313 1814 8316
rect 1756 8307 1814 8313
rect 2498 8304 2504 8316
rect 2556 8304 2562 8356
rect 3786 8353 3792 8356
rect 3780 8344 3792 8353
rect 3747 8316 3792 8344
rect 3780 8307 3792 8316
rect 3786 8304 3792 8307
rect 3844 8304 3850 8356
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 5997 8347 6055 8353
rect 5997 8344 6009 8347
rect 5408 8316 6009 8344
rect 5408 8304 5414 8316
rect 5997 8313 6009 8316
rect 6043 8313 6055 8347
rect 5997 8307 6055 8313
rect 8021 8347 8079 8353
rect 8021 8313 8033 8347
rect 8067 8344 8079 8347
rect 8846 8344 8852 8356
rect 8067 8316 8852 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 8846 8304 8852 8316
rect 8904 8304 8910 8356
rect 8938 8304 8944 8356
rect 8996 8344 9002 8356
rect 10137 8347 10195 8353
rect 10137 8344 10149 8347
rect 8996 8316 10149 8344
rect 8996 8304 9002 8316
rect 10137 8313 10149 8316
rect 10183 8344 10195 8347
rect 10962 8344 10968 8356
rect 10183 8316 10968 8344
rect 10183 8313 10195 8316
rect 10137 8307 10195 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 11112 8316 12909 8344
rect 11112 8304 11118 8316
rect 12897 8313 12909 8316
rect 12943 8344 12955 8347
rect 13449 8347 13507 8353
rect 13449 8344 13461 8347
rect 12943 8316 13461 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 13449 8313 13461 8316
rect 13495 8344 13507 8347
rect 14752 8344 14780 8384
rect 13495 8316 14780 8344
rect 14820 8347 14878 8353
rect 13495 8313 13507 8316
rect 13449 8307 13507 8313
rect 14820 8313 14832 8347
rect 14866 8344 14878 8347
rect 16666 8344 16672 8356
rect 14866 8316 16672 8344
rect 14866 8313 14878 8316
rect 14820 8307 14878 8313
rect 16666 8304 16672 8316
rect 16724 8344 16730 8356
rect 16868 8344 16896 8452
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 17788 8480 17816 8511
rect 17862 8508 17868 8560
rect 17920 8548 17926 8560
rect 18233 8551 18291 8557
rect 18233 8548 18245 8551
rect 17920 8520 18245 8548
rect 17920 8508 17926 8520
rect 18233 8517 18245 8520
rect 18279 8517 18291 8551
rect 18233 8511 18291 8517
rect 18138 8480 18144 8492
rect 17788 8452 18144 8480
rect 18138 8440 18144 8452
rect 18196 8440 18202 8492
rect 17126 8412 17132 8424
rect 17087 8384 17132 8412
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17586 8412 17592 8424
rect 17547 8384 17592 8412
rect 17586 8372 17592 8384
rect 17644 8372 17650 8424
rect 18046 8412 18052 8424
rect 18007 8384 18052 8412
rect 18046 8372 18052 8384
rect 18104 8412 18110 8424
rect 18417 8415 18475 8421
rect 18417 8412 18429 8415
rect 18104 8384 18429 8412
rect 18104 8372 18110 8384
rect 18417 8381 18429 8384
rect 18463 8381 18475 8415
rect 18417 8375 18475 8381
rect 17954 8344 17960 8356
rect 16724 8316 16896 8344
rect 17696 8316 17960 8344
rect 16724 8304 16730 8316
rect 4890 8276 4896 8288
rect 4851 8248 4896 8276
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 5534 8276 5540 8288
rect 5495 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 5902 8276 5908 8288
rect 5863 8248 5908 8276
rect 5902 8236 5908 8248
rect 5960 8276 5966 8288
rect 6730 8276 6736 8288
rect 5960 8248 6736 8276
rect 5960 8236 5966 8248
rect 6730 8236 6736 8248
rect 6788 8276 6794 8288
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6788 8248 6837 8276
rect 6788 8236 6794 8248
rect 6825 8245 6837 8248
rect 6871 8245 6883 8279
rect 7558 8276 7564 8288
rect 7519 8248 7564 8276
rect 6825 8239 6883 8245
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 8662 8276 8668 8288
rect 7708 8248 8668 8276
rect 7708 8236 7714 8248
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 10226 8276 10232 8288
rect 10187 8248 10232 8276
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 10410 8236 10416 8288
rect 10468 8276 10474 8288
rect 10689 8279 10747 8285
rect 10689 8276 10701 8279
rect 10468 8248 10701 8276
rect 10468 8236 10474 8248
rect 10689 8245 10701 8248
rect 10735 8245 10747 8279
rect 10689 8239 10747 8245
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 15562 8276 15568 8288
rect 10836 8248 15568 8276
rect 10836 8236 10842 8248
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 16761 8279 16819 8285
rect 16761 8245 16773 8279
rect 16807 8276 16819 8279
rect 17034 8276 17040 8288
rect 16807 8248 17040 8276
rect 16807 8245 16819 8248
rect 16761 8239 16819 8245
rect 17034 8236 17040 8248
rect 17092 8236 17098 8288
rect 17221 8279 17279 8285
rect 17221 8245 17233 8279
rect 17267 8276 17279 8279
rect 17696 8276 17724 8316
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 17267 8248 17724 8276
rect 17267 8245 17279 8248
rect 17221 8239 17279 8245
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8072 2743 8075
rect 3053 8075 3111 8081
rect 3053 8072 3065 8075
rect 2731 8044 3065 8072
rect 2731 8041 2743 8044
rect 2685 8035 2743 8041
rect 3053 8041 3065 8044
rect 3099 8041 3111 8075
rect 3418 8072 3424 8084
rect 3379 8044 3424 8072
rect 3053 8035 3111 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4893 8075 4951 8081
rect 4893 8072 4905 8075
rect 4571 8044 4905 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 4893 8041 4905 8044
rect 4939 8041 4951 8075
rect 4893 8035 4951 8041
rect 5353 8075 5411 8081
rect 5353 8041 5365 8075
rect 5399 8072 5411 8075
rect 5534 8072 5540 8084
rect 5399 8044 5540 8072
rect 5399 8041 5411 8044
rect 5353 8035 5411 8041
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 6178 8032 6184 8084
rect 6236 8072 6242 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 6236 8044 7297 8072
rect 6236 8032 6242 8044
rect 7285 8041 7297 8044
rect 7331 8072 7343 8075
rect 7650 8072 7656 8084
rect 7331 8044 7656 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 7837 8075 7895 8081
rect 7837 8041 7849 8075
rect 7883 8072 7895 8075
rect 8297 8075 8355 8081
rect 8297 8072 8309 8075
rect 7883 8044 8309 8072
rect 7883 8041 7895 8044
rect 7837 8035 7895 8041
rect 8297 8041 8309 8044
rect 8343 8041 8355 8075
rect 8662 8072 8668 8084
rect 8623 8044 8668 8072
rect 8297 8035 8355 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 10226 8072 10232 8084
rect 8803 8044 10232 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 11606 8072 11612 8084
rect 11567 8044 11612 8072
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 12618 8072 12624 8084
rect 12579 8044 12624 8072
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 13817 8075 13875 8081
rect 13817 8072 13829 8075
rect 13372 8044 13829 8072
rect 5988 8007 6046 8013
rect 3344 7976 4752 8004
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 2593 7939 2651 7945
rect 1719 7908 2084 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 2056 7744 2084 7908
rect 2593 7905 2605 7939
rect 2639 7936 2651 7939
rect 2958 7936 2964 7948
rect 2639 7908 2964 7936
rect 2639 7905 2651 7908
rect 2593 7899 2651 7905
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2556 7840 2881 7868
rect 2556 7828 2562 7840
rect 2869 7837 2881 7840
rect 2915 7868 2927 7871
rect 3344 7868 3372 7976
rect 3418 7896 3424 7948
rect 3476 7936 3482 7948
rect 3513 7939 3571 7945
rect 3513 7936 3525 7939
rect 3476 7908 3525 7936
rect 3476 7896 3482 7908
rect 3513 7905 3525 7908
rect 3559 7905 3571 7939
rect 4430 7936 4436 7948
rect 4391 7908 4436 7936
rect 3513 7899 3571 7905
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 2915 7840 3372 7868
rect 3697 7871 3755 7877
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3697 7837 3709 7871
rect 3743 7868 3755 7871
rect 3786 7868 3792 7880
rect 3743 7840 3792 7868
rect 3743 7837 3755 7840
rect 3697 7831 3755 7837
rect 3786 7828 3792 7840
rect 3844 7868 3850 7880
rect 4724 7877 4752 7976
rect 5988 7973 6000 8007
rect 6034 8004 6046 8007
rect 6086 8004 6092 8016
rect 6034 7976 6092 8004
rect 6034 7973 6046 7976
rect 5988 7967 6046 7973
rect 6086 7964 6092 7976
rect 6144 7964 6150 8016
rect 7558 7964 7564 8016
rect 7616 8004 7622 8016
rect 7929 8007 7987 8013
rect 7929 8004 7941 8007
rect 7616 7976 7941 8004
rect 7616 7964 7622 7976
rect 7929 7973 7941 7976
rect 7975 7973 7987 8007
rect 7929 7967 7987 7973
rect 8018 7964 8024 8016
rect 8076 8004 8082 8016
rect 10410 8004 10416 8016
rect 8076 7976 10416 8004
rect 8076 7964 8082 7976
rect 10410 7964 10416 7976
rect 10468 8013 10474 8016
rect 10468 8007 10532 8013
rect 10468 7973 10486 8007
rect 10520 7973 10532 8007
rect 12342 8004 12348 8016
rect 10468 7967 10532 7973
rect 10888 7976 12348 8004
rect 10468 7964 10474 7967
rect 5261 7939 5319 7945
rect 5261 7905 5273 7939
rect 5307 7936 5319 7939
rect 5534 7936 5540 7948
rect 5307 7908 5540 7936
rect 5307 7905 5319 7908
rect 5261 7899 5319 7905
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 5684 7908 5733 7936
rect 5684 7896 5690 7908
rect 5721 7905 5733 7908
rect 5767 7905 5779 7939
rect 5721 7899 5779 7905
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 10888 7936 10916 7976
rect 12342 7964 12348 7976
rect 12400 7964 12406 8016
rect 12529 8007 12587 8013
rect 12529 7973 12541 8007
rect 12575 8004 12587 8007
rect 12710 8004 12716 8016
rect 12575 7976 12716 8004
rect 12575 7973 12587 7976
rect 12529 7967 12587 7973
rect 12710 7964 12716 7976
rect 12768 7964 12774 8016
rect 13170 7964 13176 8016
rect 13228 8004 13234 8016
rect 13372 8013 13400 8044
rect 13817 8041 13829 8044
rect 13863 8072 13875 8075
rect 15102 8072 15108 8084
rect 13863 8044 15108 8072
rect 13863 8041 13875 8044
rect 13817 8035 13875 8041
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15470 8032 15476 8084
rect 15528 8032 15534 8084
rect 16666 8072 16672 8084
rect 16627 8044 16672 8072
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 17586 8072 17592 8084
rect 16816 8044 17592 8072
rect 16816 8032 16822 8044
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 13357 8007 13415 8013
rect 13357 8004 13369 8007
rect 13228 7976 13369 8004
rect 13228 7964 13234 7976
rect 13357 7973 13369 7976
rect 13403 7973 13415 8007
rect 13357 7967 13415 7973
rect 13722 7964 13728 8016
rect 13780 8004 13786 8016
rect 15488 8004 15516 8032
rect 13780 7976 15516 8004
rect 13780 7964 13786 7976
rect 17034 7964 17040 8016
rect 17092 8004 17098 8016
rect 17221 8007 17279 8013
rect 17221 8004 17233 8007
rect 17092 7976 17233 8004
rect 17092 7964 17098 7976
rect 17221 7973 17233 7976
rect 17267 7973 17279 8007
rect 17221 7967 17279 7973
rect 6604 7908 10916 7936
rect 6604 7896 6610 7908
rect 10962 7896 10968 7948
rect 11020 7936 11026 7948
rect 11885 7939 11943 7945
rect 11885 7936 11897 7939
rect 11020 7908 11897 7936
rect 11020 7896 11026 7908
rect 11885 7905 11897 7908
rect 11931 7905 11943 7939
rect 11885 7899 11943 7905
rect 11974 7896 11980 7948
rect 12032 7936 12038 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 12032 7908 12081 7936
rect 12032 7896 12038 7908
rect 12069 7905 12081 7908
rect 12115 7936 12127 7939
rect 13449 7939 13507 7945
rect 13449 7936 13461 7939
rect 12115 7908 13461 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 13449 7905 13461 7908
rect 13495 7936 13507 7939
rect 13630 7936 13636 7948
rect 13495 7908 13636 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 15102 7896 15108 7948
rect 15160 7936 15166 7948
rect 15545 7939 15603 7945
rect 15545 7936 15557 7939
rect 15160 7908 15557 7936
rect 15160 7896 15166 7908
rect 15545 7905 15557 7908
rect 15591 7905 15603 7939
rect 15545 7899 15603 7905
rect 16298 7896 16304 7948
rect 16356 7936 16362 7948
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 16356 7908 17141 7936
rect 16356 7896 16362 7908
rect 17129 7905 17141 7908
rect 17175 7905 17187 7939
rect 17129 7899 17187 7905
rect 17494 7896 17500 7948
rect 17552 7936 17558 7948
rect 17865 7939 17923 7945
rect 17865 7936 17877 7939
rect 17552 7908 17877 7936
rect 17552 7896 17558 7908
rect 17865 7905 17877 7908
rect 17911 7905 17923 7939
rect 18230 7936 18236 7948
rect 18191 7908 18236 7936
rect 17865 7899 17923 7905
rect 18230 7896 18236 7908
rect 18288 7896 18294 7948
rect 4709 7871 4767 7877
rect 3844 7840 4568 7868
rect 3844 7828 3850 7840
rect 4540 7744 4568 7840
rect 4709 7837 4721 7871
rect 4755 7868 4767 7871
rect 4890 7868 4896 7880
rect 4755 7840 4896 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7868 8171 7871
rect 8202 7868 8208 7880
rect 8159 7840 8208 7868
rect 8159 7837 8171 7840
rect 8113 7831 8171 7837
rect 1854 7732 1860 7744
rect 1815 7704 1860 7732
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2038 7732 2044 7744
rect 1999 7704 2044 7732
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2225 7735 2283 7741
rect 2225 7701 2237 7735
rect 2271 7732 2283 7735
rect 2314 7732 2320 7744
rect 2271 7704 2320 7732
rect 2271 7701 2283 7704
rect 2225 7695 2283 7701
rect 2314 7692 2320 7704
rect 2372 7692 2378 7744
rect 2406 7692 2412 7744
rect 2464 7732 2470 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 2464 7704 4077 7732
rect 2464 7692 2470 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4065 7695 4123 7701
rect 4522 7692 4528 7744
rect 4580 7732 4586 7744
rect 5460 7732 5488 7831
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 8754 7868 8760 7880
rect 8628 7840 8760 7868
rect 8628 7828 8634 7840
rect 8754 7828 8760 7840
rect 8812 7868 8818 7880
rect 8849 7871 8907 7877
rect 8849 7868 8861 7871
rect 8812 7840 8861 7868
rect 8812 7828 8818 7840
rect 8849 7837 8861 7840
rect 8895 7837 8907 7871
rect 8849 7831 8907 7837
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 10042 7868 10048 7880
rect 9824 7840 10048 7868
rect 9824 7828 9830 7840
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10226 7868 10232 7880
rect 10187 7840 10232 7868
rect 10226 7828 10232 7840
rect 10284 7828 10290 7880
rect 12158 7868 12164 7880
rect 11256 7840 12164 7868
rect 6730 7760 6736 7812
rect 6788 7800 6794 7812
rect 6788 7772 10088 7800
rect 6788 7760 6794 7772
rect 7101 7735 7159 7741
rect 7101 7732 7113 7735
rect 4580 7704 7113 7732
rect 4580 7692 4586 7704
rect 7101 7701 7113 7704
rect 7147 7701 7159 7735
rect 7466 7732 7472 7744
rect 7427 7704 7472 7732
rect 7101 7695 7159 7701
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 9674 7732 9680 7744
rect 8720 7704 9680 7732
rect 8720 7692 8726 7704
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10060 7732 10088 7772
rect 11256 7732 11284 7840
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 12492 7840 12725 7868
rect 12492 7828 12498 7840
rect 12713 7837 12725 7840
rect 12759 7868 12771 7871
rect 12986 7868 12992 7880
rect 12759 7840 12992 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 13538 7828 13544 7880
rect 13596 7868 13602 7880
rect 13596 7840 13689 7868
rect 13596 7828 13602 7840
rect 14918 7828 14924 7880
rect 14976 7868 14982 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 14976 7840 15301 7868
rect 14976 7828 14982 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 17218 7828 17224 7880
rect 17276 7868 17282 7880
rect 17313 7871 17371 7877
rect 17313 7868 17325 7871
rect 17276 7840 17325 7868
rect 17276 7828 17282 7840
rect 17313 7837 17325 7840
rect 17359 7837 17371 7871
rect 17313 7831 17371 7837
rect 11606 7760 11612 7812
rect 11664 7800 11670 7812
rect 13556 7800 13584 7828
rect 11664 7772 13584 7800
rect 11664 7760 11670 7772
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 16761 7803 16819 7809
rect 16761 7800 16773 7803
rect 16632 7772 16773 7800
rect 16632 7760 16638 7772
rect 16761 7769 16773 7772
rect 16807 7769 16819 7803
rect 16761 7763 16819 7769
rect 18049 7803 18107 7809
rect 18049 7769 18061 7803
rect 18095 7800 18107 7803
rect 18506 7800 18512 7812
rect 18095 7772 18512 7800
rect 18095 7769 18107 7772
rect 18049 7763 18107 7769
rect 18506 7760 18512 7772
rect 18564 7760 18570 7812
rect 11698 7732 11704 7744
rect 10060 7704 11284 7732
rect 11659 7704 11704 7732
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 12158 7732 12164 7744
rect 12119 7704 12164 7732
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 12952 7704 13001 7732
rect 12952 7692 12958 7704
rect 12989 7701 13001 7704
rect 13035 7701 13047 7735
rect 17586 7732 17592 7744
rect 17547 7704 17592 7732
rect 12989 7695 13047 7701
rect 17586 7692 17592 7704
rect 17644 7692 17650 7744
rect 18417 7735 18475 7741
rect 18417 7701 18429 7735
rect 18463 7732 18475 7735
rect 18969 7735 19027 7741
rect 18969 7732 18981 7735
rect 18463 7704 18981 7732
rect 18463 7701 18475 7704
rect 18417 7695 18475 7701
rect 18969 7701 18981 7704
rect 19015 7701 19027 7735
rect 18969 7695 19027 7701
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 1670 7488 1676 7540
rect 1728 7528 1734 7540
rect 2130 7528 2136 7540
rect 1728 7500 2136 7528
rect 1728 7488 1734 7500
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 2958 7528 2964 7540
rect 2919 7500 2964 7528
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 3881 7531 3939 7537
rect 3881 7497 3893 7531
rect 3927 7528 3939 7531
rect 4430 7528 4436 7540
rect 3927 7500 4436 7528
rect 3927 7497 3939 7500
rect 3881 7491 3939 7497
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 5534 7528 5540 7540
rect 5495 7500 5540 7528
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 5736 7500 6469 7528
rect 3789 7463 3847 7469
rect 1596 7432 3556 7460
rect 1596 7333 1624 7432
rect 2406 7392 2412 7404
rect 2367 7364 2412 7392
rect 2406 7352 2412 7364
rect 2464 7352 2470 7404
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 2682 7392 2688 7404
rect 2639 7364 2688 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7324 1547 7327
rect 1581 7327 1639 7333
rect 1581 7324 1593 7327
rect 1535 7296 1593 7324
rect 1535 7293 1547 7296
rect 1489 7287 1547 7293
rect 1581 7293 1593 7296
rect 1627 7293 1639 7327
rect 2314 7324 2320 7336
rect 2275 7296 2320 7324
rect 1581 7287 1639 7293
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 3528 7324 3556 7432
rect 3789 7429 3801 7463
rect 3835 7460 3847 7463
rect 5736 7460 5764 7500
rect 6457 7497 6469 7500
rect 6503 7528 6515 7531
rect 6503 7500 6960 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 3835 7432 5764 7460
rect 3835 7429 3847 7432
rect 3789 7423 3847 7429
rect 6270 7420 6276 7472
rect 6328 7460 6334 7472
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 6328 7432 6837 7460
rect 6328 7420 6334 7432
rect 6825 7429 6837 7432
rect 6871 7429 6883 7463
rect 6932 7460 6960 7500
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 9861 7531 9919 7537
rect 9861 7528 9873 7531
rect 8260 7500 9873 7528
rect 8260 7488 8266 7500
rect 9861 7497 9873 7500
rect 9907 7497 9919 7531
rect 11514 7528 11520 7540
rect 9861 7491 9919 7497
rect 9968 7500 11520 7528
rect 6932 7432 8340 7460
rect 6825 7423 6883 7429
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 4522 7392 4528 7404
rect 3651 7364 4528 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 4522 7352 4528 7364
rect 4580 7352 4586 7404
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 5626 7392 5632 7404
rect 5399 7364 5632 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 5626 7352 5632 7364
rect 5684 7392 5690 7404
rect 6086 7392 6092 7404
rect 5684 7364 6092 7392
rect 5684 7352 5690 7364
rect 6086 7352 6092 7364
rect 6144 7352 6150 7404
rect 6638 7392 6644 7404
rect 6599 7364 6644 7392
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 8018 7392 8024 7404
rect 7423 7364 8024 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 8202 7392 8208 7404
rect 8163 7364 8208 7392
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 8312 7392 8340 7432
rect 9876 7392 9904 7491
rect 9968 7472 9996 7500
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 12342 7488 12348 7540
rect 12400 7528 12406 7540
rect 12400 7500 15056 7528
rect 12400 7488 12406 7500
rect 9950 7420 9956 7472
rect 10008 7420 10014 7472
rect 13170 7460 13176 7472
rect 11808 7432 13176 7460
rect 8312 7364 8616 7392
rect 9876 7364 10088 7392
rect 5902 7324 5908 7336
rect 3528 7296 5908 7324
rect 5902 7284 5908 7296
rect 5960 7284 5966 7336
rect 5997 7327 6055 7333
rect 5997 7293 6009 7327
rect 6043 7324 6055 7327
rect 6454 7324 6460 7336
rect 6043 7296 6460 7324
rect 6043 7293 6055 7296
rect 5997 7287 6055 7293
rect 6454 7284 6460 7296
rect 6512 7284 6518 7336
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 7466 7324 7472 7336
rect 7331 7296 7472 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 2038 7216 2044 7268
rect 2096 7256 2102 7268
rect 3421 7259 3479 7265
rect 3421 7256 3433 7259
rect 2096 7228 3433 7256
rect 2096 7216 2102 7228
rect 3421 7225 3433 7228
rect 3467 7256 3479 7259
rect 3789 7259 3847 7265
rect 3789 7256 3801 7259
rect 3467 7228 3801 7256
rect 3467 7225 3479 7228
rect 3421 7219 3479 7225
rect 3789 7225 3801 7228
rect 3835 7225 3847 7259
rect 3789 7219 3847 7225
rect 4154 7216 4160 7268
rect 4212 7256 4218 7268
rect 4249 7259 4307 7265
rect 4249 7256 4261 7259
rect 4212 7228 4261 7256
rect 4212 7216 4218 7228
rect 4249 7225 4261 7228
rect 4295 7256 4307 7259
rect 4614 7256 4620 7268
rect 4295 7228 4620 7256
rect 4295 7225 4307 7228
rect 4249 7219 4307 7225
rect 4614 7216 4620 7228
rect 4672 7216 4678 7268
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5350 7256 5356 7268
rect 5123 7228 5356 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5350 7216 5356 7228
rect 5408 7216 5414 7268
rect 8386 7256 8392 7268
rect 5736 7228 8392 7256
rect 1762 7188 1768 7200
rect 1723 7160 1768 7188
rect 1762 7148 1768 7160
rect 1820 7148 1826 7200
rect 1946 7188 1952 7200
rect 1907 7160 1952 7188
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 2682 7148 2688 7200
rect 2740 7188 2746 7200
rect 2777 7191 2835 7197
rect 2777 7188 2789 7191
rect 2740 7160 2789 7188
rect 2740 7148 2746 7160
rect 2777 7157 2789 7160
rect 2823 7157 2835 7191
rect 3326 7188 3332 7200
rect 3287 7160 3332 7188
rect 2777 7151 2835 7157
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4709 7191 4767 7197
rect 4709 7188 4721 7191
rect 4387 7160 4721 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4709 7157 4721 7160
rect 4755 7157 4767 7191
rect 5166 7188 5172 7200
rect 5127 7160 5172 7188
rect 4709 7151 4767 7157
rect 5166 7148 5172 7160
rect 5224 7188 5230 7200
rect 5736 7188 5764 7228
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 5224 7160 5764 7188
rect 5224 7148 5230 7160
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 5868 7160 5917 7188
rect 5868 7148 5874 7160
rect 5905 7157 5917 7160
rect 5951 7188 5963 7191
rect 6638 7188 6644 7200
rect 5951 7160 6644 7188
rect 5951 7157 5963 7160
rect 5905 7151 5963 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 7193 7191 7251 7197
rect 7193 7157 7205 7191
rect 7239 7188 7251 7191
rect 7653 7191 7711 7197
rect 7653 7188 7665 7191
rect 7239 7160 7665 7188
rect 7239 7157 7251 7160
rect 7193 7151 7251 7157
rect 7653 7157 7665 7160
rect 7699 7157 7711 7191
rect 8018 7188 8024 7200
rect 7979 7160 8024 7188
rect 7653 7151 7711 7157
rect 8018 7148 8024 7160
rect 8076 7148 8082 7200
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 8496 7188 8524 7287
rect 8588 7256 8616 7364
rect 8754 7333 8760 7336
rect 8748 7324 8760 7333
rect 8715 7296 8760 7324
rect 8748 7287 8760 7296
rect 8754 7284 8760 7287
rect 8812 7284 8818 7336
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9732 7296 9965 7324
rect 9732 7284 9738 7296
rect 9953 7293 9965 7296
rect 9999 7293 10011 7327
rect 10060 7324 10088 7364
rect 10209 7327 10267 7333
rect 10209 7324 10221 7327
rect 10060 7296 10221 7324
rect 9953 7287 10011 7293
rect 10209 7293 10221 7296
rect 10255 7293 10267 7327
rect 10209 7287 10267 7293
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 11808 7324 11836 7432
rect 13170 7420 13176 7432
rect 13228 7420 13234 7472
rect 15028 7460 15056 7500
rect 15102 7488 15108 7540
rect 15160 7528 15166 7540
rect 15197 7531 15255 7537
rect 15197 7528 15209 7531
rect 15160 7500 15209 7528
rect 15160 7488 15166 7500
rect 15197 7497 15209 7500
rect 15243 7497 15255 7531
rect 15197 7491 15255 7497
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 15841 7531 15899 7537
rect 15841 7528 15853 7531
rect 15528 7500 15853 7528
rect 15528 7488 15534 7500
rect 15841 7497 15853 7500
rect 15887 7528 15899 7531
rect 15933 7531 15991 7537
rect 15933 7528 15945 7531
rect 15887 7500 15945 7528
rect 15887 7497 15899 7500
rect 15841 7491 15899 7497
rect 15933 7497 15945 7500
rect 15979 7497 15991 7531
rect 16482 7528 16488 7540
rect 16443 7500 16488 7528
rect 15933 7491 15991 7497
rect 16482 7488 16488 7500
rect 16540 7488 16546 7540
rect 16301 7463 16359 7469
rect 16301 7460 16313 7463
rect 15028 7432 16313 7460
rect 16301 7429 16313 7432
rect 16347 7460 16359 7463
rect 17034 7460 17040 7472
rect 16347 7432 17040 7460
rect 16347 7429 16359 7432
rect 16301 7423 16359 7429
rect 17034 7420 17040 7432
rect 17092 7460 17098 7472
rect 18230 7460 18236 7472
rect 17092 7432 18236 7460
rect 17092 7420 17098 7432
rect 18230 7420 18236 7432
rect 18288 7460 18294 7472
rect 18417 7463 18475 7469
rect 18417 7460 18429 7463
rect 18288 7432 18429 7460
rect 18288 7420 18294 7432
rect 18417 7429 18429 7432
rect 18463 7429 18475 7463
rect 18417 7423 18475 7429
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7392 12127 7395
rect 12342 7392 12348 7404
rect 12115 7364 12348 7392
rect 12115 7361 12127 7364
rect 12069 7355 12127 7361
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 12894 7392 12900 7404
rect 12855 7364 12900 7392
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 15841 7395 15899 7401
rect 13044 7364 13089 7392
rect 13044 7352 13050 7364
rect 15841 7361 15853 7395
rect 15887 7392 15899 7395
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 15887 7364 16957 7392
rect 15887 7361 15899 7364
rect 15841 7355 15899 7361
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17310 7392 17316 7404
rect 17175 7364 17316 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17310 7352 17316 7364
rect 17368 7352 17374 7404
rect 10560 7296 11836 7324
rect 11885 7327 11943 7333
rect 10560 7284 10566 7296
rect 11885 7293 11897 7327
rect 11931 7324 11943 7327
rect 11931 7296 12480 7324
rect 11931 7293 11943 7296
rect 11885 7287 11943 7293
rect 10778 7256 10784 7268
rect 8588 7228 10784 7256
rect 10778 7216 10784 7228
rect 10836 7216 10842 7268
rect 11977 7259 12035 7265
rect 11977 7225 11989 7259
rect 12023 7256 12035 7259
rect 12158 7256 12164 7268
rect 12023 7228 12164 7256
rect 12023 7225 12035 7228
rect 11977 7219 12035 7225
rect 12158 7216 12164 7228
rect 12216 7216 12222 7268
rect 9674 7188 9680 7200
rect 8168 7160 8213 7188
rect 8496 7160 9680 7188
rect 8168 7148 8174 7160
rect 9674 7148 9680 7160
rect 9732 7188 9738 7200
rect 10226 7188 10232 7200
rect 9732 7160 10232 7188
rect 9732 7148 9738 7160
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 10468 7160 11345 7188
rect 10468 7148 10474 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11514 7188 11520 7200
rect 11475 7160 11520 7188
rect 11333 7151 11391 7157
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 12452 7197 12480 7296
rect 12710 7284 12716 7336
rect 12768 7324 12774 7336
rect 13004 7324 13032 7352
rect 12768 7296 13032 7324
rect 13817 7327 13875 7333
rect 12768 7284 12774 7296
rect 13817 7293 13829 7327
rect 13863 7324 13875 7327
rect 13906 7324 13912 7336
rect 13863 7296 13912 7324
rect 13863 7293 13875 7296
rect 13817 7287 13875 7293
rect 13906 7284 13912 7296
rect 13964 7284 13970 7336
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 15654 7324 15660 7336
rect 14700 7296 15660 7324
rect 14700 7284 14706 7296
rect 15654 7284 15660 7296
rect 15712 7324 15718 7336
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 15712 7296 16129 7324
rect 15712 7284 15718 7296
rect 16117 7293 16129 7296
rect 16163 7324 16175 7327
rect 17218 7324 17224 7336
rect 16163 7296 17224 7324
rect 16163 7293 16175 7296
rect 16117 7287 16175 7293
rect 17218 7284 17224 7296
rect 17276 7284 17282 7336
rect 17586 7324 17592 7336
rect 17547 7296 17592 7324
rect 17586 7284 17592 7296
rect 17644 7284 17650 7336
rect 17954 7284 17960 7336
rect 18012 7324 18018 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 18012 7296 18061 7324
rect 18012 7284 18018 7296
rect 18049 7293 18061 7296
rect 18095 7324 18107 7327
rect 18414 7324 18420 7336
rect 18095 7296 18420 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18414 7284 18420 7296
rect 18472 7284 18478 7336
rect 12802 7256 12808 7268
rect 12715 7228 12808 7256
rect 12802 7216 12808 7228
rect 12860 7256 12866 7268
rect 14084 7259 14142 7265
rect 12860 7228 13676 7256
rect 12860 7216 12866 7228
rect 13648 7200 13676 7228
rect 14084 7225 14096 7259
rect 14130 7256 14142 7259
rect 16666 7256 16672 7268
rect 14130 7228 16672 7256
rect 14130 7225 14142 7228
rect 14084 7219 14142 7225
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 16853 7259 16911 7265
rect 16853 7225 16865 7259
rect 16899 7256 16911 7259
rect 17313 7259 17371 7265
rect 17313 7256 17325 7259
rect 16899 7228 17325 7256
rect 16899 7225 16911 7228
rect 16853 7219 16911 7225
rect 17313 7225 17325 7228
rect 17359 7225 17371 7259
rect 17313 7219 17371 7225
rect 12437 7191 12495 7197
rect 12437 7157 12449 7191
rect 12483 7157 12495 7191
rect 12437 7151 12495 7157
rect 13265 7191 13323 7197
rect 13265 7157 13277 7191
rect 13311 7188 13323 7191
rect 13354 7188 13360 7200
rect 13311 7160 13360 7188
rect 13311 7157 13323 7160
rect 13265 7151 13323 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 13630 7188 13636 7200
rect 13591 7160 13636 7188
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13722 7148 13728 7200
rect 13780 7188 13786 7200
rect 17586 7188 17592 7200
rect 13780 7160 17592 7188
rect 13780 7148 13786 7160
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 17770 7188 17776 7200
rect 17731 7160 17776 7188
rect 17770 7148 17776 7160
rect 17828 7148 17834 7200
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 18233 7191 18291 7197
rect 18233 7188 18245 7191
rect 17920 7160 18245 7188
rect 17920 7148 17926 7160
rect 18233 7157 18245 7160
rect 18279 7157 18291 7191
rect 18233 7151 18291 7157
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 18966 7052 18972 7064
rect 1104 7024 18860 7046
rect 18927 7024 18972 7052
rect 18966 7012 18972 7024
rect 19024 7012 19030 7064
rect 2682 6944 2688 6996
rect 2740 6984 2746 6996
rect 3326 6984 3332 6996
rect 2740 6956 3188 6984
rect 3287 6956 3332 6984
rect 2740 6944 2746 6956
rect 2498 6876 2504 6928
rect 2556 6916 2562 6928
rect 3160 6916 3188 6956
rect 3326 6944 3332 6956
rect 3384 6944 3390 6996
rect 4157 6987 4215 6993
rect 4157 6953 4169 6987
rect 4203 6984 4215 6987
rect 4338 6984 4344 6996
rect 4203 6956 4344 6984
rect 4203 6953 4215 6956
rect 4157 6947 4215 6953
rect 4338 6944 4344 6956
rect 4396 6984 4402 6996
rect 5166 6984 5172 6996
rect 4396 6956 5172 6984
rect 4396 6944 4402 6956
rect 5166 6944 5172 6956
rect 5224 6944 5230 6996
rect 5626 6984 5632 6996
rect 5587 6956 5632 6984
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 5813 6987 5871 6993
rect 5813 6953 5825 6987
rect 5859 6984 5871 6987
rect 6454 6984 6460 6996
rect 5859 6956 6460 6984
rect 5859 6953 5871 6956
rect 5813 6947 5871 6953
rect 6454 6944 6460 6956
rect 6512 6944 6518 6996
rect 8110 6984 8116 6996
rect 8071 6956 8116 6984
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 10502 6984 10508 6996
rect 8220 6956 10508 6984
rect 2556 6888 2820 6916
rect 3160 6888 5304 6916
rect 2556 6876 2562 6888
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6817 1731 6851
rect 1673 6811 1731 6817
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6817 2099 6851
rect 2041 6811 2099 6817
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2682 6848 2688 6860
rect 2455 6820 2688 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 1688 6712 1716 6811
rect 2056 6780 2084 6811
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 2792 6857 2820 6888
rect 2777 6851 2835 6857
rect 2777 6817 2789 6851
rect 2823 6817 2835 6851
rect 2777 6811 2835 6817
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6848 3847 6851
rect 4154 6848 4160 6860
rect 3835 6820 4160 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4522 6857 4528 6860
rect 4516 6848 4528 6857
rect 4483 6820 4528 6848
rect 4516 6811 4528 6820
rect 4522 6808 4528 6811
rect 4580 6808 4586 6860
rect 2056 6752 2912 6780
rect 2038 6712 2044 6724
rect 1627 6684 2044 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2038 6672 2044 6684
rect 2096 6672 2102 6724
rect 2222 6712 2228 6724
rect 2183 6684 2228 6712
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 2593 6715 2651 6721
rect 2593 6681 2605 6715
rect 2639 6712 2651 6715
rect 2774 6712 2780 6724
rect 2639 6684 2780 6712
rect 2639 6681 2651 6684
rect 2593 6675 2651 6681
rect 2774 6672 2780 6684
rect 2832 6672 2838 6724
rect 1854 6644 1860 6656
rect 1815 6616 1860 6644
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 2884 6644 2912 6752
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 4249 6783 4307 6789
rect 4249 6780 4261 6783
rect 3752 6752 4261 6780
rect 3752 6740 3758 6752
rect 4249 6749 4261 6752
rect 4295 6749 4307 6783
rect 5276 6780 5304 6888
rect 5350 6876 5356 6928
rect 5408 6916 5414 6928
rect 7009 6919 7067 6925
rect 7009 6916 7021 6919
rect 5408 6888 7021 6916
rect 5408 6876 5414 6888
rect 7009 6885 7021 6888
rect 7055 6916 7067 6919
rect 8220 6916 8248 6956
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 10594 6944 10600 6996
rect 10652 6984 10658 6996
rect 13354 6984 13360 6996
rect 10652 6956 13216 6984
rect 13315 6956 13360 6984
rect 10652 6944 10658 6956
rect 7055 6888 8248 6916
rect 7055 6885 7067 6888
rect 7009 6879 7067 6885
rect 8386 6876 8392 6928
rect 8444 6916 8450 6928
rect 11974 6916 11980 6928
rect 8444 6888 11980 6916
rect 8444 6876 8450 6888
rect 11974 6876 11980 6888
rect 12032 6876 12038 6928
rect 12434 6916 12440 6928
rect 12268 6888 12440 6916
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 6086 6848 6092 6860
rect 5500 6820 6092 6848
rect 5500 6808 5506 6820
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6848 6331 6851
rect 6822 6848 6828 6860
rect 6319 6820 6828 6848
rect 6319 6817 6331 6820
rect 6273 6811 6331 6817
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8478 6848 8484 6860
rect 8067 6820 8484 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 10594 6848 10600 6860
rect 9048 6820 10600 6848
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 5276 6752 6377 6780
rect 4249 6743 4307 6749
rect 6365 6749 6377 6752
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 2961 6715 3019 6721
rect 2961 6681 2973 6715
rect 3007 6712 3019 6715
rect 3326 6712 3332 6724
rect 3007 6684 3332 6712
rect 3007 6681 3019 6684
rect 2961 6675 3019 6681
rect 3326 6672 3332 6684
rect 3384 6672 3390 6724
rect 3234 6644 3240 6656
rect 2884 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 4264 6644 4292 6743
rect 5350 6672 5356 6724
rect 5408 6712 5414 6724
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 5408 6684 5917 6712
rect 5408 6672 5414 6684
rect 5905 6681 5917 6684
rect 5951 6681 5963 6715
rect 6380 6712 6408 6743
rect 6454 6740 6460 6792
rect 6512 6780 6518 6792
rect 6730 6780 6736 6792
rect 6512 6752 6557 6780
rect 6691 6752 6736 6780
rect 6512 6740 6518 6752
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 8570 6780 8576 6792
rect 7984 6752 8576 6780
rect 7984 6740 7990 6752
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 8754 6780 8760 6792
rect 8715 6752 8760 6780
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 8938 6780 8944 6792
rect 8899 6752 8944 6780
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 6748 6712 6776 6740
rect 6380 6684 6776 6712
rect 5905 6675 5963 6681
rect 7006 6672 7012 6724
rect 7064 6712 7070 6724
rect 9048 6712 9076 6820
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 10772 6851 10830 6857
rect 10772 6817 10784 6851
rect 10818 6848 10830 6851
rect 12268 6848 12296 6888
rect 12434 6876 12440 6888
rect 12492 6876 12498 6928
rect 13188 6916 13216 6956
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 13449 6987 13507 6993
rect 13449 6953 13461 6987
rect 13495 6984 13507 6987
rect 13538 6984 13544 6996
rect 13495 6956 13544 6984
rect 13495 6953 13507 6956
rect 13449 6947 13507 6953
rect 13538 6944 13544 6956
rect 13596 6984 13602 6996
rect 13909 6987 13967 6993
rect 13909 6984 13921 6987
rect 13596 6956 13921 6984
rect 13596 6944 13602 6956
rect 13909 6953 13921 6956
rect 13955 6984 13967 6987
rect 16114 6984 16120 6996
rect 13955 6956 16120 6984
rect 13955 6953 13967 6956
rect 13909 6947 13967 6953
rect 16114 6944 16120 6956
rect 16172 6944 16178 6996
rect 16482 6944 16488 6996
rect 16540 6984 16546 6996
rect 17957 6987 18015 6993
rect 17957 6984 17969 6987
rect 16540 6956 17969 6984
rect 16540 6944 16546 6956
rect 17957 6953 17969 6956
rect 18003 6953 18015 6987
rect 18414 6984 18420 6996
rect 18375 6956 18420 6984
rect 17957 6947 18015 6953
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 14642 6916 14648 6928
rect 13188 6888 14648 6916
rect 14642 6876 14648 6888
rect 14700 6876 14706 6928
rect 14737 6919 14795 6925
rect 14737 6885 14749 6919
rect 14783 6916 14795 6919
rect 17218 6916 17224 6928
rect 14783 6888 16252 6916
rect 17179 6888 17224 6916
rect 14783 6885 14795 6888
rect 14737 6879 14795 6885
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 10818 6820 12296 6848
rect 12452 6820 12541 6848
rect 10818 6817 10830 6820
rect 10772 6811 10830 6817
rect 10502 6780 10508 6792
rect 10463 6752 10508 6780
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11848 6752 11989 6780
rect 11848 6740 11854 6752
rect 11977 6749 11989 6752
rect 12023 6780 12035 6783
rect 12452 6780 12480 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 12529 6811 12587 6817
rect 12728 6820 13584 6848
rect 12728 6792 12756 6820
rect 12618 6780 12624 6792
rect 12023 6752 12480 6780
rect 12579 6752 12624 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 13556 6789 13584 6820
rect 14660 6820 15301 6848
rect 13541 6783 13599 6789
rect 12768 6752 12813 6780
rect 12768 6740 12774 6752
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 14660 6780 14688 6820
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15556 6851 15614 6857
rect 15556 6817 15568 6851
rect 15602 6848 15614 6851
rect 16114 6848 16120 6860
rect 15602 6820 16120 6848
rect 15602 6817 15614 6820
rect 15556 6811 15614 6817
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 16224 6848 16252 6888
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 16224 6820 16344 6848
rect 14056 6752 14688 6780
rect 14829 6783 14887 6789
rect 14056 6740 14062 6752
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 14918 6780 14924 6792
rect 14875 6752 14924 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15013 6783 15071 6789
rect 15013 6749 15025 6783
rect 15059 6780 15071 6783
rect 15102 6780 15108 6792
rect 15059 6752 15108 6780
rect 15059 6749 15071 6752
rect 15013 6743 15071 6749
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 9950 6712 9956 6724
rect 7064 6684 9076 6712
rect 9232 6684 9956 6712
rect 7064 6672 7070 6684
rect 5534 6644 5540 6656
rect 4264 6616 5540 6644
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 9232 6653 9260 6684
rect 9950 6672 9956 6684
rect 10008 6672 10014 6724
rect 14369 6715 14427 6721
rect 14369 6712 14381 6715
rect 11716 6684 14381 6712
rect 9217 6647 9275 6653
rect 9217 6644 9229 6647
rect 8628 6616 9229 6644
rect 8628 6604 8634 6616
rect 9217 6613 9229 6616
rect 9263 6613 9275 6647
rect 9217 6607 9275 6613
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 11716 6644 11744 6684
rect 14369 6681 14381 6684
rect 14415 6681 14427 6715
rect 14369 6675 14427 6681
rect 11882 6644 11888 6656
rect 9548 6616 11744 6644
rect 11843 6616 11888 6644
rect 9548 6604 9554 6616
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 12158 6644 12164 6656
rect 12119 6616 12164 6644
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 12989 6647 13047 6653
rect 12989 6644 13001 6647
rect 12860 6616 13001 6644
rect 12860 6604 12866 6616
rect 12989 6613 13001 6616
rect 13035 6613 13047 6647
rect 16316 6644 16344 6820
rect 17034 6808 17040 6860
rect 17092 6848 17098 6860
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 17092 6820 17141 6848
rect 17092 6808 17098 6820
rect 17129 6817 17141 6820
rect 17175 6817 17187 6851
rect 17129 6811 17187 6817
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 17460 6820 18184 6848
rect 17460 6808 17466 6820
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 18156 6789 18184 6820
rect 18049 6783 18107 6789
rect 17368 6752 17413 6780
rect 17368 6740 17374 6752
rect 18049 6749 18061 6783
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6749 18199 6783
rect 18141 6743 18199 6749
rect 16666 6712 16672 6724
rect 16627 6684 16672 6712
rect 16666 6672 16672 6684
rect 16724 6672 16730 6724
rect 16761 6715 16819 6721
rect 16761 6681 16773 6715
rect 16807 6712 16819 6715
rect 18064 6712 18092 6743
rect 16807 6684 18092 6712
rect 16807 6681 16819 6684
rect 16761 6675 16819 6681
rect 17589 6647 17647 6653
rect 17589 6644 17601 6647
rect 16316 6616 17601 6644
rect 12989 6607 13047 6613
rect 17589 6613 17601 6616
rect 17635 6613 17647 6647
rect 17589 6607 17647 6613
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1627 6412 3188 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1688 6245 1716 6412
rect 3160 6372 3188 6412
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 6638 6440 6644 6452
rect 3292 6412 4660 6440
rect 6551 6412 6644 6440
rect 3292 6400 3298 6412
rect 3602 6372 3608 6384
rect 3160 6344 3608 6372
rect 3602 6332 3608 6344
rect 3660 6332 3666 6384
rect 4632 6372 4660 6412
rect 6638 6400 6644 6412
rect 6696 6440 6702 6452
rect 7006 6440 7012 6452
rect 6696 6412 7012 6440
rect 6696 6400 6702 6412
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 8076 6412 8125 6440
rect 8076 6400 8082 6412
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 13538 6440 13544 6452
rect 8113 6403 8171 6409
rect 8220 6412 13544 6440
rect 8220 6372 8248 6412
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 14918 6400 14924 6452
rect 14976 6440 14982 6452
rect 16853 6443 16911 6449
rect 16853 6440 16865 6443
rect 14976 6412 16865 6440
rect 14976 6400 14982 6412
rect 16853 6409 16865 6412
rect 16899 6409 16911 6443
rect 17770 6440 17776 6452
rect 17683 6412 17776 6440
rect 16853 6403 16911 6409
rect 17770 6400 17776 6412
rect 17828 6440 17834 6452
rect 18598 6440 18604 6452
rect 17828 6412 18604 6440
rect 17828 6400 17834 6412
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 4632 6344 8248 6372
rect 8312 6344 8892 6372
rect 2038 6264 2044 6316
rect 2096 6304 2102 6316
rect 2096 6276 2268 6304
rect 2096 6264 2102 6276
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6205 1731 6239
rect 1673 6199 1731 6205
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6205 2191 6239
rect 2240 6236 2268 6276
rect 3344 6276 3740 6304
rect 3344 6236 3372 6276
rect 3602 6236 3608 6248
rect 2240 6208 3372 6236
rect 3436 6208 3608 6236
rect 2133 6199 2191 6205
rect 1854 6100 1860 6112
rect 1815 6072 1860 6100
rect 1854 6060 1860 6072
rect 1912 6060 1918 6112
rect 2148 6100 2176 6199
rect 2400 6171 2458 6177
rect 2400 6137 2412 6171
rect 2446 6168 2458 6171
rect 3234 6168 3240 6180
rect 2446 6140 3240 6168
rect 2446 6137 2458 6140
rect 2400 6131 2458 6137
rect 3234 6128 3240 6140
rect 3292 6128 3298 6180
rect 3436 6100 3464 6208
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 3712 6236 3740 6276
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 6273 6307 6331 6313
rect 6273 6304 6285 6307
rect 4764 6276 6285 6304
rect 4764 6264 4770 6276
rect 6273 6273 6285 6276
rect 6319 6304 6331 6307
rect 6454 6304 6460 6316
rect 6319 6276 6460 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 6822 6304 6828 6316
rect 6783 6276 6828 6304
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 8312 6304 8340 6344
rect 8754 6304 8760 6316
rect 7616 6276 8340 6304
rect 8715 6276 8760 6304
rect 7616 6264 7622 6276
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 8864 6304 8892 6344
rect 9674 6332 9680 6384
rect 9732 6372 9738 6384
rect 10137 6375 10195 6381
rect 10137 6372 10149 6375
rect 9732 6344 10149 6372
rect 9732 6332 9738 6344
rect 10137 6341 10149 6344
rect 10183 6372 10195 6375
rect 10502 6372 10508 6384
rect 10183 6344 10508 6372
rect 10183 6341 10195 6344
rect 10137 6335 10195 6341
rect 10502 6332 10508 6344
rect 10560 6372 10566 6384
rect 10560 6344 10916 6372
rect 10560 6332 10566 6344
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 8864 6276 9781 6304
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 10888 6248 10916 6344
rect 11882 6332 11888 6384
rect 11940 6372 11946 6384
rect 12342 6372 12348 6384
rect 11940 6344 12348 6372
rect 11940 6332 11946 6344
rect 12342 6332 12348 6344
rect 12400 6372 12406 6384
rect 15289 6375 15347 6381
rect 12400 6344 13032 6372
rect 12400 6332 12406 6344
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 13004 6313 13032 6344
rect 15289 6341 15301 6375
rect 15335 6372 15347 6375
rect 16114 6372 16120 6384
rect 15335 6344 16120 6372
rect 15335 6341 15347 6344
rect 15289 6335 15347 6341
rect 16114 6332 16120 6344
rect 16172 6372 16178 6384
rect 17310 6372 17316 6384
rect 16172 6344 17316 6372
rect 16172 6332 16178 6344
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12216 6276 12909 6304
rect 12216 6264 12222 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6273 13047 6307
rect 13354 6304 13360 6316
rect 13315 6276 13360 6304
rect 12989 6267 13047 6273
rect 13354 6264 13360 6276
rect 13412 6264 13418 6316
rect 13906 6304 13912 6316
rect 13867 6276 13912 6304
rect 13906 6264 13912 6276
rect 13964 6264 13970 6316
rect 16482 6264 16488 6316
rect 16540 6304 16546 6316
rect 16592 6313 16620 6344
rect 17310 6332 17316 6344
rect 17368 6332 17374 6384
rect 16577 6307 16635 6313
rect 16577 6304 16589 6307
rect 16540 6276 16589 6304
rect 16540 6264 16546 6276
rect 16577 6273 16589 6276
rect 16623 6273 16635 6307
rect 16577 6267 16635 6273
rect 16666 6264 16672 6316
rect 16724 6304 16730 6316
rect 17402 6304 17408 6316
rect 16724 6276 17408 6304
rect 16724 6264 16730 6276
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 8481 6239 8539 6245
rect 3712 6208 8156 6236
rect 3786 6128 3792 6180
rect 3844 6177 3850 6180
rect 3844 6171 3908 6177
rect 3844 6137 3862 6171
rect 3896 6137 3908 6171
rect 3844 6131 3908 6137
rect 5629 6171 5687 6177
rect 5629 6137 5641 6171
rect 5675 6168 5687 6171
rect 5675 6140 5856 6168
rect 5675 6137 5687 6140
rect 5629 6131 5687 6137
rect 3844 6128 3850 6131
rect 2148 6072 3464 6100
rect 3513 6103 3571 6109
rect 3513 6069 3525 6103
rect 3559 6100 3571 6103
rect 3804 6100 3832 6128
rect 3559 6072 3832 6100
rect 3559 6069 3571 6072
rect 3513 6063 3571 6069
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 4985 6103 5043 6109
rect 4985 6100 4997 6103
rect 4580 6072 4997 6100
rect 4580 6060 4586 6072
rect 4985 6069 4997 6072
rect 5031 6069 5043 6103
rect 5718 6100 5724 6112
rect 5679 6072 5724 6100
rect 4985 6063 5043 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 5828 6100 5856 6140
rect 5902 6128 5908 6180
rect 5960 6168 5966 6180
rect 6181 6171 6239 6177
rect 6181 6168 6193 6171
rect 5960 6140 6193 6168
rect 5960 6128 5966 6140
rect 6181 6137 6193 6140
rect 6227 6168 6239 6171
rect 6638 6168 6644 6180
rect 6227 6140 6644 6168
rect 6227 6137 6239 6140
rect 6181 6131 6239 6137
rect 6638 6128 6644 6140
rect 6696 6128 6702 6180
rect 8128 6168 8156 6208
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 8938 6236 8944 6248
rect 8527 6208 8944 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 9490 6236 9496 6248
rect 9451 6208 9496 6236
rect 9490 6196 9496 6208
rect 9548 6196 9554 6248
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6236 10379 6239
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10367 6208 10793 6236
rect 10367 6205 10379 6208
rect 10321 6199 10379 6205
rect 10781 6205 10793 6208
rect 10827 6205 10839 6239
rect 10781 6199 10839 6205
rect 10870 6196 10876 6248
rect 10928 6236 10934 6248
rect 11140 6239 11198 6245
rect 10928 6208 10973 6236
rect 10928 6196 10934 6208
rect 11140 6205 11152 6239
rect 11186 6236 11198 6239
rect 11882 6236 11888 6248
rect 11186 6208 11888 6236
rect 11186 6205 11198 6208
rect 11140 6199 11198 6205
rect 11882 6196 11888 6208
rect 11940 6196 11946 6248
rect 12802 6236 12808 6248
rect 12763 6208 12808 6236
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 15838 6196 15844 6248
rect 15896 6236 15902 6248
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 15896 6208 17325 6236
rect 15896 6196 15902 6208
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 18046 6236 18052 6248
rect 18007 6208 18052 6236
rect 17313 6199 17371 6205
rect 18046 6196 18052 6208
rect 18104 6236 18110 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 18104 6208 18429 6236
rect 18104 6196 18110 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 8573 6171 8631 6177
rect 8573 6168 8585 6171
rect 8128 6140 8585 6168
rect 8573 6137 8585 6140
rect 8619 6168 8631 6171
rect 9033 6171 9091 6177
rect 9033 6168 9045 6171
rect 8619 6140 9045 6168
rect 8619 6137 8631 6140
rect 8573 6131 8631 6137
rect 9033 6137 9045 6140
rect 9079 6168 9091 6171
rect 9079 6140 13860 6168
rect 9079 6137 9091 6140
rect 9033 6131 9091 6137
rect 6089 6103 6147 6109
rect 6089 6100 6101 6103
rect 5828 6072 6101 6100
rect 6089 6069 6101 6072
rect 6135 6100 6147 6103
rect 6546 6100 6552 6112
rect 6135 6072 6552 6100
rect 6135 6069 6147 6072
rect 6089 6063 6147 6069
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 10781 6103 10839 6109
rect 10781 6069 10793 6103
rect 10827 6100 10839 6103
rect 11698 6100 11704 6112
rect 10827 6072 11704 6100
rect 10827 6069 10839 6072
rect 10781 6063 10839 6069
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 12342 6100 12348 6112
rect 12299 6072 12348 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 13832 6100 13860 6140
rect 13998 6128 14004 6180
rect 14056 6168 14062 6180
rect 14154 6171 14212 6177
rect 14154 6168 14166 6171
rect 14056 6140 14166 6168
rect 14056 6128 14062 6140
rect 14154 6137 14166 6140
rect 14200 6137 14212 6171
rect 17221 6171 17279 6177
rect 17221 6168 17233 6171
rect 14154 6131 14212 6137
rect 16040 6140 17233 6168
rect 15286 6100 15292 6112
rect 12492 6072 12537 6100
rect 13832 6072 15292 6100
rect 12492 6060 12498 6072
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 15746 6060 15752 6112
rect 15804 6100 15810 6112
rect 15841 6103 15899 6109
rect 15841 6100 15853 6103
rect 15804 6072 15853 6100
rect 15804 6060 15810 6072
rect 15841 6069 15853 6072
rect 15887 6100 15899 6103
rect 15930 6100 15936 6112
rect 15887 6072 15936 6100
rect 15887 6069 15899 6072
rect 15841 6063 15899 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16040 6109 16068 6140
rect 17221 6137 17233 6140
rect 17267 6137 17279 6171
rect 17221 6131 17279 6137
rect 16025 6103 16083 6109
rect 16025 6069 16037 6103
rect 16071 6069 16083 6103
rect 16025 6063 16083 6069
rect 16114 6060 16120 6112
rect 16172 6100 16178 6112
rect 16393 6103 16451 6109
rect 16393 6100 16405 6103
rect 16172 6072 16405 6100
rect 16172 6060 16178 6072
rect 16393 6069 16405 6072
rect 16439 6069 16451 6103
rect 16393 6063 16451 6069
rect 16485 6103 16543 6109
rect 16485 6069 16497 6103
rect 16531 6100 16543 6103
rect 16574 6100 16580 6112
rect 16531 6072 16580 6100
rect 16531 6069 16543 6072
rect 16485 6063 16543 6069
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 18230 6100 18236 6112
rect 18191 6072 18236 6100
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 2590 5896 2596 5908
rect 2551 5868 2596 5896
rect 2590 5856 2596 5868
rect 2648 5856 2654 5908
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 3418 5896 3424 5908
rect 2832 5868 3424 5896
rect 2832 5856 2838 5868
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 4157 5899 4215 5905
rect 4157 5896 4169 5899
rect 3559 5868 4169 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 4157 5865 4169 5868
rect 4203 5865 4215 5899
rect 4157 5859 4215 5865
rect 4985 5899 5043 5905
rect 4985 5865 4997 5899
rect 5031 5896 5043 5899
rect 5074 5896 5080 5908
rect 5031 5868 5080 5896
rect 5031 5865 5043 5868
rect 4985 5859 5043 5865
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 5350 5896 5356 5908
rect 5311 5868 5356 5896
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5445 5899 5503 5905
rect 5445 5865 5457 5899
rect 5491 5896 5503 5899
rect 5718 5896 5724 5908
rect 5491 5868 5724 5896
rect 5491 5865 5503 5868
rect 5445 5859 5503 5865
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 5813 5899 5871 5905
rect 5813 5865 5825 5899
rect 5859 5865 5871 5899
rect 7374 5896 7380 5908
rect 5813 5859 5871 5865
rect 7024 5868 7380 5896
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5760 2099 5763
rect 2608 5760 2636 5856
rect 2682 5788 2688 5840
rect 2740 5828 2746 5840
rect 2740 5800 2912 5828
rect 2740 5788 2746 5800
rect 2087 5732 2636 5760
rect 2087 5729 2099 5732
rect 2041 5723 2099 5729
rect 1688 5692 1716 5723
rect 2501 5695 2559 5701
rect 2501 5692 2513 5695
rect 1688 5664 2513 5692
rect 2501 5661 2513 5664
rect 2547 5692 2559 5695
rect 2774 5692 2780 5704
rect 2547 5664 2780 5692
rect 2547 5661 2559 5664
rect 2501 5655 2559 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 2884 5633 2912 5800
rect 3234 5788 3240 5840
rect 3292 5828 3298 5840
rect 4065 5831 4123 5837
rect 4065 5828 4077 5831
rect 3292 5800 4077 5828
rect 3292 5788 3298 5800
rect 4065 5797 4077 5800
rect 4111 5797 4123 5831
rect 4525 5831 4583 5837
rect 4525 5828 4537 5831
rect 4065 5791 4123 5797
rect 4356 5800 4537 5828
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 3142 5760 3148 5772
rect 3099 5732 3148 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 3142 5720 3148 5732
rect 3200 5760 3206 5772
rect 4356 5760 4384 5800
rect 4525 5797 4537 5800
rect 4571 5828 4583 5831
rect 4571 5800 5120 5828
rect 4571 5797 4583 5800
rect 4525 5791 4583 5797
rect 5092 5760 5120 5800
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 5828 5828 5856 5859
rect 5592 5800 5856 5828
rect 5592 5788 5598 5800
rect 5997 5763 6055 5769
rect 3200 5732 4384 5760
rect 4448 5732 4752 5760
rect 5092 5732 5672 5760
rect 3200 5720 3206 5732
rect 3602 5692 3608 5704
rect 3563 5664 3608 5692
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 3786 5692 3792 5704
rect 3699 5664 3792 5692
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4448 5692 4476 5732
rect 4724 5704 4752 5732
rect 4614 5692 4620 5704
rect 4111 5664 4476 5692
rect 4575 5664 4620 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4706 5652 4712 5704
rect 4764 5692 4770 5704
rect 5537 5695 5595 5701
rect 4764 5664 4857 5692
rect 4764 5652 4770 5664
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5644 5692 5672 5732
rect 5997 5729 6009 5763
rect 6043 5760 6055 5763
rect 6362 5760 6368 5772
rect 6043 5732 6368 5760
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 6362 5720 6368 5732
rect 6420 5720 6426 5772
rect 7024 5769 7052 5868
rect 7374 5856 7380 5868
rect 7432 5896 7438 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7432 5868 7849 5896
rect 7432 5856 7438 5868
rect 7837 5865 7849 5868
rect 7883 5896 7895 5899
rect 8570 5896 8576 5908
rect 7883 5868 8576 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 11057 5899 11115 5905
rect 11057 5865 11069 5899
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 11072 5828 11100 5859
rect 11514 5856 11520 5908
rect 11572 5896 11578 5908
rect 11793 5899 11851 5905
rect 11793 5896 11805 5899
rect 11572 5868 11805 5896
rect 11572 5856 11578 5868
rect 11793 5865 11805 5868
rect 11839 5865 11851 5899
rect 12434 5896 12440 5908
rect 11793 5859 11851 5865
rect 12084 5868 12440 5896
rect 7392 5800 11100 5828
rect 11701 5831 11759 5837
rect 7392 5772 7420 5800
rect 11701 5797 11713 5831
rect 11747 5828 11759 5831
rect 12084 5828 12112 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 14185 5899 14243 5905
rect 14185 5896 14197 5899
rect 14056 5868 14197 5896
rect 14056 5856 14062 5868
rect 14185 5865 14197 5868
rect 14231 5865 14243 5899
rect 14185 5859 14243 5865
rect 14200 5828 14228 5859
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 15654 5896 15660 5908
rect 15252 5868 15660 5896
rect 15252 5856 15258 5868
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 15838 5896 15844 5908
rect 15799 5868 15844 5896
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 16209 5899 16267 5905
rect 16209 5865 16221 5899
rect 16255 5896 16267 5899
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 16255 5868 16681 5896
rect 16255 5865 16267 5868
rect 16209 5859 16267 5865
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 17494 5896 17500 5908
rect 16669 5859 16727 5865
rect 16960 5868 17264 5896
rect 17455 5868 17500 5896
rect 16960 5828 16988 5868
rect 11747 5800 12112 5828
rect 12176 5800 14136 5828
rect 14200 5800 16988 5828
rect 11747 5797 11759 5800
rect 11701 5791 11759 5797
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5729 7067 5763
rect 7374 5760 7380 5772
rect 7287 5732 7380 5760
rect 7009 5723 7067 5729
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 9944 5763 10002 5769
rect 9732 5732 9777 5760
rect 9732 5720 9738 5732
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 10318 5760 10324 5772
rect 9990 5732 10324 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 12176 5760 12204 5800
rect 10704 5732 12204 5760
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 5644 5664 6837 5692
rect 5537 5655 5595 5661
rect 6825 5661 6837 5664
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5692 7803 5695
rect 8478 5692 8484 5704
rect 7791 5664 8484 5692
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 2869 5627 2927 5633
rect 2869 5593 2881 5627
rect 2915 5624 2927 5627
rect 3804 5624 3832 5652
rect 5552 5624 5580 5655
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 2915 5596 3740 5624
rect 3804 5596 5580 5624
rect 2915 5593 2927 5596
rect 2869 5587 2927 5593
rect 1854 5556 1860 5568
rect 1815 5528 1860 5556
rect 1854 5516 1860 5528
rect 1912 5516 1918 5568
rect 2222 5556 2228 5568
rect 2183 5528 2228 5556
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 3142 5556 3148 5568
rect 3103 5528 3148 5556
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 3712 5556 3740 5596
rect 5810 5556 5816 5568
rect 3712 5528 5816 5556
rect 5810 5516 5816 5528
rect 5868 5516 5874 5568
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 10704 5556 10732 5732
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 13061 5763 13119 5769
rect 13061 5760 13073 5763
rect 12400 5732 13073 5760
rect 12400 5720 12406 5732
rect 13061 5729 13073 5732
rect 13107 5729 13119 5763
rect 14108 5760 14136 5800
rect 15746 5760 15752 5772
rect 14108 5732 15752 5760
rect 13061 5723 13119 5729
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5760 16359 5763
rect 16666 5760 16672 5772
rect 16347 5732 16672 5760
rect 16347 5729 16359 5732
rect 16301 5723 16359 5729
rect 16666 5720 16672 5732
rect 16724 5720 16730 5772
rect 17037 5763 17095 5769
rect 17037 5760 17049 5763
rect 16776 5732 17049 5760
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5661 11943 5695
rect 11885 5655 11943 5661
rect 11900 5624 11928 5655
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12805 5695 12863 5701
rect 12805 5692 12817 5695
rect 12032 5664 12817 5692
rect 12032 5652 12038 5664
rect 12805 5661 12817 5664
rect 12851 5661 12863 5695
rect 16482 5692 16488 5704
rect 16443 5664 16488 5692
rect 12805 5655 12863 5661
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 12342 5624 12348 5636
rect 11900 5596 12348 5624
rect 12342 5584 12348 5596
rect 12400 5584 12406 5636
rect 16206 5584 16212 5636
rect 16264 5624 16270 5636
rect 16776 5624 16804 5732
rect 17037 5729 17049 5732
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 17236 5704 17264 5868
rect 17494 5856 17500 5868
rect 17552 5856 17558 5908
rect 17678 5760 17684 5772
rect 17639 5732 17684 5760
rect 17678 5720 17684 5732
rect 17736 5760 17742 5772
rect 17865 5763 17923 5769
rect 17865 5760 17877 5763
rect 17736 5732 17877 5760
rect 17736 5720 17742 5732
rect 17865 5729 17877 5732
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 17126 5692 17132 5704
rect 17087 5664 17132 5692
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 17218 5652 17224 5704
rect 17276 5692 17282 5704
rect 17276 5664 17369 5692
rect 17276 5652 17282 5664
rect 18046 5624 18052 5636
rect 16264 5596 16804 5624
rect 18007 5596 18052 5624
rect 16264 5584 16270 5596
rect 18046 5584 18052 5596
rect 18104 5584 18110 5636
rect 18138 5584 18144 5636
rect 18196 5624 18202 5636
rect 18196 5596 18460 5624
rect 18196 5584 18202 5596
rect 18432 5568 18460 5596
rect 11330 5556 11336 5568
rect 6871 5528 10732 5556
rect 11291 5528 11336 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 17954 5556 17960 5568
rect 13872 5528 17960 5556
rect 13872 5516 13878 5528
rect 17954 5516 17960 5528
rect 18012 5556 18018 5568
rect 18233 5559 18291 5565
rect 18233 5556 18245 5559
rect 18012 5528 18245 5556
rect 18012 5516 18018 5528
rect 18233 5525 18245 5528
rect 18279 5525 18291 5559
rect 18414 5556 18420 5568
rect 18375 5528 18420 5556
rect 18233 5519 18291 5525
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 3602 5312 3608 5364
rect 3660 5352 3666 5364
rect 4065 5355 4123 5361
rect 4065 5352 4077 5355
rect 3660 5324 4077 5352
rect 3660 5312 3666 5324
rect 4065 5321 4077 5324
rect 4111 5321 4123 5355
rect 4065 5315 4123 5321
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 11330 5352 11336 5364
rect 4396 5324 11336 5352
rect 4396 5312 4402 5324
rect 11330 5312 11336 5324
rect 11388 5312 11394 5364
rect 16206 5352 16212 5364
rect 16167 5324 16212 5352
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 16666 5352 16672 5364
rect 16627 5324 16672 5352
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 2590 5284 2596 5296
rect 2551 5256 2596 5284
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 6454 5244 6460 5296
rect 6512 5284 6518 5296
rect 6641 5287 6699 5293
rect 6641 5284 6653 5287
rect 6512 5256 6653 5284
rect 6512 5244 6518 5256
rect 6641 5253 6653 5256
rect 6687 5253 6699 5287
rect 12437 5287 12495 5293
rect 12437 5284 12449 5287
rect 6641 5247 6699 5253
rect 11256 5256 12449 5284
rect 2608 5216 2636 5244
rect 11256 5228 11284 5256
rect 12437 5253 12449 5256
rect 12483 5253 12495 5287
rect 12437 5247 12495 5253
rect 16114 5244 16120 5296
rect 16172 5284 16178 5296
rect 18417 5287 18475 5293
rect 18417 5284 18429 5287
rect 16172 5256 18429 5284
rect 16172 5244 16178 5256
rect 2148 5188 2636 5216
rect 2148 5157 2176 5188
rect 3142 5176 3148 5228
rect 3200 5216 3206 5228
rect 3697 5219 3755 5225
rect 3697 5216 3709 5219
rect 3200 5188 3709 5216
rect 3200 5176 3206 5188
rect 3697 5185 3709 5188
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5216 3939 5219
rect 4522 5216 4528 5228
rect 3927 5188 4528 5216
rect 3927 5185 3939 5188
rect 3881 5179 3939 5185
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 4706 5216 4712 5228
rect 4667 5188 4712 5216
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 5258 5216 5264 5228
rect 5219 5188 5264 5216
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 11238 5216 11244 5228
rect 11199 5188 11244 5216
rect 11238 5176 11244 5188
rect 11296 5176 11302 5228
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 14274 5216 14280 5228
rect 12299 5188 14136 5216
rect 14235 5188 14280 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5148 1639 5151
rect 2133 5151 2191 5157
rect 1627 5120 2084 5148
rect 1627 5117 1639 5120
rect 1581 5111 1639 5117
rect 1394 5040 1400 5092
rect 1452 5080 1458 5092
rect 1857 5083 1915 5089
rect 1857 5080 1869 5083
rect 1452 5052 1869 5080
rect 1452 5040 1458 5052
rect 1857 5049 1869 5052
rect 1903 5049 1915 5083
rect 2056 5080 2084 5120
rect 2133 5117 2145 5151
rect 2179 5117 2191 5151
rect 2133 5111 2191 5117
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5148 2743 5151
rect 3605 5151 3663 5157
rect 2731 5120 3556 5148
rect 2731 5117 2743 5120
rect 2685 5111 2743 5117
rect 2056 5052 2452 5080
rect 1857 5043 1915 5049
rect 2314 5012 2320 5024
rect 2275 4984 2320 5012
rect 2314 4972 2320 4984
rect 2372 4972 2378 5024
rect 2424 5012 2452 5052
rect 2774 5040 2780 5092
rect 2832 5080 2838 5092
rect 2961 5083 3019 5089
rect 2961 5080 2973 5083
rect 2832 5052 2973 5080
rect 2832 5040 2838 5052
rect 2961 5049 2973 5052
rect 3007 5049 3019 5083
rect 3528 5080 3556 5120
rect 3605 5117 3617 5151
rect 3651 5148 3663 5151
rect 5074 5148 5080 5160
rect 3651 5120 5080 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5276 5148 5304 5176
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 5276 5120 6837 5148
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 7092 5151 7150 5157
rect 7092 5117 7104 5151
rect 7138 5148 7150 5151
rect 7374 5148 7380 5160
rect 7138 5120 7380 5148
rect 7138 5117 7150 5120
rect 7092 5111 7150 5117
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5117 9275 5151
rect 14108 5148 14136 5188
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 15562 5176 15568 5228
rect 15620 5216 15626 5228
rect 16301 5219 16359 5225
rect 16301 5216 16313 5219
rect 15620 5188 16313 5216
rect 15620 5176 15626 5188
rect 16301 5185 16313 5188
rect 16347 5216 16359 5219
rect 16482 5216 16488 5228
rect 16347 5188 16488 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 16577 5219 16635 5225
rect 16577 5185 16589 5219
rect 16623 5216 16635 5219
rect 16942 5216 16948 5228
rect 16623 5188 16948 5216
rect 16623 5185 16635 5188
rect 16577 5179 16635 5185
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 17218 5216 17224 5228
rect 17179 5188 17224 5216
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 17770 5176 17776 5228
rect 17828 5176 17834 5228
rect 17402 5148 17408 5160
rect 14108 5120 17408 5148
rect 9217 5111 9275 5117
rect 4338 5080 4344 5092
rect 3528 5052 4344 5080
rect 2961 5043 3019 5049
rect 4338 5040 4344 5052
rect 4396 5040 4402 5092
rect 4433 5083 4491 5089
rect 4433 5049 4445 5083
rect 4479 5080 4491 5083
rect 5350 5080 5356 5092
rect 4479 5052 5356 5080
rect 4479 5049 4491 5052
rect 4433 5043 4491 5049
rect 5350 5040 5356 5052
rect 5408 5040 5414 5092
rect 5442 5040 5448 5092
rect 5500 5089 5506 5092
rect 5500 5083 5564 5089
rect 5500 5049 5518 5083
rect 5552 5049 5564 5083
rect 5500 5043 5564 5049
rect 5500 5040 5506 5043
rect 3237 5015 3295 5021
rect 3237 5012 3249 5015
rect 2424 4984 3249 5012
rect 3237 4981 3249 4984
rect 3283 4981 3295 5015
rect 3237 4975 3295 4981
rect 4522 4972 4528 5024
rect 4580 5012 4586 5024
rect 4580 4984 4625 5012
rect 4580 4972 4586 4984
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 7524 4984 8217 5012
rect 7524 4972 7530 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 9232 5012 9260 5111
rect 17402 5108 17408 5120
rect 17460 5108 17466 5160
rect 17494 5108 17500 5160
rect 17552 5148 17558 5160
rect 17589 5151 17647 5157
rect 17589 5148 17601 5151
rect 17552 5120 17601 5148
rect 17552 5108 17558 5120
rect 17589 5117 17601 5120
rect 17635 5117 17647 5151
rect 17589 5111 17647 5117
rect 9484 5083 9542 5089
rect 9484 5049 9496 5083
rect 9530 5080 9542 5083
rect 9766 5080 9772 5092
rect 9530 5052 9772 5080
rect 9530 5049 9542 5052
rect 9484 5043 9542 5049
rect 9766 5040 9772 5052
rect 9824 5040 9830 5092
rect 10962 5040 10968 5092
rect 11020 5080 11026 5092
rect 11333 5083 11391 5089
rect 11333 5080 11345 5083
rect 11020 5052 11345 5080
rect 11020 5040 11026 5052
rect 11333 5049 11345 5052
rect 11379 5080 11391 5083
rect 13265 5083 13323 5089
rect 11379 5052 13216 5080
rect 11379 5049 11391 5052
rect 11333 5043 11391 5049
rect 13188 5024 13216 5052
rect 13265 5049 13277 5083
rect 13311 5049 13323 5083
rect 13265 5043 13323 5049
rect 9674 5012 9680 5024
rect 9232 4984 9680 5012
rect 8205 4975 8263 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 10594 5012 10600 5024
rect 10555 4984 10600 5012
rect 10594 4972 10600 4984
rect 10652 4972 10658 5024
rect 13170 4972 13176 5024
rect 13228 4972 13234 5024
rect 13280 5012 13308 5043
rect 13354 5040 13360 5092
rect 13412 5080 13418 5092
rect 17037 5083 17095 5089
rect 13412 5052 13457 5080
rect 13412 5040 13418 5052
rect 17037 5049 17049 5083
rect 17083 5080 17095 5083
rect 17788 5080 17816 5176
rect 18064 5157 18092 5256
rect 18417 5253 18429 5256
rect 18463 5253 18475 5287
rect 18417 5247 18475 5253
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 17083 5052 17816 5080
rect 17083 5049 17095 5052
rect 17037 5043 17095 5049
rect 13538 5012 13544 5024
rect 13280 4984 13544 5012
rect 13538 4972 13544 4984
rect 13596 5012 13602 5024
rect 14369 5015 14427 5021
rect 14369 5012 14381 5015
rect 13596 4984 14381 5012
rect 13596 4972 13602 4984
rect 14369 4981 14381 4984
rect 14415 4981 14427 5015
rect 14369 4975 14427 4981
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17129 5015 17187 5021
rect 17129 5012 17141 5015
rect 17000 4984 17141 5012
rect 17000 4972 17006 4984
rect 17129 4981 17141 4984
rect 17175 5012 17187 5015
rect 17494 5012 17500 5024
rect 17175 4984 17500 5012
rect 17175 4981 17187 4984
rect 17129 4975 17187 4981
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 2222 4808 2228 4820
rect 2183 4780 2228 4808
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 4522 4808 4528 4820
rect 4483 4780 4528 4808
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4808 4951 4811
rect 5166 4808 5172 4820
rect 4939 4780 5172 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 5350 4808 5356 4820
rect 5311 4780 5356 4808
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4808 5871 4811
rect 6086 4808 6092 4820
rect 5859 4780 6092 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 6086 4768 6092 4780
rect 6144 4808 6150 4820
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 6144 4780 6193 4808
rect 6144 4768 6150 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 6181 4771 6239 4777
rect 9769 4811 9827 4817
rect 9769 4777 9781 4811
rect 9815 4808 9827 4811
rect 10318 4808 10324 4820
rect 9815 4780 10324 4808
rect 9815 4777 9827 4780
rect 9769 4771 9827 4777
rect 10318 4768 10324 4780
rect 10376 4808 10382 4820
rect 10686 4808 10692 4820
rect 10376 4780 10692 4808
rect 10376 4768 10382 4780
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 12066 4808 12072 4820
rect 12027 4780 12072 4808
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12158 4768 12164 4820
rect 12216 4808 12222 4820
rect 12216 4780 12388 4808
rect 12216 4768 12222 4780
rect 10496 4743 10554 4749
rect 4264 4712 8524 4740
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4672 1731 4675
rect 1719 4644 2176 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 1854 4468 1860 4480
rect 1815 4440 1860 4468
rect 1854 4428 1860 4440
rect 1912 4428 1918 4480
rect 2148 4477 2176 4644
rect 2133 4471 2191 4477
rect 2133 4437 2145 4471
rect 2179 4468 2191 4471
rect 4264 4468 4292 4712
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 4798 4672 4804 4684
rect 4479 4644 4804 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 4798 4632 4804 4644
rect 4856 4672 4862 4684
rect 8294 4681 8300 4684
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4856 4644 4997 4672
rect 4856 4632 4862 4644
rect 4985 4641 4997 4644
rect 5031 4641 5043 4675
rect 5721 4675 5779 4681
rect 5721 4672 5733 4675
rect 4985 4635 5043 4641
rect 5092 4644 5733 4672
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 5092 4604 5120 4644
rect 5721 4641 5733 4644
rect 5767 4672 5779 4675
rect 6549 4675 6607 4681
rect 6549 4672 6561 4675
rect 5767 4644 6561 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 6549 4641 6561 4644
rect 6595 4641 6607 4675
rect 6549 4635 6607 4641
rect 8288 4635 8300 4681
rect 8352 4672 8358 4684
rect 8496 4672 8524 4712
rect 10496 4709 10508 4743
rect 10542 4740 10554 4743
rect 10594 4740 10600 4752
rect 10542 4712 10600 4740
rect 10542 4709 10554 4712
rect 10496 4703 10554 4709
rect 10594 4700 10600 4712
rect 10652 4700 10658 4752
rect 12084 4740 12112 4768
rect 12360 4749 12388 4780
rect 13354 4768 13360 4820
rect 13412 4808 13418 4820
rect 13495 4811 13553 4817
rect 13495 4808 13507 4811
rect 13412 4780 13507 4808
rect 13412 4768 13418 4780
rect 13495 4777 13507 4780
rect 13541 4777 13553 4811
rect 16574 4808 16580 4820
rect 16535 4780 16580 4808
rect 13495 4771 13553 4777
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 16942 4808 16948 4820
rect 16903 4780 16948 4808
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 12253 4743 12311 4749
rect 12253 4740 12265 4743
rect 12084 4712 12265 4740
rect 12253 4709 12265 4712
rect 12299 4709 12311 4743
rect 12253 4703 12311 4709
rect 12354 4743 12412 4749
rect 12354 4709 12366 4743
rect 12400 4709 12412 4743
rect 15470 4740 15476 4752
rect 15431 4712 15476 4740
rect 12354 4703 12412 4709
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 16390 4740 16396 4752
rect 16351 4712 16396 4740
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 16482 4700 16488 4752
rect 16540 4740 16546 4752
rect 16850 4740 16856 4752
rect 16540 4712 16856 4740
rect 16540 4700 16546 4712
rect 16850 4700 16856 4712
rect 16908 4740 16914 4752
rect 17037 4743 17095 4749
rect 17037 4740 17049 4743
rect 16908 4712 17049 4740
rect 16908 4700 16914 4712
rect 17037 4709 17049 4712
rect 17083 4709 17095 4743
rect 17037 4703 17095 4709
rect 8352 4644 8388 4672
rect 8496 4644 11284 4672
rect 8294 4632 8300 4635
rect 8352 4632 8358 4644
rect 4948 4576 5120 4604
rect 5169 4607 5227 4613
rect 4948 4564 4954 4576
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5350 4604 5356 4616
rect 5215 4576 5356 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 5350 4564 5356 4576
rect 5408 4604 5414 4616
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5408 4576 6009 4604
rect 5408 4564 5414 4576
rect 5997 4573 6009 4576
rect 6043 4604 6055 4607
rect 6086 4604 6092 4616
rect 6043 4576 6092 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7156 4576 8033 4604
rect 7156 4564 7162 4576
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 8021 4567 8079 4573
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9732 4576 10241 4604
rect 9732 4564 9738 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 4522 4496 4528 4548
rect 4580 4536 4586 4548
rect 7926 4536 7932 4548
rect 4580 4508 7932 4536
rect 4580 4496 4586 4508
rect 7926 4496 7932 4508
rect 7984 4496 7990 4548
rect 9401 4539 9459 4545
rect 9401 4505 9413 4539
rect 9447 4536 9459 4539
rect 9766 4536 9772 4548
rect 9447 4508 9772 4536
rect 9447 4505 9459 4508
rect 9401 4499 9459 4505
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 11256 4536 11284 4644
rect 13170 4632 13176 4684
rect 13228 4672 13234 4684
rect 13392 4675 13450 4681
rect 13392 4672 13404 4675
rect 13228 4644 13404 4672
rect 13228 4632 13234 4644
rect 13392 4641 13404 4644
rect 13438 4641 13450 4675
rect 13392 4635 13450 4641
rect 13998 4632 14004 4684
rect 14056 4672 14062 4684
rect 14220 4675 14278 4681
rect 14220 4672 14232 4675
rect 14056 4644 14232 4672
rect 14056 4632 14062 4644
rect 14220 4641 14232 4644
rect 14266 4641 14278 4675
rect 17402 4672 17408 4684
rect 17363 4644 17408 4672
rect 14220 4635 14278 4641
rect 17402 4632 17408 4644
rect 17460 4632 17466 4684
rect 17865 4675 17923 4681
rect 17865 4641 17877 4675
rect 17911 4672 17923 4675
rect 17954 4672 17960 4684
rect 17911 4644 17960 4672
rect 17911 4641 17923 4644
rect 17865 4635 17923 4641
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4672 18291 4675
rect 18414 4672 18420 4684
rect 18279 4644 18420 4672
rect 18279 4641 18291 4644
rect 18233 4635 18291 4641
rect 18414 4632 18420 4644
rect 18472 4632 18478 4684
rect 13265 4607 13323 4613
rect 13265 4573 13277 4607
rect 13311 4604 13323 4607
rect 14918 4604 14924 4616
rect 13311 4576 14924 4604
rect 13311 4573 13323 4576
rect 13265 4567 13323 4573
rect 14918 4564 14924 4576
rect 14976 4564 14982 4616
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 15028 4576 15393 4604
rect 12618 4536 12624 4548
rect 11256 4508 12624 4536
rect 12618 4496 12624 4508
rect 12676 4496 12682 4548
rect 2179 4440 4292 4468
rect 2179 4437 2191 4440
rect 2133 4431 2191 4437
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 6365 4471 6423 4477
rect 6365 4468 6377 4471
rect 5224 4440 6377 4468
rect 5224 4428 5230 4440
rect 6365 4437 6377 4440
rect 6411 4437 6423 4471
rect 11606 4468 11612 4480
rect 11567 4440 11612 4468
rect 6365 4431 6423 4437
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 14274 4428 14280 4480
rect 14332 4477 14338 4480
rect 14332 4471 14381 4477
rect 14332 4437 14335 4471
rect 14369 4437 14381 4471
rect 14332 4431 14381 4437
rect 14332 4428 14338 4431
rect 14642 4428 14648 4480
rect 14700 4468 14706 4480
rect 15028 4477 15056 4576
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 17218 4604 17224 4616
rect 17179 4576 17224 4604
rect 15381 4567 15439 4573
rect 17218 4564 17224 4576
rect 17276 4564 17282 4616
rect 17589 4539 17647 4545
rect 17589 4505 17601 4539
rect 17635 4536 17647 4539
rect 18138 4536 18144 4548
rect 17635 4508 18144 4536
rect 17635 4505 17647 4508
rect 17589 4499 17647 4505
rect 18138 4496 18144 4508
rect 18196 4496 18202 4548
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 14700 4440 15025 4468
rect 14700 4428 14706 4440
rect 15013 4437 15025 4440
rect 15059 4437 15071 4471
rect 15013 4431 15071 4437
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 18049 4471 18107 4477
rect 18049 4468 18061 4471
rect 17920 4440 18061 4468
rect 17920 4428 17926 4440
rect 18049 4437 18061 4440
rect 18095 4437 18107 4471
rect 18414 4468 18420 4480
rect 18375 4440 18420 4468
rect 18049 4431 18107 4437
rect 18414 4428 18420 4440
rect 18472 4428 18478 4480
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 5166 4264 5172 4276
rect 3988 4236 5172 4264
rect 2222 4196 2228 4208
rect 1596 4168 2228 4196
rect 1596 4069 1624 4168
rect 2222 4156 2228 4168
rect 2280 4156 2286 4208
rect 2685 4199 2743 4205
rect 2685 4165 2697 4199
rect 2731 4196 2743 4199
rect 2731 4168 3188 4196
rect 2731 4165 2743 4168
rect 2685 4159 2743 4165
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 3050 4128 3056 4140
rect 1903 4100 3056 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 3160 4128 3188 4168
rect 3234 4128 3240 4140
rect 3160 4100 3240 4128
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3988 4128 4016 4236
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 5350 4264 5356 4276
rect 5311 4236 5356 4264
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 5920 4236 6469 4264
rect 3896 4100 4016 4128
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4029 1639 4063
rect 1581 4023 1639 4029
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4029 2191 4063
rect 2133 4023 2191 4029
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 2961 4063 3019 4069
rect 2961 4060 2973 4063
rect 2547 4032 2973 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 2961 4029 2973 4032
rect 3007 4060 3019 4063
rect 3896 4060 3924 4100
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 5920 4137 5948 4236
rect 6457 4233 6469 4236
rect 6503 4233 6515 4267
rect 6457 4227 6515 4233
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 8352 4236 8493 4264
rect 8352 4224 8358 4236
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 8481 4227 8539 4233
rect 11256 4236 11468 4264
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5776 4100 5917 4128
rect 5776 4088 5782 4100
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 6086 4128 6092 4140
rect 6047 4100 6092 4128
rect 5905 4091 5963 4097
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 8496 4128 8524 4227
rect 8570 4156 8576 4208
rect 8628 4196 8634 4208
rect 9401 4199 9459 4205
rect 9401 4196 9413 4199
rect 8628 4168 9413 4196
rect 8628 4156 8634 4168
rect 9401 4165 9413 4168
rect 9447 4165 9459 4199
rect 10778 4196 10784 4208
rect 9401 4159 9459 4165
rect 9784 4168 10784 4196
rect 9784 4128 9812 4168
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 8496 4100 8984 4128
rect 3007 4032 3924 4060
rect 3973 4063 4031 4069
rect 3007 4029 3019 4032
rect 2961 4023 3019 4029
rect 3973 4029 3985 4063
rect 4019 4060 4031 4063
rect 5258 4060 5264 4072
rect 4019 4032 5264 4060
rect 4019 4029 4031 4032
rect 3973 4023 4031 4029
rect 2148 3992 2176 4023
rect 5258 4020 5264 4032
rect 5316 4060 5322 4072
rect 6638 4060 6644 4072
rect 5316 4032 6644 4060
rect 5316 4020 5322 4032
rect 6638 4020 6644 4032
rect 6696 4060 6702 4072
rect 7098 4060 7104 4072
rect 6696 4032 7104 4060
rect 6696 4020 6702 4032
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 8956 4069 8984 4100
rect 9048 4100 9812 4128
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 3053 3995 3111 4001
rect 3053 3992 3065 3995
rect 2148 3964 3065 3992
rect 3053 3961 3065 3964
rect 3099 3961 3111 3995
rect 3053 3955 3111 3961
rect 4240 3995 4298 4001
rect 4240 3961 4252 3995
rect 4286 3992 4298 3995
rect 4430 3992 4436 4004
rect 4286 3964 4436 3992
rect 4286 3961 4298 3964
rect 4240 3955 4298 3961
rect 2314 3924 2320 3936
rect 2275 3896 2320 3924
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 3068 3924 3096 3955
rect 4430 3952 4436 3964
rect 4488 3992 4494 4004
rect 6273 3995 6331 4001
rect 6273 3992 6285 3995
rect 4488 3964 6285 3992
rect 4488 3952 4494 3964
rect 6273 3961 6285 3964
rect 6319 3961 6331 3995
rect 6273 3955 6331 3961
rect 7368 3995 7426 4001
rect 7368 3961 7380 3995
rect 7414 3992 7426 3995
rect 8018 3992 8024 4004
rect 7414 3964 8024 3992
rect 7414 3961 7426 3964
rect 7368 3955 7426 3961
rect 8018 3952 8024 3964
rect 8076 3952 8082 4004
rect 4522 3924 4528 3936
rect 3068 3896 4528 3924
rect 4522 3884 4528 3896
rect 4580 3884 4586 3936
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 5445 3927 5503 3933
rect 5445 3924 5457 3927
rect 4672 3896 5457 3924
rect 4672 3884 4678 3896
rect 5445 3893 5457 3896
rect 5491 3893 5503 3927
rect 5810 3924 5816 3936
rect 5723 3896 5816 3924
rect 5445 3887 5503 3893
rect 5810 3884 5816 3896
rect 5868 3924 5874 3936
rect 6917 3927 6975 3933
rect 6917 3924 6929 3927
rect 5868 3896 6929 3924
rect 5868 3884 5874 3896
rect 6917 3893 6929 3896
rect 6963 3924 6975 3927
rect 9048 3924 9076 4100
rect 9858 4088 9864 4140
rect 9916 4128 9922 4140
rect 10965 4131 11023 4137
rect 10965 4128 10977 4131
rect 9916 4100 10977 4128
rect 9916 4088 9922 4100
rect 10965 4097 10977 4100
rect 11011 4128 11023 4131
rect 11256 4128 11284 4236
rect 11011 4100 11284 4128
rect 11440 4128 11468 4236
rect 14366 4224 14372 4276
rect 14424 4224 14430 4276
rect 11514 4156 11520 4208
rect 11572 4196 11578 4208
rect 11977 4199 12035 4205
rect 11977 4196 11989 4199
rect 11572 4168 11989 4196
rect 11572 4156 11578 4168
rect 11977 4165 11989 4168
rect 12023 4165 12035 4199
rect 13998 4196 14004 4208
rect 11977 4159 12035 4165
rect 12820 4168 14004 4196
rect 12820 4128 12848 4168
rect 13998 4156 14004 4168
rect 14056 4156 14062 4208
rect 14384 4196 14412 4224
rect 14384 4168 14964 4196
rect 11440 4100 12848 4128
rect 12897 4131 12955 4137
rect 11011 4097 11023 4100
rect 10965 4091 11023 4097
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13078 4128 13084 4140
rect 12943 4100 13084 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13354 4128 13360 4140
rect 13315 4100 13360 4128
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 14185 4131 14243 4137
rect 14185 4097 14197 4131
rect 14231 4128 14243 4131
rect 14366 4128 14372 4140
rect 14231 4100 14372 4128
rect 14231 4097 14243 4100
rect 14185 4091 14243 4097
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 14826 4128 14832 4140
rect 14787 4100 14832 4128
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 14936 4128 14964 4168
rect 16298 4128 16304 4140
rect 14936 4100 16304 4128
rect 16298 4088 16304 4100
rect 16356 4128 16362 4140
rect 16577 4131 16635 4137
rect 16577 4128 16589 4131
rect 16356 4100 16589 4128
rect 16356 4088 16362 4100
rect 16577 4097 16589 4100
rect 16623 4097 16635 4131
rect 17218 4128 17224 4140
rect 17179 4100 17224 4128
rect 16577 4091 16635 4097
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 9766 4060 9772 4072
rect 9727 4032 9772 4060
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 10321 4063 10379 4069
rect 10321 4060 10333 4063
rect 10192 4032 10333 4060
rect 10192 4020 10198 4032
rect 10321 4029 10333 4032
rect 10367 4060 10379 4063
rect 10502 4060 10508 4072
rect 10367 4032 10508 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 10689 4063 10747 4069
rect 10689 4060 10701 4063
rect 10652 4032 10701 4060
rect 10652 4020 10658 4032
rect 10689 4029 10701 4032
rect 10735 4029 10747 4063
rect 10689 4023 10747 4029
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 11149 4063 11207 4069
rect 11149 4060 11161 4063
rect 10836 4032 11161 4060
rect 10836 4020 10842 4032
rect 11149 4029 11161 4032
rect 11195 4060 11207 4063
rect 11422 4060 11428 4072
rect 11195 4032 11428 4060
rect 11195 4029 11207 4032
rect 11149 4023 11207 4029
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 11517 4063 11575 4069
rect 11517 4029 11529 4063
rect 11563 4060 11575 4063
rect 11606 4060 11612 4072
rect 11563 4032 11612 4060
rect 11563 4029 11575 4032
rect 11517 4023 11575 4029
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 12158 4060 12164 4072
rect 11716 4032 12164 4060
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 9272 3964 9321 3992
rect 9272 3952 9278 3964
rect 9309 3961 9321 3964
rect 9355 3992 9367 3995
rect 11716 3992 11744 4032
rect 12158 4020 12164 4032
rect 12216 4060 12222 4072
rect 12564 4063 12622 4069
rect 12564 4060 12576 4063
rect 12216 4032 12576 4060
rect 12216 4020 12222 4032
rect 12564 4029 12576 4032
rect 12610 4029 12622 4063
rect 12564 4023 12622 4029
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17552 4032 18061 4060
rect 17552 4020 17558 4032
rect 18049 4029 18061 4032
rect 18095 4060 18107 4063
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 18095 4032 18429 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 11882 3992 11888 4004
rect 9355 3964 11744 3992
rect 11843 3964 11888 3992
rect 9355 3961 9367 3964
rect 9309 3955 9367 3961
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 12989 3995 13047 4001
rect 12989 3961 13001 3995
rect 13035 3961 13047 3995
rect 12989 3955 13047 3961
rect 6963 3896 9076 3924
rect 6963 3893 6975 3896
rect 6917 3887 6975 3893
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9824 3896 9873 3924
rect 9824 3884 9830 3896
rect 9861 3893 9873 3896
rect 9907 3924 9919 3927
rect 10962 3924 10968 3936
rect 9907 3896 10968 3924
rect 9907 3893 9919 3896
rect 9861 3887 9919 3893
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 11204 3896 12173 3924
rect 11204 3884 11210 3896
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 12161 3887 12219 3893
rect 12667 3927 12725 3933
rect 12667 3893 12679 3927
rect 12713 3924 12725 3927
rect 13004 3924 13032 3955
rect 14274 3952 14280 4004
rect 14332 3992 14338 4004
rect 14332 3964 14377 3992
rect 14332 3952 14338 3964
rect 14734 3952 14740 4004
rect 14792 3992 14798 4004
rect 15381 3995 15439 4001
rect 15381 3992 15393 3995
rect 14792 3964 15393 3992
rect 14792 3952 14798 3964
rect 15381 3961 15393 3964
rect 15427 3961 15439 3995
rect 15381 3955 15439 3961
rect 15473 3995 15531 4001
rect 15473 3961 15485 3995
rect 15519 3961 15531 3995
rect 16390 3992 16396 4004
rect 16351 3964 16396 3992
rect 15473 3955 15531 3961
rect 12713 3896 13032 3924
rect 12713 3893 12725 3896
rect 12667 3887 12725 3893
rect 13998 3884 14004 3936
rect 14056 3924 14062 3936
rect 15488 3924 15516 3955
rect 16390 3952 16396 3964
rect 16448 3952 16454 4004
rect 16669 3995 16727 4001
rect 16669 3961 16681 3995
rect 16715 3961 16727 3995
rect 18690 3992 18696 4004
rect 16669 3955 16727 3961
rect 17788 3964 18696 3992
rect 14056 3896 15516 3924
rect 14056 3884 14062 3896
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 16684 3924 16712 3955
rect 17788 3936 17816 3964
rect 18690 3952 18696 3964
rect 18748 3952 18754 4004
rect 17770 3924 17776 3936
rect 16172 3896 16712 3924
rect 17731 3896 17776 3924
rect 16172 3884 16178 3896
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18230 3924 18236 3936
rect 18191 3896 18236 3924
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 2133 3723 2191 3729
rect 2133 3720 2145 3723
rect 1728 3692 2145 3720
rect 1728 3680 1734 3692
rect 2133 3689 2145 3692
rect 2179 3720 2191 3723
rect 2406 3720 2412 3732
rect 2179 3692 2412 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 7282 3720 7288 3732
rect 3620 3692 7288 3720
rect 2317 3655 2375 3661
rect 2317 3652 2329 3655
rect 1688 3624 2329 3652
rect 1688 3593 1716 3624
rect 2317 3621 2329 3624
rect 2363 3652 2375 3655
rect 3620 3652 3648 3692
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 8018 3720 8024 3732
rect 7979 3692 8024 3720
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 8570 3720 8576 3732
rect 8168 3692 8576 3720
rect 8168 3680 8174 3692
rect 8570 3680 8576 3692
rect 8628 3720 8634 3732
rect 9309 3723 9367 3729
rect 9309 3720 9321 3723
rect 8628 3692 9321 3720
rect 8628 3680 8634 3692
rect 9309 3689 9321 3692
rect 9355 3720 9367 3723
rect 10134 3720 10140 3732
rect 9355 3692 10140 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 12069 3723 12127 3729
rect 12069 3720 12081 3723
rect 10284 3692 12081 3720
rect 10284 3680 10290 3692
rect 12069 3689 12081 3692
rect 12115 3689 12127 3723
rect 12069 3683 12127 3689
rect 12158 3680 12164 3732
rect 12216 3720 12222 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 12216 3692 12909 3720
rect 12216 3680 12222 3692
rect 12897 3689 12909 3692
rect 12943 3720 12955 3723
rect 13446 3720 13452 3732
rect 12943 3692 13452 3720
rect 12943 3689 12955 3692
rect 12897 3683 12955 3689
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 15841 3723 15899 3729
rect 15841 3720 15853 3723
rect 14424 3692 15853 3720
rect 14424 3680 14430 3692
rect 15841 3689 15853 3692
rect 15887 3689 15899 3723
rect 16850 3720 16856 3732
rect 16811 3692 16856 3720
rect 15841 3683 15899 3689
rect 16850 3680 16856 3692
rect 16908 3720 16914 3732
rect 17494 3720 17500 3732
rect 16908 3692 17500 3720
rect 16908 3680 16914 3692
rect 17494 3680 17500 3692
rect 17552 3680 17558 3732
rect 2363 3624 3648 3652
rect 5436 3655 5494 3661
rect 2363 3621 2375 3624
rect 2317 3615 2375 3621
rect 5436 3621 5448 3655
rect 5482 3652 5494 3655
rect 7466 3652 7472 3664
rect 5482 3624 7472 3652
rect 5482 3621 5494 3624
rect 5436 3615 5494 3621
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3553 1731 3587
rect 1673 3547 1731 3553
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3584 5227 3587
rect 5258 3584 5264 3596
rect 5215 3556 5264 3584
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 6908 3587 6966 3593
rect 6908 3584 6920 3587
rect 6472 3556 6920 3584
rect 1854 3448 1860 3460
rect 1815 3420 1860 3448
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 6472 3448 6500 3556
rect 6908 3553 6920 3556
rect 6954 3584 6966 3587
rect 7282 3584 7288 3596
rect 6954 3556 7288 3584
rect 6954 3553 6966 3556
rect 6908 3547 6966 3553
rect 7282 3544 7288 3556
rect 7340 3544 7346 3596
rect 8036 3584 8064 3680
rect 10410 3652 10416 3664
rect 8588 3624 10416 3652
rect 8481 3587 8539 3593
rect 8481 3584 8493 3587
rect 8036 3556 8493 3584
rect 8481 3553 8493 3556
rect 8527 3553 8539 3587
rect 8481 3547 8539 3553
rect 6638 3516 6644 3528
rect 6599 3488 6644 3516
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 8110 3516 8116 3528
rect 8071 3488 8116 3516
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 6549 3451 6607 3457
rect 6549 3448 6561 3451
rect 6472 3420 6561 3448
rect 6549 3417 6561 3420
rect 6595 3417 6607 3451
rect 6549 3411 6607 3417
rect 5166 3340 5172 3392
rect 5224 3380 5230 3392
rect 8588 3380 8616 3624
rect 10410 3612 10416 3624
rect 10468 3612 10474 3664
rect 10680 3655 10738 3661
rect 10680 3621 10692 3655
rect 10726 3652 10738 3655
rect 11606 3652 11612 3664
rect 10726 3624 11612 3652
rect 10726 3621 10738 3624
rect 10680 3615 10738 3621
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 16114 3652 16120 3664
rect 11900 3624 16120 3652
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3584 8999 3587
rect 9214 3584 9220 3596
rect 8987 3556 9220 3584
rect 8987 3553 8999 3556
rect 8941 3547 8999 3553
rect 9214 3544 9220 3556
rect 9272 3544 9278 3596
rect 9674 3544 9680 3596
rect 9732 3544 9738 3596
rect 9858 3584 9864 3596
rect 9819 3556 9864 3584
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 10134 3544 10140 3596
rect 10192 3584 10198 3596
rect 10229 3587 10287 3593
rect 10229 3584 10241 3587
rect 10192 3556 10241 3584
rect 10192 3544 10198 3556
rect 10229 3553 10241 3556
rect 10275 3553 10287 3587
rect 10428 3584 10456 3612
rect 11900 3596 11928 3624
rect 11882 3584 11888 3596
rect 10428 3556 11468 3584
rect 11843 3556 11888 3584
rect 10229 3547 10287 3553
rect 8846 3516 8852 3528
rect 8807 3488 8852 3516
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9692 3516 9720 3544
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 9692 3488 10425 3516
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 8754 3408 8760 3460
rect 8812 3448 8818 3460
rect 9677 3451 9735 3457
rect 9677 3448 9689 3451
rect 8812 3420 9689 3448
rect 8812 3408 8818 3420
rect 9677 3417 9689 3420
rect 9723 3448 9735 3451
rect 11440 3448 11468 3556
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 11974 3544 11980 3596
rect 12032 3584 12038 3596
rect 12288 3587 12346 3593
rect 12288 3584 12300 3587
rect 12032 3556 12300 3584
rect 12032 3544 12038 3556
rect 12288 3553 12300 3556
rect 12334 3553 12346 3587
rect 12288 3547 12346 3553
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 12596 3587 12654 3593
rect 12596 3584 12608 3587
rect 12492 3556 12608 3584
rect 12492 3544 12498 3556
rect 12596 3553 12608 3556
rect 12642 3584 12654 3587
rect 12986 3584 12992 3596
rect 12642 3556 12992 3584
rect 12642 3553 12654 3556
rect 12596 3547 12654 3553
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 13909 3587 13967 3593
rect 13909 3553 13921 3587
rect 13955 3584 13967 3587
rect 14090 3584 14096 3596
rect 13955 3556 14096 3584
rect 13955 3553 13967 3556
rect 13909 3547 13967 3553
rect 14090 3544 14096 3556
rect 14148 3544 14154 3596
rect 14550 3544 14556 3596
rect 14608 3544 14614 3596
rect 14734 3544 14740 3596
rect 14792 3584 14798 3596
rect 15013 3587 15071 3593
rect 15013 3584 15025 3587
rect 14792 3556 15025 3584
rect 14792 3544 14798 3556
rect 15013 3553 15025 3556
rect 15059 3553 15071 3587
rect 15212 3584 15240 3624
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 16390 3612 16396 3664
rect 16448 3652 16454 3664
rect 16448 3624 18276 3652
rect 16448 3612 16454 3624
rect 15470 3593 15476 3596
rect 15324 3587 15382 3593
rect 15324 3584 15336 3587
rect 15212 3556 15336 3584
rect 15013 3547 15071 3553
rect 15324 3553 15336 3556
rect 15370 3553 15382 3587
rect 15324 3547 15382 3553
rect 15427 3587 15476 3593
rect 15427 3553 15439 3587
rect 15473 3553 15476 3587
rect 15427 3547 15476 3553
rect 15470 3544 15476 3547
rect 15528 3544 15534 3596
rect 15632 3587 15690 3593
rect 15632 3553 15644 3587
rect 15678 3584 15690 3587
rect 16206 3584 16212 3596
rect 15678 3556 16212 3584
rect 15678 3553 15690 3556
rect 15632 3547 15690 3553
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 16298 3544 16304 3596
rect 16356 3584 16362 3596
rect 16669 3587 16727 3593
rect 16356 3556 16401 3584
rect 16356 3544 16362 3556
rect 16669 3553 16681 3587
rect 16715 3584 16727 3587
rect 16758 3584 16764 3596
rect 16715 3556 16764 3584
rect 16715 3553 16727 3556
rect 16669 3547 16727 3553
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 16945 3587 17003 3593
rect 16945 3553 16957 3587
rect 16991 3553 17003 3587
rect 16945 3547 17003 3553
rect 14568 3516 14596 3544
rect 14826 3516 14832 3528
rect 14568 3488 14832 3516
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 16960 3516 16988 3547
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 17276 3556 17325 3584
rect 17276 3544 17282 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17770 3544 17776 3596
rect 17828 3584 17834 3596
rect 18248 3593 18276 3624
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17828 3556 17877 3584
rect 17828 3544 17834 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3553 18291 3587
rect 18233 3547 18291 3553
rect 14976 3488 16988 3516
rect 14976 3476 14982 3488
rect 11793 3451 11851 3457
rect 11793 3448 11805 3451
rect 9723 3420 10364 3448
rect 11440 3420 11805 3448
rect 9723 3417 9735 3420
rect 9677 3411 9735 3417
rect 5224 3352 8616 3380
rect 5224 3340 5230 3352
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 9125 3383 9183 3389
rect 9125 3380 9137 3383
rect 8720 3352 9137 3380
rect 8720 3340 8726 3352
rect 9125 3349 9137 3352
rect 9171 3349 9183 3383
rect 9125 3343 9183 3349
rect 9766 3340 9772 3392
rect 9824 3380 9830 3392
rect 10045 3383 10103 3389
rect 10045 3380 10057 3383
rect 9824 3352 10057 3380
rect 9824 3340 9830 3352
rect 10045 3349 10057 3352
rect 10091 3349 10103 3383
rect 10336 3380 10364 3420
rect 11793 3417 11805 3420
rect 11839 3417 11851 3451
rect 11793 3411 11851 3417
rect 13170 3408 13176 3460
rect 13228 3448 13234 3460
rect 14001 3451 14059 3457
rect 14001 3448 14013 3451
rect 13228 3420 14013 3448
rect 13228 3408 13234 3420
rect 14001 3417 14013 3420
rect 14047 3417 14059 3451
rect 14001 3411 14059 3417
rect 15194 3408 15200 3460
rect 15252 3448 15258 3460
rect 16025 3451 16083 3457
rect 16025 3448 16037 3451
rect 15252 3420 16037 3448
rect 15252 3408 15258 3420
rect 16025 3417 16037 3420
rect 16071 3417 16083 3451
rect 16025 3411 16083 3417
rect 17497 3451 17555 3457
rect 17497 3417 17509 3451
rect 17543 3448 17555 3451
rect 19150 3448 19156 3460
rect 17543 3420 19156 3448
rect 17543 3417 17555 3420
rect 17497 3411 17555 3417
rect 19150 3408 19156 3420
rect 19208 3408 19214 3460
rect 11146 3380 11152 3392
rect 10336 3352 11152 3380
rect 10045 3343 10103 3349
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 11882 3340 11888 3392
rect 11940 3380 11946 3392
rect 12710 3389 12716 3392
rect 12391 3383 12449 3389
rect 12391 3380 12403 3383
rect 11940 3352 12403 3380
rect 11940 3340 11946 3352
rect 12391 3349 12403 3352
rect 12437 3349 12449 3383
rect 12391 3343 12449 3349
rect 12667 3383 12716 3389
rect 12667 3349 12679 3383
rect 12713 3349 12716 3383
rect 12667 3343 12716 3349
rect 12710 3340 12716 3343
rect 12768 3340 12774 3392
rect 13630 3380 13636 3392
rect 13591 3352 13636 3380
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 15654 3340 15660 3392
rect 15712 3389 15718 3392
rect 15712 3383 15761 3389
rect 15712 3349 15715 3383
rect 15749 3349 15761 3383
rect 15712 3343 15761 3349
rect 17129 3383 17187 3389
rect 17129 3349 17141 3383
rect 17175 3380 17187 3383
rect 17402 3380 17408 3392
rect 17175 3352 17408 3380
rect 17175 3349 17187 3352
rect 17129 3343 17187 3349
rect 15712 3340 15718 3343
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 17681 3383 17739 3389
rect 17681 3380 17693 3383
rect 17644 3352 17693 3380
rect 17644 3340 17650 3352
rect 17681 3349 17693 3352
rect 17727 3349 17739 3383
rect 18046 3380 18052 3392
rect 18007 3352 18052 3380
rect 17681 3343 17739 3349
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 18417 3383 18475 3389
rect 18417 3349 18429 3383
rect 18463 3380 18475 3383
rect 18598 3380 18604 3392
rect 18463 3352 18604 3380
rect 18463 3349 18475 3352
rect 18417 3343 18475 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 2958 3176 2964 3188
rect 2516 3148 2728 3176
rect 2919 3148 2964 3176
rect 2222 3108 2228 3120
rect 2183 3080 2228 3108
rect 2222 3068 2228 3080
rect 2280 3068 2286 3120
rect 1670 2972 1676 2984
rect 1631 2944 1676 2972
rect 1670 2932 1676 2944
rect 1728 2932 1734 2984
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2941 2099 2975
rect 2041 2935 2099 2941
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 2516 2972 2544 3148
rect 2593 3111 2651 3117
rect 2593 3077 2605 3111
rect 2639 3077 2651 3111
rect 2700 3108 2728 3148
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 7558 3176 7564 3188
rect 3200 3148 7564 3176
rect 3200 3136 3206 3148
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 8021 3179 8079 3185
rect 8021 3145 8033 3179
rect 8067 3176 8079 3179
rect 8110 3176 8116 3188
rect 8067 3148 8116 3176
rect 8067 3145 8079 3148
rect 8021 3139 8079 3145
rect 2869 3111 2927 3117
rect 2869 3108 2881 3111
rect 2700 3080 2881 3108
rect 2593 3071 2651 3077
rect 2869 3077 2881 3080
rect 2915 3108 2927 3111
rect 5810 3108 5816 3120
rect 2915 3080 5816 3108
rect 2915 3077 2927 3080
rect 2869 3071 2927 3077
rect 2455 2944 2544 2972
rect 2608 2972 2636 3071
rect 5810 3068 5816 3080
rect 5868 3068 5874 3120
rect 6730 3068 6736 3120
rect 6788 3108 6794 3120
rect 7009 3111 7067 3117
rect 7009 3108 7021 3111
rect 6788 3080 7021 3108
rect 6788 3068 6794 3080
rect 7009 3077 7021 3080
rect 7055 3108 7067 3111
rect 7101 3111 7159 3117
rect 7101 3108 7113 3111
rect 7055 3080 7113 3108
rect 7055 3077 7067 3080
rect 7009 3071 7067 3077
rect 7101 3077 7113 3080
rect 7147 3108 7159 3111
rect 8036 3108 8064 3139
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 12434 3176 12440 3188
rect 8444 3148 12440 3176
rect 8444 3136 8450 3148
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 12894 3136 12900 3188
rect 12952 3176 12958 3188
rect 12952 3148 17356 3176
rect 12952 3136 12958 3148
rect 8481 3111 8539 3117
rect 8481 3108 8493 3111
rect 7147 3080 8493 3108
rect 7147 3077 7159 3080
rect 7101 3071 7159 3077
rect 8481 3077 8493 3080
rect 8527 3077 8539 3111
rect 8481 3071 8539 3077
rect 8570 3068 8576 3120
rect 8628 3108 8634 3120
rect 8846 3108 8852 3120
rect 8628 3080 8852 3108
rect 8628 3068 8634 3080
rect 8846 3068 8852 3080
rect 8904 3108 8910 3120
rect 14274 3108 14280 3120
rect 8904 3080 14280 3108
rect 8904 3068 8910 3080
rect 14274 3068 14280 3080
rect 14332 3068 14338 3120
rect 14826 3068 14832 3120
rect 14884 3108 14890 3120
rect 15749 3111 15807 3117
rect 14884 3080 15675 3108
rect 14884 3068 14890 3080
rect 8754 3040 8760 3052
rect 8715 3012 8760 3040
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 9582 3040 9588 3052
rect 9543 3012 9588 3040
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 10594 3040 10600 3052
rect 9784 3012 10600 3040
rect 2866 2972 2872 2984
rect 2608 2944 2872 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 1394 2836 1400 2848
rect 256 2808 1400 2836
rect 256 2796 262 2808
rect 1394 2796 1400 2808
rect 1452 2796 1458 2848
rect 1854 2836 1860 2848
rect 1815 2808 1860 2836
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 2056 2836 2084 2935
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 7466 2972 7472 2984
rect 7427 2944 7472 2972
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 2222 2864 2228 2916
rect 2280 2904 2286 2916
rect 5534 2904 5540 2916
rect 2280 2876 5540 2904
rect 2280 2864 2286 2876
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 7837 2907 7895 2913
rect 7837 2873 7849 2907
rect 7883 2873 7895 2907
rect 7837 2867 7895 2873
rect 2958 2836 2964 2848
rect 2056 2808 2964 2836
rect 2958 2796 2964 2808
rect 3016 2796 3022 2848
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 7852 2836 7880 2867
rect 8846 2864 8852 2916
rect 8904 2904 8910 2916
rect 9784 2904 9812 3012
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11238 3040 11244 3052
rect 11195 3012 11244 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3040 12219 3043
rect 15647 3040 15675 3080
rect 15749 3077 15761 3111
rect 15795 3108 15807 3111
rect 16114 3108 16120 3120
rect 15795 3080 16120 3108
rect 15795 3077 15807 3080
rect 15749 3071 15807 3077
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 16025 3043 16083 3049
rect 16025 3040 16037 3043
rect 12207 3012 15608 3040
rect 15647 3012 16037 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 15580 2981 15608 3012
rect 16025 3009 16037 3012
rect 16071 3009 16083 3043
rect 17328 3040 17356 3148
rect 17405 3111 17463 3117
rect 17405 3077 17417 3111
rect 17451 3108 17463 3111
rect 19610 3108 19616 3120
rect 17451 3080 19616 3108
rect 17451 3077 17463 3080
rect 17405 3071 17463 3077
rect 19610 3068 19616 3080
rect 19668 3068 19674 3120
rect 17328 3012 18092 3040
rect 16025 3003 16083 3009
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12400 2944 12449 2972
rect 12400 2932 12406 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 12437 2935 12495 2941
rect 14835 2944 15117 2972
rect 9950 2904 9956 2916
rect 8904 2876 8949 2904
rect 9048 2876 9812 2904
rect 9911 2876 9956 2904
rect 8904 2864 8910 2876
rect 9048 2836 9076 2876
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 10045 2907 10103 2913
rect 10045 2873 10057 2907
rect 10091 2873 10103 2907
rect 10045 2867 10103 2873
rect 10965 2907 11023 2913
rect 10965 2873 10977 2907
rect 11011 2873 11023 2907
rect 10965 2867 11023 2873
rect 11241 2907 11299 2913
rect 11241 2873 11253 2907
rect 11287 2904 11299 2907
rect 11330 2904 11336 2916
rect 11287 2876 11336 2904
rect 11287 2873 11299 2876
rect 11241 2867 11299 2873
rect 7800 2808 9076 2836
rect 7800 2796 7806 2808
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 10060 2836 10088 2867
rect 9180 2808 10088 2836
rect 10980 2836 11008 2867
rect 11330 2864 11336 2876
rect 11388 2864 11394 2916
rect 12158 2864 12164 2916
rect 12216 2904 12222 2916
rect 12713 2907 12771 2913
rect 12713 2904 12725 2907
rect 12216 2876 12725 2904
rect 12216 2864 12222 2876
rect 12713 2873 12725 2876
rect 12759 2873 12771 2907
rect 12713 2867 12771 2873
rect 12805 2907 12863 2913
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 12986 2904 12992 2916
rect 12851 2876 12992 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 12986 2864 12992 2876
rect 13044 2864 13050 2916
rect 13725 2907 13783 2913
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 13814 2904 13820 2916
rect 13771 2876 13820 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 13814 2864 13820 2876
rect 13872 2864 13878 2916
rect 13998 2904 14004 2916
rect 13959 2876 14004 2904
rect 13998 2864 14004 2876
rect 14056 2864 14062 2916
rect 14093 2907 14151 2913
rect 14093 2873 14105 2907
rect 14139 2904 14151 2907
rect 14274 2904 14280 2916
rect 14139 2876 14280 2904
rect 14139 2873 14151 2876
rect 14093 2867 14151 2873
rect 14274 2864 14280 2876
rect 14332 2904 14338 2916
rect 14550 2904 14556 2916
rect 14332 2876 14556 2904
rect 14332 2864 14338 2876
rect 14550 2864 14556 2876
rect 14608 2864 14614 2916
rect 14835 2836 14863 2944
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 15565 2975 15623 2981
rect 15565 2941 15577 2975
rect 15611 2941 15623 2975
rect 15565 2935 15623 2941
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 15013 2907 15071 2913
rect 15013 2873 15025 2907
rect 15059 2904 15071 2907
rect 15746 2904 15752 2916
rect 15059 2876 15752 2904
rect 15059 2873 15071 2876
rect 15013 2867 15071 2873
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 16117 2907 16175 2913
rect 16117 2873 16129 2907
rect 16163 2904 16175 2907
rect 16206 2904 16212 2916
rect 16163 2876 16212 2904
rect 16163 2873 16175 2876
rect 16117 2867 16175 2873
rect 16206 2864 16212 2876
rect 16264 2864 16270 2916
rect 17037 2907 17095 2913
rect 17037 2873 17049 2907
rect 17083 2904 17095 2907
rect 17236 2904 17264 2935
rect 17494 2932 17500 2984
rect 17552 2972 17558 2984
rect 18064 2981 18092 3012
rect 17589 2975 17647 2981
rect 17589 2972 17601 2975
rect 17552 2944 17601 2972
rect 17552 2932 17558 2944
rect 17589 2941 17601 2944
rect 17635 2941 17647 2975
rect 17589 2935 17647 2941
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2972 18107 2975
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 18095 2944 18429 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18417 2941 18429 2944
rect 18463 2941 18475 2975
rect 18417 2935 18475 2941
rect 17083 2876 17264 2904
rect 17083 2873 17095 2876
rect 17037 2867 17095 2873
rect 10980 2808 14863 2836
rect 15289 2839 15347 2845
rect 9180 2796 9186 2808
rect 15289 2805 15301 2839
rect 15335 2836 15347 2839
rect 15562 2836 15568 2848
rect 15335 2808 15568 2836
rect 15335 2805 15347 2808
rect 15289 2799 15347 2805
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 17770 2836 17776 2848
rect 17731 2808 17776 2836
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 17862 2796 17868 2848
rect 17920 2836 17926 2848
rect 18233 2839 18291 2845
rect 18233 2836 18245 2839
rect 17920 2808 18245 2836
rect 17920 2796 17926 2808
rect 18233 2805 18245 2808
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 4890 2632 4896 2644
rect 3283 2604 4896 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2496 1639 2499
rect 1946 2496 1952 2508
rect 1627 2468 1952 2496
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2130 2496 2136 2508
rect 2091 2468 2136 2496
rect 2130 2456 2136 2468
rect 2188 2456 2194 2508
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 3252 2496 3280 2595
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 7650 2592 7656 2644
rect 7708 2632 7714 2644
rect 8297 2635 8355 2641
rect 8297 2632 8309 2635
rect 7708 2604 8309 2632
rect 7708 2592 7714 2604
rect 8297 2601 8309 2604
rect 8343 2601 8355 2635
rect 8297 2595 8355 2601
rect 8478 2592 8484 2644
rect 8536 2592 8542 2644
rect 8846 2592 8852 2644
rect 8904 2632 8910 2644
rect 8987 2635 9045 2641
rect 8987 2632 8999 2635
rect 8904 2604 8999 2632
rect 8904 2592 8910 2604
rect 8987 2601 8999 2604
rect 9033 2601 9045 2635
rect 15151 2635 15209 2641
rect 15151 2632 15163 2635
rect 8987 2595 9045 2601
rect 14016 2604 15163 2632
rect 3510 2524 3516 2576
rect 3568 2524 3574 2576
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 5629 2567 5687 2573
rect 5629 2564 5641 2567
rect 5592 2536 5641 2564
rect 5592 2524 5598 2536
rect 5629 2533 5641 2536
rect 5675 2533 5687 2567
rect 8496 2564 8524 2592
rect 11333 2567 11391 2573
rect 5629 2527 5687 2533
rect 6472 2536 8800 2564
rect 2823 2468 3280 2496
rect 3329 2499 3387 2505
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 3329 2465 3341 2499
rect 3375 2496 3387 2499
rect 3528 2496 3556 2524
rect 3375 2468 3556 2496
rect 4065 2499 4123 2505
rect 3375 2465 3387 2468
rect 3329 2459 3387 2465
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 5258 2496 5264 2508
rect 4111 2468 5264 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 5353 2499 5411 2505
rect 5353 2465 5365 2499
rect 5399 2496 5411 2499
rect 6270 2496 6276 2508
rect 5399 2468 6276 2496
rect 5399 2465 5411 2468
rect 5353 2459 5411 2465
rect 6270 2456 6276 2468
rect 6328 2456 6334 2508
rect 6472 2505 6500 2536
rect 6457 2499 6515 2505
rect 6457 2465 6469 2499
rect 6503 2465 6515 2499
rect 6457 2459 6515 2465
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6788 2468 6929 2496
rect 6788 2456 6794 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 7282 2496 7288 2508
rect 7243 2468 7288 2496
rect 6917 2459 6975 2465
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 7742 2496 7748 2508
rect 7703 2468 7748 2496
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8386 2496 8392 2508
rect 8159 2468 8392 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 658 2388 664 2440
rect 716 2428 722 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 716 2400 1777 2428
rect 716 2388 722 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 1118 2320 1124 2372
rect 1176 2360 1182 2372
rect 2332 2360 2360 2391
rect 3528 2360 3556 2391
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 4249 2431 4307 2437
rect 4249 2428 4261 2431
rect 3660 2400 4261 2428
rect 3660 2388 3666 2400
rect 4249 2397 4261 2400
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 8128 2428 8156 2459
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 8570 2496 8576 2508
rect 8527 2468 8576 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 8772 2496 8800 2536
rect 9968 2536 10824 2564
rect 8884 2499 8942 2505
rect 8884 2496 8896 2499
rect 8772 2468 8896 2496
rect 8884 2465 8896 2468
rect 8930 2496 8942 2499
rect 9122 2496 9128 2508
rect 8930 2468 9128 2496
rect 8930 2465 8942 2468
rect 8884 2459 8942 2465
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 9674 2496 9680 2508
rect 9263 2468 9680 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 9968 2505 9996 2536
rect 9953 2499 10011 2505
rect 9953 2465 9965 2499
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 10410 2456 10416 2508
rect 10468 2496 10474 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 10468 2468 10701 2496
rect 10468 2456 10474 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 10689 2459 10747 2465
rect 7699 2400 8156 2428
rect 9769 2431 9827 2437
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 9769 2397 9781 2431
rect 9815 2428 9827 2431
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9815 2400 10333 2428
rect 9815 2397 9827 2400
rect 9769 2391 9827 2397
rect 10321 2397 10333 2400
rect 10367 2428 10379 2431
rect 10502 2428 10508 2440
rect 10367 2400 10508 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 1176 2332 2360 2360
rect 2792 2332 3556 2360
rect 1176 2320 1182 2332
rect 1670 2252 1676 2304
rect 1728 2292 1734 2304
rect 2792 2292 2820 2332
rect 7098 2320 7104 2372
rect 7156 2360 7162 2372
rect 7929 2363 7987 2369
rect 7929 2360 7941 2363
rect 7156 2332 7941 2360
rect 7156 2320 7162 2332
rect 7929 2329 7941 2332
rect 7975 2329 7987 2363
rect 7929 2323 7987 2329
rect 8110 2320 8116 2372
rect 8168 2360 8174 2372
rect 8665 2363 8723 2369
rect 8665 2360 8677 2363
rect 8168 2332 8677 2360
rect 8168 2320 8174 2332
rect 8665 2329 8677 2332
rect 8711 2329 8723 2363
rect 8665 2323 8723 2329
rect 10796 2304 10824 2536
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 11882 2564 11888 2576
rect 11379 2536 11888 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 11882 2524 11888 2536
rect 11940 2524 11946 2576
rect 12250 2564 12256 2576
rect 12211 2536 12256 2564
rect 12250 2524 12256 2536
rect 12308 2524 12314 2576
rect 12710 2524 12716 2576
rect 12768 2564 12774 2576
rect 14016 2573 14044 2604
rect 15151 2601 15163 2604
rect 15197 2601 15209 2635
rect 15151 2595 15209 2601
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 12768 2536 12817 2564
rect 12768 2524 12774 2536
rect 12805 2533 12817 2536
rect 12851 2533 12863 2567
rect 12805 2527 12863 2533
rect 14001 2567 14059 2573
rect 14001 2533 14013 2567
rect 14047 2533 14059 2567
rect 14001 2527 14059 2533
rect 14550 2524 14556 2576
rect 14608 2564 14614 2576
rect 15654 2564 15660 2576
rect 14608 2536 15091 2564
rect 15615 2536 15660 2564
rect 14608 2524 14614 2536
rect 15063 2505 15091 2536
rect 15654 2524 15660 2536
rect 15712 2524 15718 2576
rect 15746 2524 15752 2576
rect 15804 2564 15810 2576
rect 15804 2536 17080 2564
rect 15804 2524 15810 2536
rect 17052 2505 17080 2536
rect 17126 2524 17132 2576
rect 17184 2564 17190 2576
rect 18325 2567 18383 2573
rect 18325 2564 18337 2567
rect 17184 2536 18337 2564
rect 17184 2524 17190 2536
rect 15048 2499 15106 2505
rect 15048 2465 15060 2499
rect 15094 2465 15106 2499
rect 15048 2459 15106 2465
rect 16669 2499 16727 2505
rect 16669 2465 16681 2499
rect 16715 2465 16727 2499
rect 16669 2459 16727 2465
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2465 17095 2499
rect 17037 2459 17095 2465
rect 17405 2499 17463 2505
rect 17405 2465 17417 2499
rect 17451 2496 17463 2499
rect 17586 2496 17592 2508
rect 17451 2468 17592 2496
rect 17451 2465 17463 2468
rect 17405 2459 17463 2465
rect 11241 2431 11299 2437
rect 11241 2397 11253 2431
rect 11287 2428 11299 2431
rect 11606 2428 11612 2440
rect 11287 2400 11612 2428
rect 11287 2397 11299 2400
rect 11241 2391 11299 2397
rect 11606 2388 11612 2400
rect 11664 2428 11670 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 11664 2400 12357 2428
rect 11664 2388 11670 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12492 2400 12725 2428
rect 12492 2388 12498 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 12526 2320 12532 2372
rect 12584 2360 12590 2372
rect 13004 2360 13032 2391
rect 13630 2388 13636 2440
rect 13688 2428 13694 2440
rect 13909 2431 13967 2437
rect 13909 2428 13921 2431
rect 13688 2400 13921 2428
rect 13688 2388 13694 2400
rect 13909 2397 13921 2400
rect 13955 2397 13967 2431
rect 13909 2391 13967 2397
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14185 2431 14243 2437
rect 14185 2428 14197 2431
rect 14056 2400 14197 2428
rect 14056 2388 14062 2400
rect 14185 2397 14197 2400
rect 14231 2397 14243 2431
rect 14185 2391 14243 2397
rect 15194 2388 15200 2440
rect 15252 2428 15258 2440
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 15252 2400 15577 2428
rect 15252 2388 15258 2400
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2397 15899 2431
rect 16684 2428 16712 2459
rect 17586 2456 17592 2468
rect 17644 2456 17650 2508
rect 17788 2505 17816 2536
rect 18325 2533 18337 2536
rect 18371 2533 18383 2567
rect 18325 2527 18383 2533
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2465 17831 2499
rect 17773 2459 17831 2465
rect 15841 2391 15899 2397
rect 15948 2400 16712 2428
rect 12584 2332 13032 2360
rect 12584 2320 12590 2332
rect 15378 2320 15384 2372
rect 15436 2360 15442 2372
rect 15856 2360 15884 2391
rect 15436 2332 15884 2360
rect 15436 2320 15442 2332
rect 2958 2292 2964 2304
rect 1728 2264 2820 2292
rect 2919 2264 2964 2292
rect 1728 2252 1734 2264
rect 2958 2252 2964 2264
rect 3016 2252 3022 2304
rect 6638 2292 6644 2304
rect 6599 2264 6644 2292
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 9122 2252 9128 2304
rect 9180 2292 9186 2304
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 9180 2264 9413 2292
rect 9180 2252 9186 2264
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 9401 2255 9459 2261
rect 10137 2295 10195 2301
rect 10137 2261 10149 2295
rect 10183 2292 10195 2295
rect 10594 2292 10600 2304
rect 10183 2264 10600 2292
rect 10183 2261 10195 2264
rect 10137 2255 10195 2261
rect 10594 2252 10600 2264
rect 10652 2252 10658 2304
rect 10778 2292 10784 2304
rect 10739 2264 10784 2292
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 13814 2252 13820 2304
rect 13872 2292 13878 2304
rect 15948 2292 15976 2400
rect 13872 2264 15976 2292
rect 13872 2252 13878 2264
rect 16666 2252 16672 2304
rect 16724 2292 16730 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16724 2264 16865 2292
rect 16724 2252 16730 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 17126 2252 17132 2304
rect 17184 2292 17190 2304
rect 17221 2295 17279 2301
rect 17221 2292 17233 2295
rect 17184 2264 17233 2292
rect 17184 2252 17190 2264
rect 17221 2261 17233 2264
rect 17267 2261 17279 2295
rect 17586 2292 17592 2304
rect 17547 2264 17592 2292
rect 17221 2255 17279 2261
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 17957 2295 18015 2301
rect 17957 2292 17969 2295
rect 17920 2264 17969 2292
rect 17920 2252 17926 2264
rect 17957 2261 17969 2264
rect 18003 2261 18015 2295
rect 17957 2255 18015 2261
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 10778 2048 10784 2100
rect 10836 2088 10842 2100
rect 16206 2088 16212 2100
rect 10836 2060 16212 2088
rect 10836 2048 10842 2060
rect 16206 2048 16212 2060
rect 16264 2048 16270 2100
rect 5258 1980 5264 2032
rect 5316 2020 5322 2032
rect 14458 2020 14464 2032
rect 5316 1992 14464 2020
rect 5316 1980 5322 1992
rect 14458 1980 14464 1992
rect 14516 1980 14522 2032
rect 12618 1708 12624 1760
rect 12676 1748 12682 1760
rect 13630 1748 13636 1760
rect 12676 1720 13636 1748
rect 12676 1708 12682 1720
rect 13630 1708 13636 1720
rect 13688 1708 13694 1760
<< via1 >>
rect 3332 15240 3384 15292
rect 6184 15240 6236 15292
rect 3240 15172 3292 15224
rect 6552 15172 6604 15224
rect 10968 15172 11020 15224
rect 15844 15172 15896 15224
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 4068 14424 4120 14476
rect 8484 14424 8536 14476
rect 3332 14356 3384 14408
rect 11796 14356 11848 14408
rect 3792 14288 3844 14340
rect 14188 14288 14240 14340
rect 14280 14288 14332 14340
rect 19616 14288 19668 14340
rect 2412 14220 2464 14272
rect 3608 14220 3660 14272
rect 12440 14220 12492 14272
rect 18328 14220 18380 14272
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 296 14016 348 14068
rect 1584 13948 1636 14000
rect 2872 14016 2924 14068
rect 3608 14059 3660 14068
rect 3608 14025 3617 14059
rect 3617 14025 3651 14059
rect 3651 14025 3660 14059
rect 3608 14016 3660 14025
rect 3792 14059 3844 14068
rect 3792 14025 3801 14059
rect 3801 14025 3835 14059
rect 3835 14025 3844 14059
rect 3792 14016 3844 14025
rect 2228 13948 2280 14000
rect 940 13880 992 13932
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 2412 13855 2464 13864
rect 2412 13821 2421 13855
rect 2421 13821 2455 13855
rect 2455 13821 2464 13855
rect 2412 13812 2464 13821
rect 6000 13948 6052 14000
rect 6736 14016 6788 14068
rect 10876 13948 10928 14000
rect 15752 13948 15804 14000
rect 13268 13880 13320 13932
rect 14280 13880 14332 13932
rect 6092 13812 6144 13864
rect 6276 13812 6328 13864
rect 14372 13812 14424 13864
rect 15108 13812 15160 13864
rect 15660 13880 15712 13932
rect 15568 13855 15620 13864
rect 15568 13821 15577 13855
rect 15577 13821 15611 13855
rect 15611 13821 15620 13855
rect 15568 13812 15620 13821
rect 16396 13812 16448 13864
rect 4252 13744 4304 13796
rect 8668 13676 8720 13728
rect 10692 13676 10744 13728
rect 13820 13719 13872 13728
rect 13820 13685 13829 13719
rect 13829 13685 13863 13719
rect 13863 13685 13872 13719
rect 13820 13676 13872 13685
rect 15384 13719 15436 13728
rect 15384 13685 15393 13719
rect 15393 13685 15427 13719
rect 15427 13685 15436 13719
rect 15384 13676 15436 13685
rect 15476 13676 15528 13728
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 3332 13472 3384 13524
rect 4436 13472 4488 13524
rect 9312 13472 9364 13524
rect 11152 13472 11204 13524
rect 2044 13404 2096 13456
rect 4804 13404 4856 13456
rect 15384 13472 15436 13524
rect 13176 13404 13228 13456
rect 14372 13404 14424 13456
rect 12256 13336 12308 13388
rect 11244 13268 11296 13320
rect 12072 13268 12124 13320
rect 12532 13336 12584 13388
rect 14740 13336 14792 13388
rect 17684 13336 17736 13388
rect 15660 13268 15712 13320
rect 16396 13268 16448 13320
rect 1676 13200 1728 13252
rect 9404 13200 9456 13252
rect 17040 13200 17092 13252
rect 10600 13132 10652 13184
rect 14096 13132 14148 13184
rect 14188 13132 14240 13184
rect 18972 13132 19024 13184
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 2780 12928 2832 12980
rect 2504 12792 2556 12844
rect 10232 12928 10284 12980
rect 13452 12928 13504 12980
rect 5448 12860 5500 12912
rect 15476 12860 15528 12912
rect 3148 12835 3200 12844
rect 3148 12801 3157 12835
rect 3157 12801 3191 12835
rect 3191 12801 3200 12835
rect 3148 12792 3200 12801
rect 3516 12792 3568 12844
rect 13820 12792 13872 12844
rect 10784 12724 10836 12776
rect 11244 12724 11296 12776
rect 11888 12724 11940 12776
rect 2320 12631 2372 12640
rect 2320 12597 2329 12631
rect 2329 12597 2363 12631
rect 2363 12597 2372 12631
rect 2320 12588 2372 12597
rect 2412 12588 2464 12640
rect 10876 12588 10928 12640
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 2320 12384 2372 12436
rect 2228 12316 2280 12368
rect 7748 12384 7800 12436
rect 8024 12384 8076 12436
rect 13912 12384 13964 12436
rect 14556 12384 14608 12436
rect 2504 12316 2556 12368
rect 3240 12316 3292 12368
rect 10968 12316 11020 12368
rect 2320 12248 2372 12300
rect 2596 12248 2648 12300
rect 6368 12248 6420 12300
rect 1860 12044 1912 12096
rect 4988 12180 5040 12232
rect 3516 12112 3568 12164
rect 3792 12044 3844 12096
rect 16580 12112 16632 12164
rect 7288 12044 7340 12096
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 2320 11883 2372 11892
rect 2320 11849 2329 11883
rect 2329 11849 2363 11883
rect 2363 11849 2372 11883
rect 2320 11840 2372 11849
rect 2688 11840 2740 11892
rect 2504 11704 2556 11756
rect 3240 11747 3292 11756
rect 3240 11713 3249 11747
rect 3249 11713 3283 11747
rect 3283 11713 3292 11747
rect 3240 11704 3292 11713
rect 7748 11840 7800 11892
rect 15568 11840 15620 11892
rect 16212 11840 16264 11892
rect 8392 11747 8444 11756
rect 1860 11679 1912 11688
rect 1860 11645 1869 11679
rect 1869 11645 1903 11679
rect 1903 11645 1912 11679
rect 1860 11636 1912 11645
rect 3148 11636 3200 11688
rect 3240 11568 3292 11620
rect 3792 11679 3844 11688
rect 3792 11645 3826 11679
rect 3826 11645 3844 11679
rect 3792 11636 3844 11645
rect 4988 11679 5040 11688
rect 4988 11645 4997 11679
rect 4997 11645 5031 11679
rect 5031 11645 5040 11679
rect 4988 11636 5040 11645
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 7748 11679 7800 11688
rect 7748 11645 7757 11679
rect 7757 11645 7791 11679
rect 7791 11645 7800 11679
rect 7748 11636 7800 11645
rect 14648 11636 14700 11688
rect 1676 11500 1728 11552
rect 1860 11500 1912 11552
rect 2596 11500 2648 11552
rect 6368 11543 6420 11552
rect 6368 11509 6377 11543
rect 6377 11509 6411 11543
rect 6411 11509 6420 11543
rect 6368 11500 6420 11509
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 1952 11296 2004 11348
rect 1584 11228 1636 11280
rect 3240 11296 3292 11348
rect 3516 11339 3568 11348
rect 3516 11305 3525 11339
rect 3525 11305 3559 11339
rect 3559 11305 3568 11339
rect 3516 11296 3568 11305
rect 3700 11296 3752 11348
rect 17316 11296 17368 11348
rect 2228 11203 2280 11212
rect 2228 11169 2237 11203
rect 2237 11169 2271 11203
rect 2271 11169 2280 11203
rect 2228 11160 2280 11169
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 3792 11228 3844 11280
rect 4988 11228 5040 11280
rect 6828 11228 6880 11280
rect 7288 11228 7340 11280
rect 2780 11024 2832 11076
rect 3516 11160 3568 11212
rect 6644 11203 6696 11212
rect 6644 11169 6653 11203
rect 6653 11169 6687 11203
rect 6687 11169 6696 11203
rect 6644 11160 6696 11169
rect 10416 11160 10468 11212
rect 11336 11160 11388 11212
rect 12624 11160 12676 11212
rect 13268 11160 13320 11212
rect 4344 11092 4396 11144
rect 5908 11092 5960 11144
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 3240 11024 3292 11076
rect 3424 11024 3476 11076
rect 6092 11024 6144 11076
rect 5724 10999 5776 11008
rect 5724 10965 5733 10999
rect 5733 10965 5767 10999
rect 5767 10965 5776 10999
rect 5724 10956 5776 10965
rect 8208 10999 8260 11008
rect 8208 10965 8217 10999
rect 8217 10965 8251 10999
rect 8251 10965 8260 10999
rect 8208 10956 8260 10965
rect 8300 10956 8352 11008
rect 11888 10956 11940 11008
rect 13544 11092 13596 11144
rect 15200 11092 15252 11144
rect 13636 11024 13688 11076
rect 16120 11024 16172 11076
rect 17776 11024 17828 11076
rect 16304 10956 16356 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 2228 10752 2280 10804
rect 1768 10684 1820 10736
rect 2688 10752 2740 10804
rect 3056 10752 3108 10804
rect 3792 10752 3844 10804
rect 6184 10752 6236 10804
rect 6644 10752 6696 10804
rect 8760 10727 8812 10736
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 8760 10693 8769 10727
rect 8769 10693 8803 10727
rect 8803 10693 8812 10727
rect 8760 10684 8812 10693
rect 5264 10659 5316 10668
rect 1860 10455 1912 10464
rect 1860 10421 1869 10455
rect 1869 10421 1903 10455
rect 1903 10421 1912 10455
rect 1860 10412 1912 10421
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 3240 10480 3292 10532
rect 4068 10480 4120 10532
rect 4896 10480 4948 10532
rect 5724 10616 5776 10668
rect 6184 10616 6236 10668
rect 10784 10752 10836 10804
rect 18052 10752 18104 10804
rect 11336 10616 11388 10668
rect 13636 10684 13688 10736
rect 12716 10616 12768 10668
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 13544 10616 13596 10625
rect 16580 10616 16632 10668
rect 6828 10548 6880 10600
rect 7380 10591 7432 10600
rect 7380 10557 7389 10591
rect 7389 10557 7423 10591
rect 7423 10557 7432 10591
rect 7380 10548 7432 10557
rect 8208 10548 8260 10600
rect 11888 10548 11940 10600
rect 12624 10548 12676 10600
rect 13820 10548 13872 10600
rect 14924 10548 14976 10600
rect 2504 10412 2556 10464
rect 3056 10412 3108 10464
rect 4804 10412 4856 10464
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 10416 10480 10468 10532
rect 11060 10523 11112 10532
rect 11060 10489 11069 10523
rect 11069 10489 11103 10523
rect 11103 10489 11112 10523
rect 11060 10480 11112 10489
rect 11704 10480 11756 10532
rect 5908 10412 5960 10464
rect 7472 10412 7524 10464
rect 10140 10412 10192 10464
rect 10324 10412 10376 10464
rect 10508 10412 10560 10464
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 12164 10412 12216 10464
rect 13268 10480 13320 10532
rect 15016 10480 15068 10532
rect 15568 10480 15620 10532
rect 17776 10523 17828 10532
rect 17776 10489 17785 10523
rect 17785 10489 17819 10523
rect 17819 10489 17828 10523
rect 17776 10480 17828 10489
rect 13360 10412 13412 10464
rect 13544 10412 13596 10464
rect 13728 10412 13780 10464
rect 16304 10455 16356 10464
rect 16304 10421 16313 10455
rect 16313 10421 16347 10455
rect 16347 10421 16356 10455
rect 16304 10412 16356 10421
rect 16672 10455 16724 10464
rect 16672 10421 16681 10455
rect 16681 10421 16715 10455
rect 16715 10421 16724 10455
rect 16672 10412 16724 10421
rect 16948 10412 17000 10464
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 18328 10412 18380 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 2320 10208 2372 10260
rect 4068 10208 4120 10260
rect 1860 10140 1912 10192
rect 2872 10140 2924 10192
rect 5080 10208 5132 10260
rect 5724 10208 5776 10260
rect 6276 10208 6328 10260
rect 6644 10251 6696 10260
rect 6644 10217 6653 10251
rect 6653 10217 6687 10251
rect 6687 10217 6696 10251
rect 6644 10208 6696 10217
rect 3700 10072 3752 10124
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 3516 9868 3568 9920
rect 4344 9868 4396 9920
rect 4620 9911 4672 9920
rect 4620 9877 4629 9911
rect 4629 9877 4663 9911
rect 4663 9877 4672 9911
rect 4620 9868 4672 9877
rect 5540 10140 5592 10192
rect 5908 10140 5960 10192
rect 5632 10072 5684 10124
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 6276 10072 6328 10124
rect 6460 10072 6512 10124
rect 8300 10208 8352 10260
rect 10876 10208 10928 10260
rect 11704 10208 11756 10260
rect 12164 10208 12216 10260
rect 14924 10208 14976 10260
rect 15016 10208 15068 10260
rect 16580 10208 16632 10260
rect 16948 10251 17000 10260
rect 16948 10217 16957 10251
rect 16957 10217 16991 10251
rect 16991 10217 17000 10251
rect 16948 10208 17000 10217
rect 17408 10251 17460 10260
rect 17408 10217 17417 10251
rect 17417 10217 17451 10251
rect 17451 10217 17460 10251
rect 17408 10208 17460 10217
rect 17500 10208 17552 10260
rect 10508 10140 10560 10192
rect 10784 10140 10836 10192
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 6184 10004 6236 10056
rect 7288 10072 7340 10124
rect 7380 10072 7432 10124
rect 7840 10115 7892 10124
rect 7840 10081 7874 10115
rect 7874 10081 7892 10115
rect 7840 10072 7892 10081
rect 8760 10072 8812 10124
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 11888 10072 11940 10124
rect 13268 10072 13320 10124
rect 13820 10072 13872 10124
rect 16212 10140 16264 10192
rect 17776 10140 17828 10192
rect 11336 10004 11388 10056
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 13636 10004 13688 10056
rect 16580 10072 16632 10124
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 17960 10072 18012 10124
rect 14924 10004 14976 10056
rect 9404 9868 9456 9920
rect 9772 9911 9824 9920
rect 9772 9877 9781 9911
rect 9781 9877 9815 9911
rect 9815 9877 9824 9911
rect 9772 9868 9824 9877
rect 12164 9911 12216 9920
rect 12164 9877 12173 9911
rect 12173 9877 12207 9911
rect 12207 9877 12216 9911
rect 12164 9868 12216 9877
rect 13544 9868 13596 9920
rect 16672 9936 16724 9988
rect 16856 9868 16908 9920
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 2872 9707 2924 9716
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 3700 9707 3752 9716
rect 3700 9673 3709 9707
rect 3709 9673 3743 9707
rect 3743 9673 3752 9707
rect 3700 9664 3752 9673
rect 3792 9664 3844 9716
rect 12440 9664 12492 9716
rect 12624 9664 12676 9716
rect 13268 9664 13320 9716
rect 13820 9664 13872 9716
rect 15200 9664 15252 9716
rect 2596 9596 2648 9648
rect 3516 9596 3568 9648
rect 5448 9596 5500 9648
rect 5632 9596 5684 9648
rect 3240 9528 3292 9580
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 4712 9528 4764 9580
rect 4804 9528 4856 9580
rect 5356 9528 5408 9580
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 6644 9528 6696 9580
rect 7288 9528 7340 9580
rect 7840 9528 7892 9580
rect 9220 9528 9272 9580
rect 10324 9571 10376 9580
rect 4620 9460 4672 9512
rect 5080 9460 5132 9512
rect 7104 9460 7156 9512
rect 8024 9460 8076 9512
rect 9864 9460 9916 9512
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 11612 9528 11664 9580
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 13636 9596 13688 9648
rect 13268 9528 13320 9580
rect 13728 9528 13780 9580
rect 14464 9596 14516 9648
rect 16212 9596 16264 9648
rect 15016 9528 15068 9580
rect 11520 9460 11572 9512
rect 12164 9460 12216 9512
rect 13544 9460 13596 9512
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 16212 9460 16264 9512
rect 1860 9367 1912 9376
rect 1860 9333 1869 9367
rect 1869 9333 1903 9367
rect 1903 9333 1912 9367
rect 1860 9324 1912 9333
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 3424 9324 3476 9376
rect 3976 9324 4028 9376
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 5264 9324 5316 9376
rect 5540 9324 5592 9376
rect 5632 9324 5684 9376
rect 6460 9324 6512 9376
rect 6736 9324 6788 9376
rect 10232 9392 10284 9444
rect 13084 9435 13136 9444
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 13084 9401 13093 9435
rect 13093 9401 13127 9435
rect 13127 9401 13136 9435
rect 13084 9392 13136 9401
rect 15016 9392 15068 9444
rect 17408 9664 17460 9716
rect 16948 9596 17000 9648
rect 17684 9596 17736 9648
rect 16580 9528 16632 9580
rect 17592 9460 17644 9512
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 16488 9392 16540 9444
rect 17408 9392 17460 9444
rect 17500 9435 17552 9444
rect 17500 9401 17509 9435
rect 17509 9401 17543 9435
rect 17543 9401 17552 9435
rect 17500 9392 17552 9401
rect 17868 9392 17920 9444
rect 13636 9324 13688 9376
rect 13728 9324 13780 9376
rect 15200 9324 15252 9376
rect 16580 9324 16632 9376
rect 17224 9324 17276 9376
rect 17776 9324 17828 9376
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 3608 9163 3660 9172
rect 3608 9129 3617 9163
rect 3617 9129 3651 9163
rect 3651 9129 3660 9163
rect 3608 9120 3660 9129
rect 4160 9120 4212 9172
rect 3424 9052 3476 9104
rect 5172 9120 5224 9172
rect 5448 9120 5500 9172
rect 5908 9120 5960 9172
rect 5356 9052 5408 9104
rect 6368 9052 6420 9104
rect 6736 9120 6788 9172
rect 17592 9163 17644 9172
rect 2688 8984 2740 9036
rect 5816 8984 5868 9036
rect 1492 8916 1544 8968
rect 1768 8916 1820 8968
rect 4252 8916 4304 8968
rect 4988 8959 5040 8968
rect 4988 8925 4997 8959
rect 4997 8925 5031 8959
rect 5031 8925 5040 8959
rect 4988 8916 5040 8925
rect 5080 8916 5132 8968
rect 6276 8916 6328 8968
rect 7012 9052 7064 9104
rect 9680 9052 9732 9104
rect 10140 9095 10192 9104
rect 10140 9061 10149 9095
rect 10149 9061 10183 9095
rect 10183 9061 10192 9095
rect 10140 9052 10192 9061
rect 10232 9052 10284 9104
rect 16488 9052 16540 9104
rect 17592 9129 17601 9163
rect 17601 9129 17635 9163
rect 17635 9129 17644 9163
rect 17592 9120 17644 9129
rect 17868 9120 17920 9172
rect 18696 9120 18748 9172
rect 17500 9052 17552 9104
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 8944 8984 8996 9036
rect 9128 9027 9180 9036
rect 9128 8993 9137 9027
rect 9137 8993 9171 9027
rect 9171 8993 9180 9027
rect 9128 8984 9180 8993
rect 9956 8984 10008 9036
rect 10600 9027 10652 9036
rect 6644 8916 6696 8968
rect 9220 8959 9272 8968
rect 5540 8848 5592 8900
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 9496 8916 9548 8968
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 11612 8984 11664 9036
rect 11704 8984 11756 9036
rect 13268 8984 13320 9036
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 18144 9052 18196 9104
rect 5908 8780 5960 8832
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 8760 8823 8812 8832
rect 8760 8789 8769 8823
rect 8769 8789 8803 8823
rect 8803 8789 8812 8823
rect 8760 8780 8812 8789
rect 8944 8848 8996 8900
rect 10232 8848 10284 8900
rect 9680 8823 9732 8832
rect 9680 8789 9689 8823
rect 9689 8789 9723 8823
rect 9723 8789 9732 8823
rect 9680 8780 9732 8789
rect 9772 8780 9824 8832
rect 10416 8848 10468 8900
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 14004 8916 14056 8968
rect 15200 8916 15252 8968
rect 17316 8959 17368 8968
rect 17316 8925 17325 8959
rect 17325 8925 17359 8959
rect 17359 8925 17368 8959
rect 17316 8916 17368 8925
rect 17500 8916 17552 8968
rect 10784 8780 10836 8832
rect 12440 8780 12492 8832
rect 12716 8848 12768 8900
rect 16488 8848 16540 8900
rect 13912 8780 13964 8832
rect 14924 8780 14976 8832
rect 16304 8780 16356 8832
rect 17960 8780 18012 8832
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 2688 8576 2740 8628
rect 3424 8576 3476 8628
rect 3792 8576 3844 8628
rect 5356 8619 5408 8628
rect 5356 8585 5365 8619
rect 5365 8585 5399 8619
rect 5399 8585 5408 8619
rect 5356 8576 5408 8585
rect 11060 8576 11112 8628
rect 11520 8576 11572 8628
rect 13360 8576 13412 8628
rect 3332 8551 3384 8560
rect 3332 8517 3341 8551
rect 3341 8517 3375 8551
rect 3375 8517 3384 8551
rect 3332 8508 3384 8517
rect 4620 8508 4672 8560
rect 5908 8508 5960 8560
rect 6368 8551 6420 8560
rect 6368 8517 6377 8551
rect 6377 8517 6411 8551
rect 6411 8517 6420 8551
rect 6368 8508 6420 8517
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 6092 8483 6144 8492
rect 6092 8449 6101 8483
rect 6101 8449 6135 8483
rect 6135 8449 6144 8483
rect 6092 8440 6144 8449
rect 7380 8440 7432 8492
rect 7656 8440 7708 8492
rect 5632 8372 5684 8424
rect 7748 8372 7800 8424
rect 8760 8508 8812 8560
rect 8852 8508 8904 8560
rect 9680 8508 9732 8560
rect 12624 8508 12676 8560
rect 8576 8440 8628 8492
rect 9404 8440 9456 8492
rect 9772 8440 9824 8492
rect 10048 8440 10100 8492
rect 10416 8440 10468 8492
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 13820 8508 13872 8560
rect 13544 8483 13596 8492
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 8668 8372 8720 8424
rect 10232 8372 10284 8424
rect 10876 8372 10928 8424
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 11336 8372 11388 8424
rect 16672 8576 16724 8628
rect 17224 8576 17276 8628
rect 17132 8508 17184 8560
rect 14004 8440 14056 8492
rect 16488 8483 16540 8492
rect 16488 8449 16497 8483
rect 16497 8449 16531 8483
rect 16531 8449 16540 8483
rect 16488 8440 16540 8449
rect 16764 8440 16816 8492
rect 17316 8483 17368 8492
rect 2504 8304 2556 8356
rect 3792 8347 3844 8356
rect 3792 8313 3826 8347
rect 3826 8313 3844 8347
rect 3792 8304 3844 8313
rect 5356 8304 5408 8356
rect 8852 8304 8904 8356
rect 8944 8304 8996 8356
rect 10968 8304 11020 8356
rect 11060 8304 11112 8356
rect 16672 8304 16724 8356
rect 17316 8449 17325 8483
rect 17325 8449 17359 8483
rect 17359 8449 17368 8483
rect 17316 8440 17368 8449
rect 17868 8508 17920 8560
rect 18144 8440 18196 8492
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 17592 8415 17644 8424
rect 17592 8381 17601 8415
rect 17601 8381 17635 8415
rect 17635 8381 17644 8415
rect 17592 8372 17644 8381
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 4896 8279 4948 8288
rect 4896 8245 4905 8279
rect 4905 8245 4939 8279
rect 4939 8245 4948 8279
rect 4896 8236 4948 8245
rect 5540 8279 5592 8288
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 5540 8236 5592 8245
rect 5908 8279 5960 8288
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 5908 8236 5960 8245
rect 6736 8236 6788 8288
rect 7564 8279 7616 8288
rect 7564 8245 7573 8279
rect 7573 8245 7607 8279
rect 7607 8245 7616 8279
rect 7564 8236 7616 8245
rect 7656 8236 7708 8288
rect 8668 8236 8720 8288
rect 10232 8279 10284 8288
rect 10232 8245 10241 8279
rect 10241 8245 10275 8279
rect 10275 8245 10284 8279
rect 10232 8236 10284 8245
rect 10416 8236 10468 8288
rect 10784 8236 10836 8288
rect 15568 8236 15620 8288
rect 17040 8236 17092 8288
rect 17960 8304 18012 8356
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 5540 8032 5592 8084
rect 6184 8032 6236 8084
rect 7656 8032 7708 8084
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 10232 8032 10284 8084
rect 11612 8075 11664 8084
rect 11612 8041 11621 8075
rect 11621 8041 11655 8075
rect 11655 8041 11664 8075
rect 11612 8032 11664 8041
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 2964 7896 3016 7948
rect 2504 7828 2556 7880
rect 3424 7896 3476 7948
rect 4436 7939 4488 7948
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 3792 7828 3844 7880
rect 6092 7964 6144 8016
rect 7564 7964 7616 8016
rect 8024 7964 8076 8016
rect 10416 7964 10468 8016
rect 5540 7896 5592 7948
rect 5632 7896 5684 7948
rect 6552 7896 6604 7948
rect 12348 7964 12400 8016
rect 12716 7964 12768 8016
rect 13176 7964 13228 8016
rect 15108 8032 15160 8084
rect 15476 8032 15528 8084
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 16764 8032 16816 8084
rect 17592 8032 17644 8084
rect 13728 7964 13780 8016
rect 17040 7964 17092 8016
rect 10968 7896 11020 7948
rect 11980 7896 12032 7948
rect 13636 7896 13688 7948
rect 15108 7896 15160 7948
rect 16304 7896 16356 7948
rect 17500 7896 17552 7948
rect 18236 7939 18288 7948
rect 18236 7905 18245 7939
rect 18245 7905 18279 7939
rect 18279 7905 18288 7939
rect 18236 7896 18288 7905
rect 4896 7828 4948 7880
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 1860 7692 1912 7701
rect 2044 7735 2096 7744
rect 2044 7701 2053 7735
rect 2053 7701 2087 7735
rect 2087 7701 2096 7735
rect 2044 7692 2096 7701
rect 2320 7692 2372 7744
rect 2412 7692 2464 7744
rect 4528 7692 4580 7744
rect 8208 7828 8260 7880
rect 8576 7828 8628 7880
rect 8760 7828 8812 7880
rect 9772 7828 9824 7880
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 6736 7760 6788 7812
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 8668 7692 8720 7744
rect 9680 7692 9732 7744
rect 12164 7828 12216 7880
rect 12440 7828 12492 7880
rect 12992 7828 13044 7880
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 14924 7828 14976 7880
rect 17224 7828 17276 7880
rect 11612 7760 11664 7812
rect 16580 7760 16632 7812
rect 18512 7760 18564 7812
rect 11704 7735 11756 7744
rect 11704 7701 11713 7735
rect 11713 7701 11747 7735
rect 11747 7701 11756 7735
rect 11704 7692 11756 7701
rect 12164 7735 12216 7744
rect 12164 7701 12173 7735
rect 12173 7701 12207 7735
rect 12207 7701 12216 7735
rect 12164 7692 12216 7701
rect 12900 7692 12952 7744
rect 17592 7735 17644 7744
rect 17592 7701 17601 7735
rect 17601 7701 17635 7735
rect 17635 7701 17644 7735
rect 17592 7692 17644 7701
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 1676 7488 1728 7540
rect 2136 7488 2188 7540
rect 2964 7531 3016 7540
rect 2964 7497 2973 7531
rect 2973 7497 3007 7531
rect 3007 7497 3016 7531
rect 2964 7488 3016 7497
rect 4436 7488 4488 7540
rect 5540 7531 5592 7540
rect 5540 7497 5549 7531
rect 5549 7497 5583 7531
rect 5583 7497 5592 7531
rect 5540 7488 5592 7497
rect 2412 7395 2464 7404
rect 2412 7361 2421 7395
rect 2421 7361 2455 7395
rect 2455 7361 2464 7395
rect 2412 7352 2464 7361
rect 2688 7352 2740 7404
rect 2320 7327 2372 7336
rect 2320 7293 2329 7327
rect 2329 7293 2363 7327
rect 2363 7293 2372 7327
rect 2320 7284 2372 7293
rect 6276 7420 6328 7472
rect 8208 7488 8260 7540
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 5632 7352 5684 7404
rect 6092 7395 6144 7404
rect 6092 7361 6101 7395
rect 6101 7361 6135 7395
rect 6135 7361 6144 7395
rect 6092 7352 6144 7361
rect 6644 7395 6696 7404
rect 6644 7361 6653 7395
rect 6653 7361 6687 7395
rect 6687 7361 6696 7395
rect 6644 7352 6696 7361
rect 8024 7352 8076 7404
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 11520 7488 11572 7540
rect 12348 7488 12400 7540
rect 9956 7420 10008 7472
rect 5908 7284 5960 7336
rect 6460 7284 6512 7336
rect 7472 7284 7524 7336
rect 2044 7216 2096 7268
rect 4160 7216 4212 7268
rect 4620 7216 4672 7268
rect 5356 7216 5408 7268
rect 1768 7191 1820 7200
rect 1768 7157 1777 7191
rect 1777 7157 1811 7191
rect 1811 7157 1820 7191
rect 1768 7148 1820 7157
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 2688 7148 2740 7200
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 8392 7216 8444 7268
rect 5172 7148 5224 7157
rect 5816 7148 5868 7200
rect 6644 7148 6696 7200
rect 8024 7191 8076 7200
rect 8024 7157 8033 7191
rect 8033 7157 8067 7191
rect 8067 7157 8076 7191
rect 8024 7148 8076 7157
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8760 7327 8812 7336
rect 8760 7293 8794 7327
rect 8794 7293 8812 7327
rect 8760 7284 8812 7293
rect 9680 7284 9732 7336
rect 10508 7284 10560 7336
rect 13176 7420 13228 7472
rect 15108 7488 15160 7540
rect 15476 7488 15528 7540
rect 16488 7531 16540 7540
rect 16488 7497 16497 7531
rect 16497 7497 16531 7531
rect 16531 7497 16540 7531
rect 16488 7488 16540 7497
rect 17040 7420 17092 7472
rect 18236 7420 18288 7472
rect 12348 7352 12400 7404
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 17316 7352 17368 7404
rect 10784 7216 10836 7268
rect 12164 7216 12216 7268
rect 8116 7148 8168 7157
rect 9680 7148 9732 7200
rect 10232 7148 10284 7200
rect 10416 7148 10468 7200
rect 11520 7191 11572 7200
rect 11520 7157 11529 7191
rect 11529 7157 11563 7191
rect 11563 7157 11572 7191
rect 11520 7148 11572 7157
rect 12716 7284 12768 7336
rect 13912 7284 13964 7336
rect 14648 7284 14700 7336
rect 15660 7284 15712 7336
rect 17224 7284 17276 7336
rect 17592 7327 17644 7336
rect 17592 7293 17601 7327
rect 17601 7293 17635 7327
rect 17635 7293 17644 7327
rect 17592 7284 17644 7293
rect 17960 7284 18012 7336
rect 18420 7284 18472 7336
rect 12808 7259 12860 7268
rect 12808 7225 12817 7259
rect 12817 7225 12851 7259
rect 12851 7225 12860 7259
rect 12808 7216 12860 7225
rect 16672 7216 16724 7268
rect 13360 7148 13412 7200
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 13728 7148 13780 7200
rect 17592 7148 17644 7200
rect 17776 7191 17828 7200
rect 17776 7157 17785 7191
rect 17785 7157 17819 7191
rect 17819 7157 17828 7191
rect 17776 7148 17828 7157
rect 17868 7148 17920 7200
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 18972 7055 19024 7064
rect 18972 7021 18981 7055
rect 18981 7021 19015 7055
rect 19015 7021 19024 7055
rect 18972 7012 19024 7021
rect 2688 6944 2740 6996
rect 3332 6987 3384 6996
rect 2504 6876 2556 6928
rect 3332 6953 3341 6987
rect 3341 6953 3375 6987
rect 3375 6953 3384 6987
rect 3332 6944 3384 6953
rect 4344 6944 4396 6996
rect 5172 6944 5224 6996
rect 5632 6987 5684 6996
rect 5632 6953 5641 6987
rect 5641 6953 5675 6987
rect 5675 6953 5684 6987
rect 5632 6944 5684 6953
rect 6460 6944 6512 6996
rect 8116 6987 8168 6996
rect 8116 6953 8125 6987
rect 8125 6953 8159 6987
rect 8159 6953 8168 6987
rect 8116 6944 8168 6953
rect 2688 6808 2740 6860
rect 4160 6808 4212 6860
rect 4528 6851 4580 6860
rect 4528 6817 4562 6851
rect 4562 6817 4580 6851
rect 4528 6808 4580 6817
rect 2044 6672 2096 6724
rect 2228 6715 2280 6724
rect 2228 6681 2237 6715
rect 2237 6681 2271 6715
rect 2271 6681 2280 6715
rect 2228 6672 2280 6681
rect 2780 6672 2832 6724
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 3700 6740 3752 6792
rect 5356 6876 5408 6928
rect 10508 6944 10560 6996
rect 10600 6944 10652 6996
rect 13360 6987 13412 6996
rect 8392 6876 8444 6928
rect 11980 6876 12032 6928
rect 5448 6808 5500 6860
rect 6092 6808 6144 6860
rect 6828 6808 6880 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 3332 6672 3384 6724
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 5356 6672 5408 6724
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6736 6783 6788 6792
rect 6460 6740 6512 6749
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7932 6740 7984 6792
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 7012 6672 7064 6724
rect 10600 6808 10652 6860
rect 12440 6876 12492 6928
rect 13360 6953 13369 6987
rect 13369 6953 13403 6987
rect 13403 6953 13412 6987
rect 13360 6944 13412 6953
rect 13544 6944 13596 6996
rect 16120 6944 16172 6996
rect 16488 6944 16540 6996
rect 18420 6987 18472 6996
rect 18420 6953 18429 6987
rect 18429 6953 18463 6987
rect 18463 6953 18472 6987
rect 18420 6944 18472 6953
rect 14648 6876 14700 6928
rect 17224 6919 17276 6928
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 11796 6740 11848 6792
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 12716 6783 12768 6792
rect 12716 6749 12725 6783
rect 12725 6749 12759 6783
rect 12759 6749 12768 6783
rect 12716 6740 12768 6749
rect 14004 6740 14056 6792
rect 16120 6808 16172 6860
rect 17224 6885 17233 6919
rect 17233 6885 17267 6919
rect 17267 6885 17276 6919
rect 17224 6876 17276 6885
rect 14924 6740 14976 6792
rect 15108 6740 15160 6792
rect 5540 6604 5592 6656
rect 8576 6604 8628 6656
rect 9956 6672 10008 6724
rect 9496 6604 9548 6656
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 11888 6604 11940 6613
rect 12164 6647 12216 6656
rect 12164 6613 12173 6647
rect 12173 6613 12207 6647
rect 12207 6613 12216 6647
rect 12164 6604 12216 6613
rect 12808 6604 12860 6656
rect 17040 6808 17092 6860
rect 17408 6808 17460 6860
rect 17316 6783 17368 6792
rect 17316 6749 17325 6783
rect 17325 6749 17359 6783
rect 17359 6749 17368 6783
rect 17316 6740 17368 6749
rect 16672 6715 16724 6724
rect 16672 6681 16681 6715
rect 16681 6681 16715 6715
rect 16715 6681 16724 6715
rect 16672 6672 16724 6681
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 3240 6400 3292 6452
rect 6644 6443 6696 6452
rect 3608 6332 3660 6384
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 7012 6400 7064 6452
rect 8024 6400 8076 6452
rect 13544 6400 13596 6452
rect 14924 6400 14976 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 18604 6400 18656 6452
rect 2044 6264 2096 6316
rect 3608 6239 3660 6248
rect 1860 6103 1912 6112
rect 1860 6069 1869 6103
rect 1869 6069 1903 6103
rect 1903 6069 1912 6103
rect 1860 6060 1912 6069
rect 3240 6128 3292 6180
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 4712 6264 4764 6316
rect 6460 6264 6512 6316
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 7564 6264 7616 6316
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 9680 6332 9732 6384
rect 10508 6332 10560 6384
rect 11888 6332 11940 6384
rect 12348 6332 12400 6384
rect 12164 6264 12216 6316
rect 16120 6332 16172 6384
rect 13360 6307 13412 6316
rect 13360 6273 13369 6307
rect 13369 6273 13403 6307
rect 13403 6273 13412 6307
rect 13360 6264 13412 6273
rect 13912 6307 13964 6316
rect 13912 6273 13921 6307
rect 13921 6273 13955 6307
rect 13955 6273 13964 6307
rect 13912 6264 13964 6273
rect 16488 6264 16540 6316
rect 17316 6332 17368 6384
rect 16672 6264 16724 6316
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 3792 6128 3844 6180
rect 4528 6060 4580 6112
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 5724 6060 5776 6069
rect 5908 6128 5960 6180
rect 6644 6128 6696 6180
rect 8944 6196 8996 6248
rect 9496 6239 9548 6248
rect 9496 6205 9505 6239
rect 9505 6205 9539 6239
rect 9539 6205 9548 6239
rect 9496 6196 9548 6205
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 11888 6196 11940 6248
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 15844 6196 15896 6248
rect 18052 6239 18104 6248
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 6552 6060 6604 6112
rect 11704 6060 11756 6112
rect 12348 6060 12400 6112
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 14004 6128 14056 6180
rect 12440 6060 12492 6069
rect 15292 6060 15344 6112
rect 15752 6060 15804 6112
rect 15936 6060 15988 6112
rect 16120 6060 16172 6112
rect 16580 6060 16632 6112
rect 18236 6103 18288 6112
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 2596 5899 2648 5908
rect 2596 5865 2605 5899
rect 2605 5865 2639 5899
rect 2639 5865 2648 5899
rect 2596 5856 2648 5865
rect 2780 5856 2832 5908
rect 3424 5856 3476 5908
rect 5080 5856 5132 5908
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 5724 5856 5776 5908
rect 2688 5788 2740 5840
rect 2780 5652 2832 5704
rect 3240 5788 3292 5840
rect 3148 5720 3200 5772
rect 5540 5788 5592 5840
rect 3608 5695 3660 5704
rect 3608 5661 3617 5695
rect 3617 5661 3651 5695
rect 3651 5661 3660 5695
rect 3608 5652 3660 5661
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 6368 5720 6420 5772
rect 7380 5856 7432 5908
rect 8576 5856 8628 5908
rect 11520 5856 11572 5908
rect 12440 5856 12492 5908
rect 14004 5856 14056 5908
rect 15200 5856 15252 5908
rect 15660 5899 15712 5908
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 15844 5899 15896 5908
rect 15844 5865 15853 5899
rect 15853 5865 15887 5899
rect 15887 5865 15896 5899
rect 15844 5856 15896 5865
rect 17500 5899 17552 5908
rect 7380 5763 7432 5772
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 7380 5720 7432 5729
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 10324 5720 10376 5772
rect 8484 5652 8536 5704
rect 1860 5559 1912 5568
rect 1860 5525 1869 5559
rect 1869 5525 1903 5559
rect 1903 5525 1912 5559
rect 1860 5516 1912 5525
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 3148 5559 3200 5568
rect 3148 5525 3157 5559
rect 3157 5525 3191 5559
rect 3191 5525 3200 5559
rect 3148 5516 3200 5525
rect 5816 5516 5868 5568
rect 12348 5720 12400 5772
rect 15752 5720 15804 5772
rect 16672 5720 16724 5772
rect 11980 5652 12032 5704
rect 16488 5695 16540 5704
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 12348 5584 12400 5636
rect 16212 5584 16264 5636
rect 17500 5865 17509 5899
rect 17509 5865 17543 5899
rect 17543 5865 17552 5899
rect 17500 5856 17552 5865
rect 17684 5763 17736 5772
rect 17684 5729 17693 5763
rect 17693 5729 17727 5763
rect 17727 5729 17736 5763
rect 17684 5720 17736 5729
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 18052 5627 18104 5636
rect 18052 5593 18061 5627
rect 18061 5593 18095 5627
rect 18095 5593 18104 5627
rect 18052 5584 18104 5593
rect 18144 5584 18196 5636
rect 11336 5559 11388 5568
rect 11336 5525 11345 5559
rect 11345 5525 11379 5559
rect 11379 5525 11388 5559
rect 11336 5516 11388 5525
rect 13820 5516 13872 5568
rect 17960 5516 18012 5568
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 3608 5312 3660 5364
rect 4344 5312 4396 5364
rect 11336 5312 11388 5364
rect 16212 5355 16264 5364
rect 16212 5321 16221 5355
rect 16221 5321 16255 5355
rect 16255 5321 16264 5355
rect 16212 5312 16264 5321
rect 16672 5355 16724 5364
rect 16672 5321 16681 5355
rect 16681 5321 16715 5355
rect 16715 5321 16724 5355
rect 16672 5312 16724 5321
rect 2596 5287 2648 5296
rect 2596 5253 2605 5287
rect 2605 5253 2639 5287
rect 2639 5253 2648 5287
rect 2596 5244 2648 5253
rect 6460 5244 6512 5296
rect 16120 5244 16172 5296
rect 3148 5176 3200 5228
rect 4528 5176 4580 5228
rect 4712 5219 4764 5228
rect 4712 5185 4721 5219
rect 4721 5185 4755 5219
rect 4755 5185 4764 5219
rect 4712 5176 4764 5185
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 11244 5219 11296 5228
rect 11244 5185 11253 5219
rect 11253 5185 11287 5219
rect 11287 5185 11296 5219
rect 11244 5176 11296 5185
rect 14280 5219 14332 5228
rect 1400 5040 1452 5092
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 2780 5040 2832 5092
rect 5080 5108 5132 5160
rect 7380 5108 7432 5160
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 15568 5176 15620 5228
rect 16488 5176 16540 5228
rect 16948 5176 17000 5228
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 17776 5176 17828 5228
rect 4344 5040 4396 5092
rect 5356 5040 5408 5092
rect 5448 5040 5500 5092
rect 4528 5015 4580 5024
rect 4528 4981 4537 5015
rect 4537 4981 4571 5015
rect 4571 4981 4580 5015
rect 4528 4972 4580 4981
rect 7472 4972 7524 5024
rect 17408 5108 17460 5160
rect 17500 5108 17552 5160
rect 9772 5040 9824 5092
rect 10968 5040 11020 5092
rect 9680 4972 9732 5024
rect 10600 5015 10652 5024
rect 10600 4981 10609 5015
rect 10609 4981 10643 5015
rect 10643 4981 10652 5015
rect 10600 4972 10652 4981
rect 13176 4972 13228 5024
rect 13360 5083 13412 5092
rect 13360 5049 13369 5083
rect 13369 5049 13403 5083
rect 13403 5049 13412 5083
rect 13360 5040 13412 5049
rect 13544 4972 13596 5024
rect 16948 4972 17000 5024
rect 17500 4972 17552 5024
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 2228 4811 2280 4820
rect 2228 4777 2237 4811
rect 2237 4777 2271 4811
rect 2271 4777 2280 4811
rect 2228 4768 2280 4777
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 5172 4768 5224 4820
rect 5356 4811 5408 4820
rect 5356 4777 5365 4811
rect 5365 4777 5399 4811
rect 5399 4777 5408 4811
rect 5356 4768 5408 4777
rect 6092 4768 6144 4820
rect 10324 4768 10376 4820
rect 10692 4768 10744 4820
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 12164 4768 12216 4820
rect 1860 4471 1912 4480
rect 1860 4437 1869 4471
rect 1869 4437 1903 4471
rect 1903 4437 1912 4471
rect 1860 4428 1912 4437
rect 4804 4632 4856 4684
rect 4896 4564 4948 4616
rect 8300 4675 8352 4684
rect 8300 4641 8334 4675
rect 8334 4641 8352 4675
rect 10600 4700 10652 4752
rect 13360 4768 13412 4820
rect 16580 4811 16632 4820
rect 16580 4777 16589 4811
rect 16589 4777 16623 4811
rect 16623 4777 16632 4811
rect 16580 4768 16632 4777
rect 16948 4811 17000 4820
rect 16948 4777 16957 4811
rect 16957 4777 16991 4811
rect 16991 4777 17000 4811
rect 16948 4768 17000 4777
rect 15476 4743 15528 4752
rect 15476 4709 15485 4743
rect 15485 4709 15519 4743
rect 15519 4709 15528 4743
rect 15476 4700 15528 4709
rect 16396 4743 16448 4752
rect 16396 4709 16405 4743
rect 16405 4709 16439 4743
rect 16439 4709 16448 4743
rect 16396 4700 16448 4709
rect 16488 4700 16540 4752
rect 16856 4700 16908 4752
rect 8300 4632 8352 4641
rect 5356 4564 5408 4616
rect 6092 4564 6144 4616
rect 7104 4564 7156 4616
rect 9680 4564 9732 4616
rect 4528 4496 4580 4548
rect 7932 4496 7984 4548
rect 9772 4496 9824 4548
rect 13176 4632 13228 4684
rect 14004 4632 14056 4684
rect 17408 4675 17460 4684
rect 17408 4641 17417 4675
rect 17417 4641 17451 4675
rect 17451 4641 17460 4675
rect 17408 4632 17460 4641
rect 17960 4632 18012 4684
rect 18420 4632 18472 4684
rect 14924 4564 14976 4616
rect 12624 4496 12676 4548
rect 5172 4428 5224 4480
rect 11612 4471 11664 4480
rect 11612 4437 11621 4471
rect 11621 4437 11655 4471
rect 11655 4437 11664 4471
rect 11612 4428 11664 4437
rect 14280 4428 14332 4480
rect 14648 4428 14700 4480
rect 17224 4607 17276 4616
rect 17224 4573 17233 4607
rect 17233 4573 17267 4607
rect 17267 4573 17276 4607
rect 17224 4564 17276 4573
rect 18144 4496 18196 4548
rect 17868 4428 17920 4480
rect 18420 4471 18472 4480
rect 18420 4437 18429 4471
rect 18429 4437 18463 4471
rect 18463 4437 18472 4471
rect 18420 4428 18472 4437
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 2228 4156 2280 4208
rect 3056 4088 3108 4140
rect 3240 4088 3292 4140
rect 5172 4224 5224 4276
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 5724 4088 5776 4140
rect 8300 4224 8352 4276
rect 6092 4131 6144 4140
rect 6092 4097 6101 4131
rect 6101 4097 6135 4131
rect 6135 4097 6144 4131
rect 6092 4088 6144 4097
rect 8576 4199 8628 4208
rect 8576 4165 8585 4199
rect 8585 4165 8619 4199
rect 8619 4165 8628 4199
rect 8576 4156 8628 4165
rect 10784 4156 10836 4208
rect 5264 4020 5316 4072
rect 6644 4020 6696 4072
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 2320 3884 2372 3893
rect 4436 3952 4488 4004
rect 8024 3952 8076 4004
rect 4528 3884 4580 3936
rect 4620 3884 4672 3936
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 9864 4088 9916 4140
rect 14372 4224 14424 4276
rect 11520 4156 11572 4208
rect 14004 4156 14056 4208
rect 13084 4088 13136 4140
rect 13360 4131 13412 4140
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 14372 4088 14424 4140
rect 14832 4131 14884 4140
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 16304 4088 16356 4140
rect 17224 4131 17276 4140
rect 17224 4097 17233 4131
rect 17233 4097 17267 4131
rect 17267 4097 17276 4131
rect 17224 4088 17276 4097
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 10140 4020 10192 4072
rect 10508 4020 10560 4072
rect 10600 4020 10652 4072
rect 10784 4020 10836 4072
rect 11428 4020 11480 4072
rect 11612 4020 11664 4072
rect 9220 3952 9272 4004
rect 12164 4020 12216 4072
rect 17500 4020 17552 4072
rect 11888 3995 11940 4004
rect 11888 3961 11897 3995
rect 11897 3961 11931 3995
rect 11931 3961 11940 3995
rect 11888 3952 11940 3961
rect 9772 3884 9824 3936
rect 10968 3884 11020 3936
rect 11152 3884 11204 3936
rect 14280 3995 14332 4004
rect 14280 3961 14289 3995
rect 14289 3961 14323 3995
rect 14323 3961 14332 3995
rect 14280 3952 14332 3961
rect 14740 3952 14792 4004
rect 16396 3995 16448 4004
rect 14004 3884 14056 3936
rect 16396 3961 16405 3995
rect 16405 3961 16439 3995
rect 16439 3961 16448 3995
rect 16396 3952 16448 3961
rect 16120 3884 16172 3936
rect 18696 3952 18748 4004
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 1676 3680 1728 3732
rect 2412 3680 2464 3732
rect 7288 3680 7340 3732
rect 8024 3723 8076 3732
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 8116 3680 8168 3732
rect 8576 3680 8628 3732
rect 10140 3680 10192 3732
rect 10232 3680 10284 3732
rect 12164 3680 12216 3732
rect 13452 3680 13504 3732
rect 14372 3680 14424 3732
rect 16856 3723 16908 3732
rect 16856 3689 16865 3723
rect 16865 3689 16899 3723
rect 16899 3689 16908 3723
rect 16856 3680 16908 3689
rect 17500 3680 17552 3732
rect 7472 3612 7524 3664
rect 5264 3544 5316 3596
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 7288 3544 7340 3596
rect 6644 3519 6696 3528
rect 6644 3485 6653 3519
rect 6653 3485 6687 3519
rect 6687 3485 6696 3519
rect 6644 3476 6696 3485
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 5172 3340 5224 3392
rect 10416 3612 10468 3664
rect 11612 3612 11664 3664
rect 9220 3544 9272 3596
rect 9680 3544 9732 3596
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 9864 3544 9916 3553
rect 10140 3544 10192 3596
rect 11888 3587 11940 3596
rect 8852 3519 8904 3528
rect 8852 3485 8861 3519
rect 8861 3485 8895 3519
rect 8895 3485 8904 3519
rect 8852 3476 8904 3485
rect 8760 3408 8812 3460
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 11980 3544 12032 3596
rect 12440 3544 12492 3596
rect 12992 3544 13044 3596
rect 14096 3544 14148 3596
rect 14556 3544 14608 3596
rect 14740 3544 14792 3596
rect 16120 3612 16172 3664
rect 16396 3612 16448 3664
rect 15476 3544 15528 3596
rect 16212 3544 16264 3596
rect 16304 3587 16356 3596
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 16764 3544 16816 3596
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 14924 3476 14976 3528
rect 17224 3544 17276 3596
rect 17776 3544 17828 3596
rect 8668 3340 8720 3392
rect 9772 3340 9824 3392
rect 13176 3408 13228 3460
rect 15200 3408 15252 3460
rect 19156 3408 19208 3460
rect 11152 3340 11204 3392
rect 11888 3340 11940 3392
rect 12716 3340 12768 3392
rect 13636 3383 13688 3392
rect 13636 3349 13645 3383
rect 13645 3349 13679 3383
rect 13679 3349 13688 3383
rect 13636 3340 13688 3349
rect 15660 3340 15712 3392
rect 17408 3340 17460 3392
rect 17592 3340 17644 3392
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 18604 3340 18656 3392
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 2964 3179 3016 3188
rect 2228 3111 2280 3120
rect 2228 3077 2237 3111
rect 2237 3077 2271 3111
rect 2271 3077 2280 3111
rect 2228 3068 2280 3077
rect 1676 2975 1728 2984
rect 1676 2941 1685 2975
rect 1685 2941 1719 2975
rect 1719 2941 1728 2975
rect 1676 2932 1728 2941
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 3148 3136 3200 3188
rect 7564 3136 7616 3188
rect 8116 3179 8168 3188
rect 5816 3068 5868 3120
rect 6736 3068 6788 3120
rect 8116 3145 8125 3179
rect 8125 3145 8159 3179
rect 8159 3145 8168 3179
rect 8116 3136 8168 3145
rect 8392 3136 8444 3188
rect 12440 3136 12492 3188
rect 12900 3136 12952 3188
rect 8576 3068 8628 3120
rect 8852 3068 8904 3120
rect 14280 3068 14332 3120
rect 14832 3068 14884 3120
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 204 2796 256 2848
rect 1400 2796 1452 2848
rect 1860 2839 1912 2848
rect 1860 2805 1869 2839
rect 1869 2805 1903 2839
rect 1903 2805 1912 2839
rect 1860 2796 1912 2805
rect 2872 2932 2924 2984
rect 7472 2975 7524 2984
rect 7472 2941 7481 2975
rect 7481 2941 7515 2975
rect 7515 2941 7524 2975
rect 7472 2932 7524 2941
rect 2228 2864 2280 2916
rect 5540 2864 5592 2916
rect 2964 2796 3016 2848
rect 7748 2796 7800 2848
rect 8852 2907 8904 2916
rect 8852 2873 8861 2907
rect 8861 2873 8895 2907
rect 8895 2873 8904 2907
rect 10600 3000 10652 3052
rect 11244 3000 11296 3052
rect 16120 3068 16172 3120
rect 12348 2932 12400 2984
rect 19616 3068 19668 3120
rect 9956 2907 10008 2916
rect 8852 2864 8904 2873
rect 9956 2873 9965 2907
rect 9965 2873 9999 2907
rect 9999 2873 10008 2907
rect 9956 2864 10008 2873
rect 9128 2796 9180 2848
rect 11336 2864 11388 2916
rect 12164 2864 12216 2916
rect 12992 2864 13044 2916
rect 13820 2864 13872 2916
rect 14004 2907 14056 2916
rect 14004 2873 14013 2907
rect 14013 2873 14047 2907
rect 14047 2873 14056 2907
rect 14004 2864 14056 2873
rect 14280 2864 14332 2916
rect 14556 2864 14608 2916
rect 15752 2864 15804 2916
rect 16212 2864 16264 2916
rect 17500 2932 17552 2984
rect 15568 2796 15620 2848
rect 17776 2839 17828 2848
rect 17776 2805 17785 2839
rect 17785 2805 17819 2839
rect 17819 2805 17828 2839
rect 17776 2796 17828 2805
rect 17868 2796 17920 2848
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 1952 2456 2004 2508
rect 2136 2499 2188 2508
rect 2136 2465 2145 2499
rect 2145 2465 2179 2499
rect 2179 2465 2188 2499
rect 2136 2456 2188 2465
rect 4896 2592 4948 2644
rect 7656 2592 7708 2644
rect 8484 2592 8536 2644
rect 8852 2592 8904 2644
rect 3516 2524 3568 2576
rect 5540 2524 5592 2576
rect 5264 2456 5316 2508
rect 6276 2456 6328 2508
rect 6736 2456 6788 2508
rect 7288 2499 7340 2508
rect 7288 2465 7297 2499
rect 7297 2465 7331 2499
rect 7331 2465 7340 2499
rect 7288 2456 7340 2465
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 664 2388 716 2440
rect 1124 2320 1176 2372
rect 3608 2388 3660 2440
rect 8392 2456 8444 2508
rect 8576 2456 8628 2508
rect 9128 2456 9180 2508
rect 9680 2456 9732 2508
rect 10416 2456 10468 2508
rect 10508 2388 10560 2440
rect 1676 2252 1728 2304
rect 7104 2320 7156 2372
rect 8116 2320 8168 2372
rect 11888 2524 11940 2576
rect 12256 2567 12308 2576
rect 12256 2533 12265 2567
rect 12265 2533 12299 2567
rect 12299 2533 12308 2567
rect 12256 2524 12308 2533
rect 12716 2524 12768 2576
rect 14556 2524 14608 2576
rect 15660 2567 15712 2576
rect 15660 2533 15669 2567
rect 15669 2533 15703 2567
rect 15703 2533 15712 2567
rect 15660 2524 15712 2533
rect 15752 2524 15804 2576
rect 17132 2524 17184 2576
rect 11612 2388 11664 2440
rect 12440 2388 12492 2440
rect 12532 2320 12584 2372
rect 13636 2388 13688 2440
rect 14004 2388 14056 2440
rect 15200 2388 15252 2440
rect 17592 2456 17644 2508
rect 15384 2320 15436 2372
rect 2964 2295 3016 2304
rect 2964 2261 2973 2295
rect 2973 2261 3007 2295
rect 3007 2261 3016 2295
rect 2964 2252 3016 2261
rect 6644 2295 6696 2304
rect 6644 2261 6653 2295
rect 6653 2261 6687 2295
rect 6687 2261 6696 2295
rect 6644 2252 6696 2261
rect 9128 2252 9180 2304
rect 10600 2252 10652 2304
rect 10784 2295 10836 2304
rect 10784 2261 10793 2295
rect 10793 2261 10827 2295
rect 10827 2261 10836 2295
rect 10784 2252 10836 2261
rect 13820 2252 13872 2304
rect 16672 2252 16724 2304
rect 17132 2252 17184 2304
rect 17592 2295 17644 2304
rect 17592 2261 17601 2295
rect 17601 2261 17635 2295
rect 17635 2261 17644 2295
rect 17592 2252 17644 2261
rect 17868 2252 17920 2304
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 10784 2048 10836 2100
rect 16212 2048 16264 2100
rect 5264 1980 5316 2032
rect 14464 1980 14516 2032
rect 12624 1708 12676 1760
rect 13636 1708 13688 1760
<< metal2 >>
rect 294 16400 350 17200
rect 938 16400 994 17200
rect 1582 16400 1638 17200
rect 2226 16400 2282 17200
rect 2778 16416 2834 16425
rect 308 14074 336 16400
rect 296 14068 348 14074
rect 296 14010 348 14016
rect 952 13938 980 16400
rect 1596 14006 1624 16400
rect 2240 14006 2268 16400
rect 2870 16400 2926 17200
rect 3330 16824 3386 16833
rect 3330 16759 3386 16768
rect 2778 16351 2834 16360
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 1584 14000 1636 14006
rect 1584 13942 1636 13948
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 940 13932 992 13938
rect 940 13874 992 13880
rect 2424 13870 2452 14214
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 1688 13258 1716 13806
rect 2056 13462 2084 13806
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 2792 12986 2820 16351
rect 2884 14074 2912 16400
rect 3054 16008 3110 16017
rect 3054 15943 3110 15952
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2870 13968 2926 13977
rect 2870 13903 2926 13912
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2332 12442 2360 12582
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1872 11694 1900 12038
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1582 11384 1638 11393
rect 1582 11319 1638 11328
rect 1596 11286 1624 11319
rect 1584 11280 1636 11286
rect 1584 11222 1636 11228
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1504 8498 1532 8910
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1688 7546 1716 11494
rect 1872 11354 1900 11494
rect 2240 11370 2268 12310
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 11898 2360 12242
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2148 11342 2268 11370
rect 1768 10736 1820 10742
rect 1768 10678 1820 10684
rect 1780 8974 1808 10678
rect 1964 10674 1992 11290
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1872 10198 1900 10406
rect 1860 10192 1912 10198
rect 1860 10134 1912 10140
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1872 8129 1900 9318
rect 1858 8120 1914 8129
rect 1858 8055 1914 8064
rect 2148 7970 2176 11342
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2240 10810 2268 11154
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2332 10266 2360 11086
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2424 9500 2452 12582
rect 2516 12374 2544 12786
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2516 11762 2544 12310
rect 2596 12300 2648 12306
rect 2648 12260 2728 12288
rect 2596 12242 2648 12248
rect 2700 11898 2728 12260
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2516 10470 2544 11698
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2608 9654 2636 11494
rect 2700 10810 2728 11834
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2792 9602 2820 11018
rect 2884 10198 2912 13903
rect 2962 12744 3018 12753
rect 2962 12679 3018 12688
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2884 9722 2912 9998
rect 2976 9874 3004 12679
rect 3068 10810 3096 15943
rect 3238 15600 3294 15609
rect 3238 15535 3294 15544
rect 3252 15230 3280 15535
rect 3344 15298 3372 16759
rect 3514 16400 3570 17200
rect 4158 16400 4214 17200
rect 4802 16400 4858 17200
rect 5446 16400 5502 17200
rect 6090 16400 6146 17200
rect 6734 16400 6790 17200
rect 7378 16400 7434 17200
rect 8022 16400 8078 17200
rect 8666 16400 8722 17200
rect 9310 16400 9366 17200
rect 9954 16400 10010 17200
rect 10598 16400 10654 17200
rect 11242 16400 11298 17200
rect 11886 16400 11942 17200
rect 12530 16400 12586 17200
rect 13174 16400 13230 17200
rect 13818 16400 13874 17200
rect 14462 16400 14518 17200
rect 15106 16400 15162 17200
rect 15750 16400 15806 17200
rect 15842 16416 15898 16425
rect 3332 15292 3384 15298
rect 3332 15234 3384 15240
rect 3240 15224 3292 15230
rect 3240 15166 3292 15172
rect 3330 15192 3386 15201
rect 3330 15127 3386 15136
rect 3344 14414 3372 15127
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3330 13560 3386 13569
rect 3330 13495 3332 13504
rect 3384 13495 3386 13504
rect 3332 13466 3384 13472
rect 3330 13152 3386 13161
rect 3330 13087 3386 13096
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3160 11694 3188 12786
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 3252 11762 3280 12310
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3252 11354 3280 11562
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3344 11234 3372 13087
rect 3528 12850 3556 16400
rect 4066 14784 4122 14793
rect 4066 14719 4122 14728
rect 4080 14482 4108 14719
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3620 14074 3648 14214
rect 3804 14074 3832 14282
rect 4172 14260 4200 16400
rect 4342 14376 4398 14385
rect 4342 14311 4398 14320
rect 4172 14232 4292 14260
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 4264 13802 4292 14232
rect 4252 13796 4304 13802
rect 4252 13738 4304 13744
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3422 12336 3478 12345
rect 3422 12271 3478 12280
rect 3160 11206 3372 11234
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 3068 10062 3096 10406
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 2976 9846 3096 9874
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2792 9574 2912 9602
rect 2780 9512 2832 9518
rect 2424 9472 2636 9500
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 8537 2268 9318
rect 2226 8528 2282 8537
rect 2226 8463 2282 8472
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2148 7942 2268 7970
rect 1860 7744 1912 7750
rect 1858 7712 1860 7721
rect 2044 7744 2096 7750
rect 1912 7712 1914 7721
rect 2044 7686 2096 7692
rect 1858 7647 1914 7656
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 2056 7274 2084 7686
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1400 5092 1452 5098
rect 1400 5034 1452 5040
rect 1412 2854 1440 5034
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1688 2990 1716 3674
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 216 800 244 2790
rect 664 2440 716 2446
rect 664 2382 716 2388
rect 676 800 704 2382
rect 1124 2372 1176 2378
rect 1124 2314 1176 2320
rect 1136 800 1164 2314
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 1688 800 1716 2246
rect 1780 1057 1808 7142
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 6497 1900 6598
rect 1858 6488 1914 6497
rect 1858 6423 1914 6432
rect 1860 6112 1912 6118
rect 1858 6080 1860 6089
rect 1912 6080 1914 6089
rect 1858 6015 1914 6024
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1872 5137 1900 5510
rect 1858 5128 1914 5137
rect 1858 5063 1914 5072
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1872 4321 1900 4422
rect 1858 4312 1914 4321
rect 1858 4247 1914 4256
rect 1858 3496 1914 3505
rect 1858 3431 1860 3440
rect 1912 3431 1914 3440
rect 1860 3402 1912 3408
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1872 2689 1900 2790
rect 1858 2680 1914 2689
rect 1858 2615 1914 2624
rect 1964 2514 1992 7142
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 2056 6322 2084 6666
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2148 2514 2176 7482
rect 2240 7154 2268 7942
rect 2516 7886 2544 8298
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2332 7342 2360 7686
rect 2424 7410 2452 7686
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2240 7126 2360 7154
rect 2226 6896 2282 6905
rect 2226 6831 2282 6840
rect 2240 6730 2268 6831
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2228 5568 2280 5574
rect 2226 5536 2228 5545
rect 2280 5536 2282 5545
rect 2226 5471 2282 5480
rect 2332 5114 2360 7126
rect 2504 6928 2556 6934
rect 2410 6896 2466 6905
rect 2504 6870 2556 6876
rect 2410 6831 2466 6840
rect 2240 5086 2360 5114
rect 2240 4826 2268 5086
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2240 4214 2268 4762
rect 2332 4729 2360 4966
rect 2318 4720 2374 4729
rect 2318 4655 2374 4664
rect 2228 4208 2280 4214
rect 2228 4150 2280 4156
rect 2320 3936 2372 3942
rect 2318 3904 2320 3913
rect 2372 3904 2374 3913
rect 2318 3839 2374 3848
rect 2424 3738 2452 6831
rect 2516 5794 2544 6870
rect 2608 5914 2636 9472
rect 2780 9454 2832 9460
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2700 8634 2728 8978
rect 2792 8945 2820 9454
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2700 7410 2728 8570
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2778 7304 2834 7313
rect 2778 7239 2834 7248
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2700 7002 2728 7142
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2700 6866 2728 6938
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2792 6730 2820 7239
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2688 5840 2740 5846
rect 2516 5788 2688 5794
rect 2516 5782 2740 5788
rect 2516 5766 2728 5782
rect 2792 5710 2820 5850
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2596 5296 2648 5302
rect 2594 5264 2596 5273
rect 2648 5264 2650 5273
rect 2594 5199 2650 5208
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2228 3120 2280 3126
rect 2226 3088 2228 3097
rect 2280 3088 2282 3097
rect 2226 3023 2282 3032
rect 2228 2916 2280 2922
rect 2228 2858 2280 2864
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2136 2508 2188 2514
rect 2136 2450 2188 2456
rect 2240 1306 2268 2858
rect 2792 2802 2820 5034
rect 2884 3176 2912 9574
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7546 3004 7890
rect 3068 7585 3096 9846
rect 3054 7576 3110 7585
rect 2964 7540 3016 7546
rect 3054 7511 3110 7520
rect 2964 7482 3016 7488
rect 3160 5778 3188 11206
rect 3436 11082 3464 12271
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3528 11354 3556 12106
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3698 11928 3754 11937
rect 3698 11863 3754 11872
rect 3712 11354 3740 11863
rect 3804 11694 3832 12038
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3528 11218 3556 11290
rect 3804 11286 3832 11630
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 4356 11150 4384 14311
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3252 10538 3280 11018
rect 3514 10976 3570 10985
rect 3514 10911 3570 10920
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 3252 9586 3280 10474
rect 3330 10024 3386 10033
rect 3330 9959 3386 9968
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3252 9178 3280 9522
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3344 8566 3372 9959
rect 3528 9926 3556 10911
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3606 9752 3662 9761
rect 3712 9722 3740 10066
rect 3804 9722 3832 10746
rect 4066 10568 4122 10577
rect 4066 10503 4068 10512
rect 4120 10503 4122 10512
rect 4068 10474 4120 10480
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4080 10169 4108 10202
rect 4066 10160 4122 10169
rect 4066 10095 4122 10104
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 3606 9687 3662 9696
rect 3700 9716 3752 9722
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9110 3464 9318
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3344 7970 3372 8502
rect 3436 8090 3464 8570
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3344 7954 3464 7970
rect 3344 7948 3476 7954
rect 3344 7942 3424 7948
rect 3424 7890 3476 7896
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3344 7002 3372 7142
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 6458 3280 6598
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3252 5846 3280 6122
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3160 5234 3188 5510
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2964 3188 3016 3194
rect 2884 3148 2964 3176
rect 2964 3130 3016 3136
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2148 1278 2268 1306
rect 2700 2774 2820 2802
rect 1766 1048 1822 1057
rect 1766 983 1822 992
rect 2148 800 2176 1278
rect 2700 800 2728 2774
rect 2884 2281 2912 2926
rect 2976 2854 3004 3130
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2964 2304 3016 2310
rect 2870 2272 2926 2281
rect 2964 2246 3016 2252
rect 2870 2207 2926 2216
rect 2976 1465 3004 2246
rect 2962 1456 3018 1465
rect 2962 1391 3018 1400
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1674 0 1730 800
rect 2134 0 2190 800
rect 2686 0 2742 800
rect 3068 241 3096 4082
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3160 800 3188 3130
rect 3054 232 3110 241
rect 3054 167 3110 176
rect 3146 0 3202 800
rect 3252 649 3280 4082
rect 3344 1873 3372 6666
rect 3436 5914 3464 7890
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3528 2582 3556 9590
rect 3620 9178 3648 9687
rect 3700 9658 3752 9664
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3698 9616 3754 9625
rect 3698 9551 3754 9560
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3712 9024 3740 9551
rect 3620 8996 3740 9024
rect 3620 6390 3648 8996
rect 3804 8634 3832 9658
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 3988 8945 4016 9318
rect 4172 9178 4200 9318
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4252 8968 4304 8974
rect 3974 8936 4030 8945
rect 4252 8910 4304 8916
rect 3974 8871 4030 8880
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3804 7886 3832 8298
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4172 6866 4200 7210
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3608 6248 3660 6254
rect 3712 6236 3740 6734
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 3660 6208 3740 6236
rect 3608 6190 3660 6196
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3804 5710 3832 6122
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3620 5370 3648 5646
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 3516 2576 3568 2582
rect 3516 2518 3568 2524
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3330 1864 3386 1873
rect 3330 1799 3386 1808
rect 3620 800 3648 2382
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 4264 1306 4292 8910
rect 4356 7002 4384 9862
rect 4448 8548 4476 13466
rect 4816 13462 4844 16400
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 5460 12918 5488 16400
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 5000 11694 5028 12174
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5000 11286 5028 11630
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10674 5764 10950
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 9518 4660 9862
rect 4816 9586 4844 10406
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4620 8560 4672 8566
rect 4448 8520 4620 8548
rect 4620 8502 4672 8508
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4448 7546 4476 7890
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4540 7410 4568 7686
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4632 7274 4660 8502
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4540 6118 4568 6802
rect 4724 6474 4752 9522
rect 4908 8378 4936 10474
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5092 10266 5120 10406
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5276 10062 5304 10610
rect 5920 10470 5948 11086
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5354 9888 5410 9897
rect 5354 9823 5410 9832
rect 5262 9752 5318 9761
rect 5262 9687 5318 9696
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5092 8974 5120 9454
rect 5276 9382 5304 9687
rect 5368 9586 5396 9823
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5460 9489 5488 9590
rect 5552 9500 5580 10134
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5644 9654 5672 10066
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5446 9480 5502 9489
rect 5552 9472 5672 9500
rect 5446 9415 5502 9424
rect 5644 9382 5672 9472
rect 5264 9376 5316 9382
rect 5540 9376 5592 9382
rect 5264 9318 5316 9324
rect 5354 9344 5410 9353
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 4988 8968 5040 8974
rect 4986 8936 4988 8945
rect 5080 8968 5132 8974
rect 5040 8936 5042 8945
rect 5080 8910 5132 8916
rect 4986 8871 5042 8880
rect 4816 8350 4936 8378
rect 4816 6610 4844 8350
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 7886 4936 8230
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4816 6582 4936 6610
rect 4724 6446 4844 6474
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4356 5098 4384 5306
rect 4540 5234 4568 6054
rect 4724 5710 4752 6258
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4540 4826 4568 4966
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4448 3754 4476 3946
rect 4540 3942 4568 4490
rect 4632 3942 4660 5646
rect 4724 5234 4752 5646
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4816 4690 4844 6446
rect 4908 5817 4936 6582
rect 4894 5808 4950 5817
rect 4894 5743 4950 5752
rect 5000 5658 5028 8871
rect 5184 7290 5212 9114
rect 5276 7800 5304 9318
rect 5540 9318 5592 9324
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5354 9279 5410 9288
rect 5368 9110 5396 9279
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5356 9104 5408 9110
rect 5460 9081 5488 9114
rect 5356 9046 5408 9052
rect 5446 9072 5502 9081
rect 5368 8634 5396 9046
rect 5446 9007 5502 9016
rect 5552 8906 5580 9318
rect 5540 8900 5592 8906
rect 5592 8860 5672 8888
rect 5540 8842 5592 8848
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5368 8362 5396 8570
rect 5644 8430 5672 8860
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5552 8090 5580 8230
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5644 7954 5672 8366
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5276 7772 5488 7800
rect 5184 7262 5304 7290
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 7002 5212 7142
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4908 5630 5028 5658
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4908 4622 4936 5630
rect 5092 5166 5120 5850
rect 5276 5386 5304 7262
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5368 6934 5396 7210
rect 5356 6928 5408 6934
rect 5354 6896 5356 6905
rect 5408 6896 5410 6905
rect 5460 6866 5488 7772
rect 5552 7546 5580 7890
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5644 7002 5672 7346
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5736 6882 5764 10202
rect 5920 10198 5948 10406
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5828 9654 5856 10066
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5920 9178 5948 9998
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5828 8809 5856 8978
rect 5908 8832 5960 8838
rect 5814 8800 5870 8809
rect 5908 8774 5960 8780
rect 5814 8735 5870 8744
rect 5920 8566 5948 8774
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 7342 5948 8230
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5354 6831 5410 6840
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5644 6854 5764 6882
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5368 5914 5396 6666
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5552 5846 5580 6598
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5184 5358 5304 5386
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5184 4826 5212 5358
rect 5264 5228 5316 5234
rect 5552 5216 5580 5782
rect 5316 5188 5580 5216
rect 5264 5170 5316 5176
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4448 3726 4660 3754
rect 4172 1278 4292 1306
rect 4172 800 4200 1278
rect 4632 800 4660 3726
rect 4908 2650 4936 4558
rect 5184 4486 5212 4762
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5184 4282 5212 4422
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5276 4078 5304 5170
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5368 4826 5396 5034
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5356 4616 5408 4622
rect 5460 4604 5488 5034
rect 5408 4576 5488 4604
rect 5356 4558 5408 4564
rect 5368 4282 5396 4558
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5276 3602 5304 4014
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5184 800 5212 3334
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5552 2582 5580 2858
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5276 2038 5304 2450
rect 5264 2032 5316 2038
rect 5264 1974 5316 1980
rect 5644 800 5672 6854
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5914 5764 6054
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5722 5808 5778 5817
rect 5722 5743 5778 5752
rect 5736 4146 5764 5743
rect 5828 5574 5856 7142
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5920 5273 5948 6122
rect 5906 5264 5962 5273
rect 5906 5199 5962 5208
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3126 5856 3878
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 6012 2666 6040 13942
rect 6104 13870 6132 16400
rect 6184 15292 6236 15298
rect 6184 15234 6236 15240
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 6104 8616 6132 11018
rect 6196 10810 6224 15234
rect 6552 15224 6604 15230
rect 6552 15166 6604 15172
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6196 10062 6224 10610
rect 6288 10266 6316 13806
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6380 11558 6408 12242
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 11150 6408 11494
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6288 9738 6316 10066
rect 6196 9710 6316 9738
rect 6196 8820 6224 9710
rect 6380 9586 6408 11086
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6472 9625 6500 10066
rect 6458 9616 6514 9625
rect 6368 9580 6420 9586
rect 6458 9551 6514 9560
rect 6368 9522 6420 9528
rect 6380 9110 6408 9522
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 9217 6500 9318
rect 6458 9208 6514 9217
rect 6458 9143 6514 9152
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6276 8968 6328 8974
rect 6328 8928 6408 8956
rect 6276 8910 6328 8916
rect 6196 8792 6316 8820
rect 6104 8588 6224 8616
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6104 8022 6132 8434
rect 6196 8090 6224 8588
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6092 8016 6144 8022
rect 6288 7970 6316 8792
rect 6380 8566 6408 8928
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6092 7958 6144 7964
rect 6104 7410 6132 7958
rect 6196 7942 6316 7970
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6104 4826 6132 6802
rect 6196 5817 6224 7942
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6182 5808 6238 5817
rect 6182 5743 6238 5752
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6104 4146 6132 4558
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6012 2638 6224 2666
rect 6196 800 6224 2638
rect 6288 2514 6316 7414
rect 6380 5778 6408 8502
rect 6472 7342 6500 9143
rect 6564 7954 6592 15166
rect 6748 14074 6776 16400
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 7392 13172 7420 16400
rect 7392 13144 7696 13172
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 6642 11656 6698 11665
rect 6642 11591 6698 11600
rect 6656 11218 6684 11591
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 7300 11286 7328 12038
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 6644 11212 6696 11218
rect 6696 11172 6776 11200
rect 6644 11154 6696 11160
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6656 10266 6684 10746
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6748 9704 6776 11172
rect 6840 11150 6868 11222
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6840 10606 6868 11086
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 7300 10130 7328 11222
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7392 10130 7420 10542
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 6748 9676 6868 9704
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6656 8974 6684 9522
rect 6734 9480 6790 9489
rect 6840 9466 6868 9676
rect 7116 9518 7144 9998
rect 7300 9586 7328 10066
rect 7484 10033 7512 10406
rect 7470 10024 7526 10033
rect 7470 9959 7526 9968
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7104 9512 7156 9518
rect 6918 9480 6974 9489
rect 6840 9438 6918 9466
rect 6734 9415 6790 9424
rect 7104 9454 7156 9460
rect 7286 9480 7342 9489
rect 6918 9415 6974 9424
rect 7286 9415 7342 9424
rect 6748 9382 6776 9415
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6734 9208 6790 9217
rect 6886 9200 7182 9220
rect 6734 9143 6736 9152
rect 6788 9143 6790 9152
rect 6736 9114 6788 9120
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6472 7002 6500 7278
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6472 6322 6500 6734
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6472 5302 6500 6258
rect 6564 6118 6592 7890
rect 6656 7410 6684 8910
rect 6748 8401 6776 8978
rect 7024 8809 7052 9046
rect 7010 8800 7066 8809
rect 7010 8735 7066 8744
rect 6734 8392 6790 8401
rect 6734 8327 6790 8336
rect 6748 8294 6776 8327
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6656 7206 6684 7346
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6748 6798 6776 7754
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6656 6186 6684 6394
rect 6840 6322 6868 6802
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7024 6458 7052 6666
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7116 4078 7144 4558
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 6656 3534 6684 4014
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 7300 3738 7328 9415
rect 7668 8498 7696 13144
rect 8036 12442 8064 16400
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7760 11898 7788 12378
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7760 11694 7788 11834
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8220 10606 8248 10950
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8312 10266 8340 10950
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7852 9897 7880 10066
rect 7838 9888 7894 9897
rect 7838 9823 7894 9832
rect 7838 9752 7894 9761
rect 7838 9687 7894 9696
rect 7852 9586 7880 9687
rect 8022 9616 8078 9625
rect 7840 9580 7892 9586
rect 8022 9551 8078 9560
rect 7840 9522 7892 9528
rect 8036 9518 8064 9551
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7392 5914 7420 8434
rect 8404 8430 8432 11698
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7656 8288 7708 8294
rect 7760 8265 7788 8366
rect 7656 8230 7708 8236
rect 7746 8256 7802 8265
rect 7576 8022 7604 8230
rect 7668 8090 7696 8230
rect 7746 8191 7802 8200
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 7342 7512 7686
rect 8036 7410 8064 7958
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 7546 8248 7822
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8220 7410 8248 7482
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7392 5166 7420 5714
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7484 3670 7512 4966
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6748 2514 6776 3062
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 7300 2514 7328 3538
rect 7484 2990 7512 3606
rect 7576 3194 7604 6258
rect 7944 4554 7972 6734
rect 8036 6458 8064 7142
rect 8128 7002 8156 7142
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8404 6934 8432 7210
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8496 6866 8524 14418
rect 8680 13734 8708 16400
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 9324 13530 9352 16400
rect 9968 14260 9996 16400
rect 9968 14232 10272 14260
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9416 11098 9444 13194
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 10244 12986 10272 14232
rect 10612 13190 10640 16400
rect 10968 15224 11020 15230
rect 10968 15166 11020 15172
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 9678 11792 9734 11801
rect 9678 11727 9734 11736
rect 9586 11656 9642 11665
rect 9692 11642 9720 11727
rect 9642 11614 9720 11642
rect 9586 11591 9642 11600
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 9416 11070 9628 11098
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8772 10130 8800 10678
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 8956 8906 8984 8978
rect 9140 8945 9168 8978
rect 9232 8974 9260 9522
rect 9416 8974 9444 9862
rect 9494 9072 9550 9081
rect 9494 9007 9550 9016
rect 9508 8974 9536 9007
rect 9220 8968 9272 8974
rect 9126 8936 9182 8945
rect 8944 8900 8996 8906
rect 9220 8910 9272 8916
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9126 8871 9182 8880
rect 8944 8842 8996 8848
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8588 8498 8616 8774
rect 8772 8566 8800 8774
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8588 7886 8616 8434
rect 8668 8424 8720 8430
rect 8666 8392 8668 8401
rect 8720 8392 8722 8401
rect 8864 8362 8892 8502
rect 9416 8498 9444 8910
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 8666 8327 8722 8336
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8668 8288 8720 8294
rect 8956 8265 8984 8298
rect 8668 8230 8720 8236
rect 8942 8256 8998 8265
rect 8680 8090 8708 8230
rect 8942 8191 8998 8200
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8680 7750 8708 8026
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8772 7342 8800 7822
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8496 6225 8524 6802
rect 8772 6798 8800 7278
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8588 6662 8616 6734
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8772 6322 8800 6734
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8956 6254 8984 6734
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6254 9536 6598
rect 8944 6248 8996 6254
rect 8482 6216 8538 6225
rect 8944 6190 8996 6196
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 8482 6151 8538 6160
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 8312 4282 8340 4626
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 8036 3738 8064 3946
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8128 3534 8156 3674
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8128 3194 8156 3470
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 6276 2508 6328 2514
rect 6276 2450 6328 2456
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6656 800 6684 2246
rect 7116 800 7144 2314
rect 7668 800 7696 2586
rect 7760 2514 7788 2790
rect 8404 2514 8432 3130
rect 8496 2650 8524 5646
rect 8588 4214 8616 5850
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8588 3738 8616 4150
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 9232 3602 9260 3946
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8588 2514 8616 3062
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8128 800 8156 2314
rect 8680 800 8708 3334
rect 8772 3058 8800 3402
rect 8864 3126 8892 3470
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 9600 3058 9628 11070
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 10138 10568 10194 10577
rect 10428 10538 10456 11154
rect 10138 10503 10194 10512
rect 10416 10532 10468 10538
rect 10152 10470 10180 10503
rect 10416 10474 10468 10480
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9784 9602 9812 9862
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 9784 9574 9904 9602
rect 10336 9586 10364 10406
rect 9876 9518 9904 9574
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 9110 9720 9318
rect 10244 9194 10272 9386
rect 10152 9166 10272 9194
rect 10152 9110 10180 9166
rect 9680 9104 9732 9110
rect 10140 9104 10192 9110
rect 9680 9046 9732 9052
rect 9954 9072 10010 9081
rect 10140 9046 10192 9052
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 9954 9007 9956 9016
rect 10008 9007 10010 9016
rect 9956 8978 10008 8984
rect 10244 8906 10272 9046
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9692 8566 9720 8774
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9784 8498 9812 8774
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 10230 8528 10286 8537
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 10048 8492 10100 8498
rect 10230 8463 10286 8472
rect 10048 8434 10100 8440
rect 9678 8392 9734 8401
rect 9678 8327 9734 8336
rect 9692 7750 9720 8327
rect 10060 7886 10088 8434
rect 10244 8430 10272 8463
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10244 8090 10272 8230
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 7206 9720 7278
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6390 9720 7142
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9692 5778 9720 6326
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9692 5030 9720 5714
rect 9784 5681 9812 7822
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9968 6730 9996 7414
rect 10244 7206 10272 7822
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 10336 5778 10364 9522
rect 10428 8906 10456 10474
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 10198 10548 10406
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 10598 9480 10654 9489
rect 10598 9415 10654 9424
rect 10612 9042 10640 9415
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10428 8294 10456 8434
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10428 7206 10456 7958
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10520 7002 10548 7278
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10612 6866 10640 6938
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10520 6390 10548 6734
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 9770 5672 9826 5681
rect 9770 5607 9826 5616
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9692 4622 9720 4966
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9692 3602 9720 4558
rect 9784 4554 9812 5034
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9784 4078 9812 4490
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9784 3482 9812 3878
rect 9876 3602 9904 4082
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10152 3738 10180 4014
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10152 3602 10180 3674
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 9692 3454 9812 3482
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8864 2650 8892 2858
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 9140 2514 9168 2790
rect 9692 2514 9720 3454
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 800 9168 2246
rect 9784 1034 9812 3334
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 9954 2952 10010 2961
rect 9954 2887 9956 2896
rect 10008 2887 10010 2896
rect 9956 2858 10008 2864
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 10244 1442 10272 3674
rect 10336 2961 10364 4762
rect 10612 4758 10640 4966
rect 10704 4826 10732 13670
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10796 10810 10824 12718
rect 10888 12646 10916 13942
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10796 10198 10824 10746
rect 10888 10266 10916 12582
rect 10980 12374 11008 15166
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10980 11370 11008 12310
rect 10980 11342 11100 11370
rect 11072 10538 11100 11342
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10980 9586 11008 10406
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10782 9072 10838 9081
rect 10782 9007 10784 9016
rect 10836 9007 10838 9016
rect 10784 8978 10836 8984
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8498 10824 8774
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 7274 10824 8230
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10888 7154 10916 8366
rect 11072 8362 11100 8570
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10980 7954 11008 8298
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10796 7126 10916 7154
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10600 4752 10652 4758
rect 10600 4694 10652 4700
rect 10612 4078 10640 4694
rect 10796 4214 10824 7126
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10888 6089 10916 6190
rect 10874 6080 10930 6089
rect 10874 6015 10930 6024
rect 10874 5536 10930 5545
rect 10874 5471 10930 5480
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10520 3924 10548 4014
rect 10796 3924 10824 4014
rect 10520 3896 10824 3924
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10322 2952 10378 2961
rect 10322 2887 10378 2896
rect 10428 2514 10456 3606
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10520 2446 10548 3896
rect 10598 3360 10654 3369
rect 10598 3295 10654 3304
rect 10612 3058 10640 3295
rect 10888 3097 10916 5471
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10980 3942 11008 5034
rect 11164 3942 11192 13466
rect 11256 13326 11284 16400
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11256 5234 11284 12718
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11348 10674 11376 11154
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11348 10062 11376 10610
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11532 9518 11560 10406
rect 11716 10266 11744 10474
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11610 9752 11666 9761
rect 11610 9687 11666 9696
rect 11624 9586 11652 9687
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11334 8528 11390 8537
rect 11334 8463 11390 8472
rect 11348 8430 11376 8463
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11532 7546 11560 8570
rect 11624 8090 11652 8978
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11624 7818 11652 8026
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11716 7750 11744 8978
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11532 5914 11560 7142
rect 11716 6118 11744 7686
rect 11808 7290 11836 14350
rect 11900 12782 11928 16400
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10606 11928 10950
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11900 10130 11928 10542
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11900 9586 11928 10066
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11886 7304 11942 7313
rect 11808 7262 11886 7290
rect 11808 6798 11836 7262
rect 11886 7239 11942 7248
rect 11992 6934 12020 7890
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11900 6390 11928 6598
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11900 6254 11928 6326
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11978 6080 12034 6089
rect 11978 6015 12034 6024
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11992 5710 12020 6015
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 11348 5370 11376 5510
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 12084 4826 12112 13262
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12176 10266 12204 10406
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 9518 12204 9862
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12164 7880 12216 7886
rect 12162 7848 12164 7857
rect 12216 7848 12218 7857
rect 12162 7783 12218 7792
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12176 7274 12204 7686
rect 12164 7268 12216 7274
rect 12164 7210 12216 7216
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6322 12204 6598
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11520 4208 11572 4214
rect 11440 4156 11520 4162
rect 11440 4150 11572 4156
rect 11440 4134 11560 4150
rect 11440 4078 11468 4134
rect 11624 4078 11652 4422
rect 12176 4078 12204 4762
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 11152 3936 11204 3942
rect 11204 3896 11284 3924
rect 11152 3878 11204 3884
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 10874 3088 10930 3097
rect 10600 3052 10652 3058
rect 10874 3023 10930 3032
rect 10600 2994 10652 3000
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 9692 1006 9812 1034
rect 10152 1414 10272 1442
rect 9692 800 9720 1006
rect 10152 800 10180 1414
rect 10612 800 10640 2246
rect 10796 2106 10824 2246
rect 10784 2100 10836 2106
rect 10784 2042 10836 2048
rect 11164 800 11192 3334
rect 11256 3058 11284 3896
rect 11624 3670 11652 4014
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11900 3602 11928 3946
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11888 3392 11940 3398
rect 11334 3360 11390 3369
rect 11992 3369 12020 3538
rect 11888 3334 11940 3340
rect 11978 3360 12034 3369
rect 11334 3295 11390 3304
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11348 2922 11376 3295
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11900 2582 11928 3334
rect 11978 3295 12034 3304
rect 12176 2922 12204 3674
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 12268 2582 12296 13330
rect 12452 12322 12480 14214
rect 12544 13394 12572 16400
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 13188 13462 13216 16400
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 13280 13172 13308 13874
rect 13832 13818 13860 16400
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 13832 13790 13952 13818
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13188 13144 13308 13172
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 12452 12294 12572 12322
rect 12438 10024 12494 10033
rect 12438 9959 12494 9968
rect 12452 9722 12480 9959
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 12360 7546 12388 7958
rect 12452 7886 12480 8774
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12360 6390 12388 7346
rect 12452 6934 12480 7822
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12360 5778 12388 6054
rect 12452 5914 12480 6054
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12360 5642 12388 5714
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12452 3194 12480 3538
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 11888 2576 11940 2582
rect 11888 2518 11940 2524
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 11612 2440 11664 2446
rect 12360 2394 12388 2926
rect 12440 2440 12492 2446
rect 11612 2382 11664 2388
rect 12176 2388 12440 2394
rect 12176 2382 12492 2388
rect 11624 800 11652 2382
rect 12176 2366 12480 2382
rect 12544 2378 12572 12294
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12636 10606 12664 11154
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9722 12664 9998
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12728 9024 12756 10610
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 13082 9480 13138 9489
rect 13082 9415 13084 9424
rect 13136 9415 13138 9424
rect 13084 9386 13136 9392
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 12728 8996 12848 9024
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12636 8090 12664 8502
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12728 8022 12756 8842
rect 12820 8401 12848 8996
rect 12806 8392 12862 8401
rect 12806 8327 12862 8336
rect 13188 8242 13216 13144
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13280 10674 13308 11154
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13280 10538 13308 10610
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13280 9722 13308 10066
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13280 9042 13308 9522
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13372 8634 13400 10406
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13188 8214 13308 8242
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12806 7440 12862 7449
rect 12912 7410 12940 7686
rect 13004 7410 13032 7822
rect 13188 7478 13216 7958
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 12806 7375 12862 7384
rect 12900 7404 12952 7410
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12728 6798 12756 7278
rect 12820 7274 12848 7375
rect 12900 7346 12952 7352
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12636 6361 12664 6734
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12622 6352 12678 6361
rect 12622 6287 12678 6296
rect 12636 4554 12664 6287
rect 12820 6254 12848 6598
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 13188 4690 13216 4966
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 13084 4140 13136 4146
rect 13280 4128 13308 8214
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 7002 13400 7142
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13358 6352 13414 6361
rect 13358 6287 13360 6296
rect 13412 6287 13414 6296
rect 13360 6258 13412 6264
rect 13360 5092 13412 5098
rect 13360 5034 13412 5040
rect 13372 4826 13400 5034
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13360 4140 13412 4146
rect 13136 4100 13216 4128
rect 13280 4100 13360 4128
rect 13084 4082 13136 4088
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12728 2582 12756 3334
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 12912 3097 12940 3130
rect 12898 3088 12954 3097
rect 12898 3023 12954 3032
rect 13004 2922 13032 3538
rect 13188 3466 13216 4100
rect 13360 4082 13412 4088
rect 13464 3738 13492 12922
rect 13832 12850 13860 13670
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13924 12442 13952 13790
rect 14200 13190 14228 14282
rect 14292 13938 14320 14282
rect 14476 13954 14504 16400
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14384 13926 14504 13954
rect 14384 13870 14412 13926
rect 15120 13870 15148 16400
rect 15290 15600 15346 15609
rect 15290 15535 15346 15544
rect 15198 14784 15254 14793
rect 15198 14719 15254 14728
rect 14372 13864 14424 13870
rect 14292 13812 14372 13818
rect 15108 13864 15160 13870
rect 14292 13806 14424 13812
rect 15028 13824 15108 13852
rect 14292 13790 14412 13806
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13556 10674 13584 11086
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13648 10742 13676 11018
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13556 10470 13584 10610
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13648 10062 13676 10678
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13556 9761 13584 9862
rect 13542 9752 13598 9761
rect 13542 9687 13598 9696
rect 13556 9518 13584 9687
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13648 9382 13676 9590
rect 13740 9586 13768 10406
rect 13832 10130 13860 10542
rect 13820 10124 13872 10130
rect 13872 10084 13952 10112
rect 13820 10066 13872 10072
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 9081 13768 9318
rect 13726 9072 13782 9081
rect 13726 9007 13782 9016
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 8498 13584 8910
rect 13832 8566 13860 9658
rect 13924 8838 13952 10084
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14016 8974 14044 9454
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13912 8832 13964 8838
rect 13964 8792 14044 8820
rect 13912 8774 13964 8780
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 14016 8498 14044 8792
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13556 7886 13584 8434
rect 13818 8392 13874 8401
rect 13818 8327 13874 8336
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13648 7732 13676 7890
rect 13740 7857 13768 7958
rect 13726 7848 13782 7857
rect 13726 7783 13782 7792
rect 13648 7704 13768 7732
rect 13740 7206 13768 7704
rect 13636 7200 13688 7206
rect 13634 7168 13636 7177
rect 13728 7200 13780 7206
rect 13688 7168 13690 7177
rect 13728 7142 13780 7148
rect 13634 7103 13690 7112
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13556 6458 13584 6938
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13832 5574 13860 8327
rect 13912 7336 13964 7342
rect 14016 7324 14044 8434
rect 13964 7296 14044 7324
rect 13912 7278 13964 7284
rect 14016 6798 14044 7296
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13912 6316 13964 6322
rect 14016 6304 14044 6734
rect 13964 6276 14044 6304
rect 13912 6258 13964 6264
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 14016 5914 14044 6122
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13176 3460 13228 3466
rect 13176 3402 13228 3408
rect 12992 2916 13044 2922
rect 12992 2858 13044 2864
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12532 2372 12584 2378
rect 12176 800 12204 2366
rect 12532 2314 12584 2320
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12636 800 12664 1702
rect 13188 800 13216 3402
rect 13556 1306 13584 4966
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14016 4214 14044 4626
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 14016 3942 14044 4150
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 14108 3602 14136 13126
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 2446 13676 3334
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 14004 2916 14056 2922
rect 14108 2904 14136 3538
rect 14056 2876 14136 2904
rect 14004 2858 14056 2864
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13648 1766 13676 2382
rect 13832 2310 13860 2858
rect 14200 2564 14228 13126
rect 14292 5234 14320 13790
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4010 14320 4422
rect 14384 4282 14412 13398
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14384 3738 14412 4082
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14292 2922 14320 3062
rect 14280 2916 14332 2922
rect 14280 2858 14332 2864
rect 14016 2536 14228 2564
rect 14016 2446 14044 2536
rect 14384 2496 14412 3674
rect 14108 2468 14412 2496
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13636 1760 13688 1766
rect 13636 1702 13688 1708
rect 13556 1278 13676 1306
rect 13648 800 13676 1278
rect 14108 800 14136 2468
rect 14476 2038 14504 9590
rect 14568 3602 14596 12378
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14660 8537 14688 11630
rect 14646 8528 14702 8537
rect 14646 8463 14702 8472
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14660 6934 14688 7278
rect 14648 6928 14700 6934
rect 14648 6870 14700 6876
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14568 2582 14596 2858
rect 14556 2576 14608 2582
rect 14556 2518 14608 2524
rect 14464 2032 14516 2038
rect 14464 1974 14516 1980
rect 14660 800 14688 4422
rect 14752 4010 14780 13330
rect 15028 12322 15056 13824
rect 15108 13806 15160 13812
rect 15212 12458 15240 14719
rect 15304 12617 15332 15535
rect 15764 14362 15792 16400
rect 16394 16400 16450 17200
rect 16486 16824 16542 16833
rect 16486 16759 16542 16768
rect 15842 16351 15898 16360
rect 15856 15230 15884 16351
rect 16210 16008 16266 16017
rect 16210 15943 16266 15952
rect 15844 15224 15896 15230
rect 15844 15166 15896 15172
rect 15672 14334 15792 14362
rect 15672 13938 15700 14334
rect 15782 14172 16078 14192
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15396 13530 15424 13670
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15488 12918 15516 13670
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15580 12730 15608 13806
rect 15672 13326 15700 13874
rect 15764 13841 15792 13942
rect 15750 13832 15806 13841
rect 15750 13767 15806 13776
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15658 12880 15714 12889
rect 15658 12815 15714 12824
rect 15396 12702 15608 12730
rect 15290 12608 15346 12617
rect 15290 12543 15346 12552
rect 15212 12430 15332 12458
rect 14844 12294 15056 12322
rect 14844 4146 14872 12294
rect 15198 12200 15254 12209
rect 15198 12135 15254 12144
rect 15212 11150 15240 12135
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15106 10704 15162 10713
rect 15106 10639 15162 10648
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14936 10266 14964 10542
rect 15016 10532 15068 10538
rect 15016 10474 15068 10480
rect 15028 10266 15056 10474
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14936 8838 14964 9998
rect 15028 9586 15056 10202
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15014 9480 15070 9489
rect 15014 9415 15016 9424
rect 15068 9415 15070 9424
rect 15016 9386 15068 9392
rect 15028 8945 15056 9386
rect 15014 8936 15070 8945
rect 15014 8871 15070 8880
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14936 7886 14964 8774
rect 15120 8090 15148 10639
rect 15198 10432 15254 10441
rect 15198 10367 15254 10376
rect 15212 9722 15240 10367
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15198 9480 15254 9489
rect 15198 9415 15254 9424
rect 15212 9382 15240 9415
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15120 7546 15148 7890
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15120 6798 15148 7482
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14936 6458 14964 6734
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 15212 5914 15240 8910
rect 15304 6118 15332 12430
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14752 3602 14780 3946
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14936 3534 14964 4558
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14844 3126 14872 3470
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 14832 3120 14884 3126
rect 14832 3062 14884 3068
rect 15212 2446 15240 3402
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15212 1714 15240 2382
rect 15396 2378 15424 12702
rect 15474 12336 15530 12345
rect 15474 12271 15530 12280
rect 15488 8090 15516 12271
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15580 10538 15608 11834
rect 15672 10792 15700 12815
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 16224 11898 16252 15943
rect 16302 14240 16358 14249
rect 16302 14175 16358 14184
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 15672 10764 15792 10792
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 8294 15608 10474
rect 15764 9908 15792 10764
rect 15672 9880 15792 9908
rect 15672 9704 15700 9880
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 15672 9676 15792 9704
rect 15764 8820 15792 9676
rect 16132 9568 16160 11018
rect 16316 11014 16344 14175
rect 16408 13870 16436 16400
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16210 10296 16266 10305
rect 16210 10231 16266 10240
rect 16224 10198 16252 10231
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 16224 9654 16252 10134
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 15672 8792 15792 8820
rect 16040 9540 16160 9568
rect 16040 8820 16068 9540
rect 16212 9512 16264 9518
rect 16118 9480 16174 9489
rect 16316 9500 16344 10406
rect 16264 9472 16344 9500
rect 16212 9454 16264 9460
rect 16118 9415 16174 9424
rect 16132 8888 16160 9415
rect 16132 8860 16252 8888
rect 16040 8792 16160 8820
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15566 8120 15622 8129
rect 15476 8084 15528 8090
rect 15566 8055 15622 8064
rect 15476 8026 15528 8032
rect 15488 7546 15516 8026
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15580 5234 15608 8055
rect 15672 7342 15700 8792
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 16132 7002 16160 8792
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 16132 6390 16160 6802
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15672 5681 15700 5850
rect 15764 5778 15792 6054
rect 15856 5914 15884 6190
rect 15936 6112 15988 6118
rect 16120 6112 16172 6118
rect 15988 6072 16120 6100
rect 15936 6054 15988 6060
rect 16120 6054 16172 6060
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15658 5672 15714 5681
rect 15658 5607 15714 5616
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 16132 5302 16160 6054
rect 16224 5642 16252 8860
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16316 7954 16344 8774
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 16224 5370 16252 5578
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 16408 4758 16436 13262
rect 16500 9625 16528 16759
rect 17038 16400 17094 17200
rect 17682 16400 17738 17200
rect 18326 16400 18382 17200
rect 18970 16400 19026 17200
rect 19614 16400 19670 17200
rect 17052 13258 17080 16400
rect 17406 13424 17462 13433
rect 17696 13394 17724 16400
rect 17774 15192 17830 15201
rect 17774 15127 17830 15136
rect 17406 13359 17462 13368
rect 17684 13388 17736 13394
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16592 11257 16620 12106
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 16578 11248 16634 11257
rect 16578 11183 16634 11192
rect 16762 11248 16818 11257
rect 16762 11183 16818 11192
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16592 10305 16620 10610
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16578 10296 16634 10305
rect 16578 10231 16580 10240
rect 16632 10231 16634 10240
rect 16580 10202 16632 10208
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16486 9616 16542 9625
rect 16592 9586 16620 10066
rect 16684 9994 16712 10406
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16486 9551 16542 9560
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16592 9466 16620 9522
rect 16488 9444 16540 9450
rect 16592 9438 16712 9466
rect 16488 9386 16540 9392
rect 16500 9110 16528 9386
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16500 8498 16528 8842
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16592 7818 16620 9318
rect 16684 8634 16712 9438
rect 16776 9024 16804 11183
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16960 10266 16988 10406
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16868 10033 16896 10066
rect 16854 10024 16910 10033
rect 16854 9959 16910 9968
rect 17130 10024 17186 10033
rect 17130 9959 17186 9968
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16868 9217 16896 9862
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 16960 9466 16988 9590
rect 16960 9438 17080 9466
rect 16854 9208 16910 9217
rect 16854 9143 16910 9152
rect 16776 8996 16896 9024
rect 16762 8936 16818 8945
rect 16762 8871 16818 8880
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16776 8498 16804 8871
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16684 8090 16712 8298
rect 16776 8090 16804 8434
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16500 7002 16528 7482
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16684 6730 16712 7210
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 16684 6322 16712 6666
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16500 5710 16528 6258
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16500 4758 16528 5170
rect 16592 4826 16620 6054
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16684 5370 16712 5714
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16868 4842 16896 8996
rect 17052 8378 17080 9438
rect 17144 9042 17172 9959
rect 17328 9568 17356 11290
rect 17420 10577 17448 13359
rect 17684 13330 17736 13336
rect 17788 11082 17816 15127
rect 18340 14278 18368 16400
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18984 13190 19012 16400
rect 19628 14346 19656 16400
rect 19616 14340 19668 14346
rect 19616 14282 19668 14288
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18142 11792 18198 11801
rect 18142 11727 18198 11736
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17406 10568 17462 10577
rect 17406 10503 17462 10512
rect 17776 10532 17828 10538
rect 17420 10266 17448 10503
rect 17776 10474 17828 10480
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 10266 17540 10406
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17420 9722 17448 10202
rect 17788 10198 17816 10474
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17328 9540 17540 9568
rect 17512 9450 17540 9540
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17500 9444 17552 9450
rect 17500 9386 17552 9392
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17236 8786 17264 9318
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17144 8758 17264 8786
rect 17144 8566 17172 8758
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17144 8430 17172 8502
rect 16960 8350 17080 8378
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 16960 5234 16988 8350
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 17052 8022 17080 8230
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17236 7886 17264 8570
rect 17328 8498 17356 8910
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17420 7562 17448 9386
rect 17604 9178 17632 9454
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17512 8974 17540 9046
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17512 7954 17540 8910
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17604 8090 17632 8366
rect 17696 8265 17724 9590
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 9217 17816 9318
rect 17774 9208 17830 9217
rect 17880 9178 17908 9386
rect 17972 9330 18000 10066
rect 18064 9518 18092 10746
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17972 9302 18092 9330
rect 17774 9143 17830 9152
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17682 8256 17738 8265
rect 17682 8191 17738 8200
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17420 7534 17540 7562
rect 17040 7472 17092 7478
rect 17040 7414 17092 7420
rect 17052 6866 17080 7414
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17236 6934 17264 7278
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17328 6798 17356 7346
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17328 6390 17356 6734
rect 17316 6384 17368 6390
rect 17316 6326 17368 6332
rect 17420 6322 17448 6802
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17512 5914 17540 7534
rect 17604 7342 17632 7686
rect 17880 7449 17908 8502
rect 17972 8362 18000 8774
rect 18064 8430 18092 9302
rect 18156 9110 18184 11727
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17866 7440 17922 7449
rect 17866 7375 17922 7384
rect 17972 7342 18000 8298
rect 18156 7857 18184 8434
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18142 7848 18198 7857
rect 18142 7783 18198 7792
rect 18248 7478 18276 7890
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 17592 7336 17644 7342
rect 17590 7304 17592 7313
rect 17960 7336 18012 7342
rect 17644 7304 17646 7313
rect 17960 7278 18012 7284
rect 17590 7239 17646 7248
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 18142 7168 18198 7177
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17132 5704 17184 5710
rect 17130 5672 17132 5681
rect 17224 5704 17276 5710
rect 17184 5672 17186 5681
rect 17224 5646 17276 5652
rect 17130 5607 17186 5616
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16960 5030 16988 5170
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16776 4826 16988 4842
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16776 4820 17000 4826
rect 16776 4814 16948 4820
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 15488 3602 15516 4694
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16132 3670 16160 3878
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16316 3602 16344 4082
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16408 3670 16436 3946
rect 16396 3664 16448 3670
rect 16396 3606 16448 3612
rect 16776 3602 16804 4814
rect 16948 4762 17000 4768
rect 16856 4752 16908 4758
rect 16856 4694 16908 4700
rect 16868 3738 16896 4694
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 15120 1686 15240 1714
rect 15120 800 15148 1686
rect 15580 898 15608 2790
rect 15672 2582 15700 3334
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 15764 2582 15792 2858
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 15752 2576 15804 2582
rect 15752 2518 15804 2524
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 15580 870 15700 898
rect 15672 800 15700 870
rect 16132 800 16160 3062
rect 16224 2922 16252 3538
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16224 2106 16252 2858
rect 17144 2582 17172 5607
rect 17236 5234 17264 5646
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17236 4622 17264 5170
rect 17512 5166 17540 5850
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17420 4690 17448 5102
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17236 3602 17264 4082
rect 17512 4078 17540 4966
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 16684 800 16712 2246
rect 17144 800 17172 2246
rect 17420 1306 17448 3334
rect 17512 2990 17540 3674
rect 17604 3398 17632 7142
rect 17788 6633 17816 7142
rect 17774 6624 17830 6633
rect 17774 6559 17830 6568
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17682 5808 17738 5817
rect 17682 5743 17684 5752
rect 17736 5743 17738 5752
rect 17684 5714 17736 5720
rect 17788 5234 17816 6394
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17880 5114 17908 7142
rect 18142 7103 18198 7112
rect 18052 6248 18104 6254
rect 18050 6216 18052 6225
rect 18104 6216 18106 6225
rect 18050 6151 18106 6160
rect 18050 5672 18106 5681
rect 18156 5642 18184 7103
rect 18234 6216 18290 6225
rect 18234 6151 18290 6160
rect 18248 6118 18276 6151
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18050 5607 18052 5616
rect 18104 5607 18106 5616
rect 18144 5636 18196 5642
rect 18052 5578 18104 5584
rect 18144 5578 18196 5584
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17696 5086 17908 5114
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17604 2514 17632 3334
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 17592 2304 17644 2310
rect 17590 2272 17592 2281
rect 17644 2272 17646 2281
rect 17590 2207 17646 2216
rect 17420 1278 17632 1306
rect 17604 800 17632 1278
rect 3238 640 3294 649
rect 3238 575 3294 584
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5170 0 5226 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11610 0 11666 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13634 0 13690 800
rect 14094 0 14150 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17130 0 17186 800
rect 17590 0 17646 800
rect 17696 649 17724 5086
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 4865 17816 4966
rect 17774 4856 17830 4865
rect 17774 4791 17830 4800
rect 17972 4690 18000 5510
rect 18340 5273 18368 10406
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18602 8800 18658 8809
rect 18602 8735 18658 8744
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18432 7002 18460 7278
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18326 5264 18382 5273
rect 18326 5199 18382 5208
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17788 3602 17816 3878
rect 17880 3641 17908 4422
rect 17866 3632 17922 3641
rect 17776 3596 17828 3602
rect 17866 3567 17922 3576
rect 17776 3538 17828 3544
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 3233 18092 3334
rect 18050 3224 18106 3233
rect 18050 3159 18106 3168
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17788 2689 17816 2790
rect 17774 2680 17830 2689
rect 17774 2615 17830 2624
rect 17880 2394 17908 2790
rect 17788 2366 17908 2394
rect 17788 1873 17816 2366
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17774 1864 17830 1873
rect 17774 1799 17830 1808
rect 17880 1057 17908 2246
rect 17866 1048 17922 1057
rect 17866 983 17922 992
rect 18156 800 18184 4490
rect 18248 4457 18276 4966
rect 18432 4690 18460 5510
rect 18420 4684 18472 4690
rect 18420 4626 18472 4632
rect 18420 4480 18472 4486
rect 18234 4448 18290 4457
rect 18420 4422 18472 4428
rect 18234 4383 18290 4392
rect 18432 4049 18460 4422
rect 18418 4040 18474 4049
rect 18418 3975 18474 3984
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 17682 640 17738 649
rect 17682 575 17738 584
rect 18142 0 18198 800
rect 18248 241 18276 3878
rect 18524 1465 18552 7754
rect 18616 6458 18644 8735
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18708 4010 18736 9114
rect 18972 7064 19024 7070
rect 18970 7032 18972 7041
rect 19024 7032 19026 7041
rect 18970 6967 19026 6976
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18510 1456 18566 1465
rect 18510 1391 18566 1400
rect 18616 800 18644 3334
rect 19168 800 19196 3402
rect 19616 3120 19668 3126
rect 19616 3062 19668 3068
rect 19628 800 19656 3062
rect 18234 232 18290 241
rect 18234 167 18290 176
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19614 0 19670 800
<< via2 >>
rect 2778 16360 2834 16416
rect 3330 16768 3386 16824
rect 3054 15952 3110 16008
rect 2870 13912 2926 13968
rect 1582 11328 1638 11384
rect 1858 8064 1914 8120
rect 2962 12688 3018 12744
rect 3238 15544 3294 15600
rect 3330 15136 3386 15192
rect 3330 13524 3386 13560
rect 3330 13504 3332 13524
rect 3332 13504 3384 13524
rect 3384 13504 3386 13524
rect 3330 13096 3386 13152
rect 4066 14728 4122 14784
rect 4342 14320 4398 14376
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3422 12280 3478 12336
rect 2226 8472 2282 8528
rect 1858 7692 1860 7712
rect 1860 7692 1912 7712
rect 1912 7692 1914 7712
rect 1858 7656 1914 7692
rect 1858 6432 1914 6488
rect 1858 6060 1860 6080
rect 1860 6060 1912 6080
rect 1912 6060 1914 6080
rect 1858 6024 1914 6060
rect 1858 5072 1914 5128
rect 1858 4256 1914 4312
rect 1858 3460 1914 3496
rect 1858 3440 1860 3460
rect 1860 3440 1912 3460
rect 1912 3440 1914 3460
rect 1858 2624 1914 2680
rect 2226 6840 2282 6896
rect 2226 5516 2228 5536
rect 2228 5516 2280 5536
rect 2280 5516 2282 5536
rect 2226 5480 2282 5516
rect 2410 6840 2466 6896
rect 2318 4664 2374 4720
rect 2318 3884 2320 3904
rect 2320 3884 2372 3904
rect 2372 3884 2374 3904
rect 2318 3848 2374 3884
rect 2778 8880 2834 8936
rect 2778 7248 2834 7304
rect 2594 5244 2596 5264
rect 2596 5244 2648 5264
rect 2648 5244 2650 5264
rect 2594 5208 2650 5244
rect 2226 3068 2228 3088
rect 2228 3068 2280 3088
rect 2280 3068 2282 3088
rect 2226 3032 2282 3068
rect 3054 7520 3110 7576
rect 3698 11872 3754 11928
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3514 10920 3570 10976
rect 3330 9968 3386 10024
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 3606 9696 3662 9752
rect 4066 10532 4122 10568
rect 4066 10512 4068 10532
rect 4068 10512 4120 10532
rect 4120 10512 4122 10532
rect 4066 10104 4122 10160
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 1766 992 1822 1048
rect 2870 2216 2926 2272
rect 2962 1400 3018 1456
rect 3054 176 3110 232
rect 3698 9560 3754 9616
rect 3974 8880 4030 8936
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 3330 1808 3386 1864
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 5354 9832 5410 9888
rect 5262 9696 5318 9752
rect 5446 9424 5502 9480
rect 4986 8916 4988 8936
rect 4988 8916 5040 8936
rect 5040 8916 5042 8936
rect 4986 8880 5042 8916
rect 4894 5752 4950 5808
rect 5354 9288 5410 9344
rect 5446 9016 5502 9072
rect 5354 6876 5356 6896
rect 5356 6876 5408 6896
rect 5408 6876 5410 6896
rect 5354 6840 5410 6876
rect 5814 8744 5870 8800
rect 5722 5752 5778 5808
rect 5906 5208 5962 5264
rect 6458 9560 6514 9616
rect 6458 9152 6514 9208
rect 6182 5752 6238 5808
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6642 11600 6698 11656
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 6734 9424 6790 9480
rect 7470 9968 7526 10024
rect 6918 9424 6974 9480
rect 7286 9424 7342 9480
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 6734 9172 6790 9208
rect 6734 9152 6736 9172
rect 6736 9152 6788 9172
rect 6788 9152 6790 9172
rect 7010 8744 7066 8800
rect 6734 8336 6790 8392
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 7838 9832 7894 9888
rect 7838 9696 7894 9752
rect 8022 9560 8078 9616
rect 7746 8200 7802 8256
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9678 11736 9734 11792
rect 9586 11600 9642 11656
rect 9494 9016 9550 9072
rect 9126 8880 9182 8936
rect 8666 8372 8668 8392
rect 8668 8372 8720 8392
rect 8720 8372 8722 8392
rect 8666 8336 8722 8372
rect 8942 8200 8998 8256
rect 8482 6160 8538 6216
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 10138 10512 10194 10568
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9954 9036 10010 9072
rect 9954 9016 9956 9036
rect 9956 9016 10008 9036
rect 10008 9016 10010 9036
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10230 8472 10286 8528
rect 9678 8336 9734 8392
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 10598 9424 10654 9480
rect 9770 5616 9826 5672
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 9954 2916 10010 2952
rect 9954 2896 9956 2916
rect 9956 2896 10008 2916
rect 10008 2896 10010 2916
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 10782 9036 10838 9072
rect 10782 9016 10784 9036
rect 10784 9016 10836 9036
rect 10836 9016 10838 9036
rect 10874 6024 10930 6080
rect 10874 5480 10930 5536
rect 10322 2896 10378 2952
rect 10598 3304 10654 3360
rect 11610 9696 11666 9752
rect 11334 8472 11390 8528
rect 11886 7248 11942 7304
rect 11978 6024 12034 6080
rect 12162 7828 12164 7848
rect 12164 7828 12216 7848
rect 12216 7828 12218 7848
rect 12162 7792 12218 7828
rect 10874 3032 10930 3088
rect 11334 3304 11390 3360
rect 11978 3304 12034 3360
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12438 9968 12494 10024
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 13082 9444 13138 9480
rect 13082 9424 13084 9444
rect 13084 9424 13136 9444
rect 13136 9424 13138 9444
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 12806 8336 12862 8392
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 12806 7384 12862 7440
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 12622 6296 12678 6352
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 13358 6316 13414 6352
rect 13358 6296 13360 6316
rect 13360 6296 13412 6316
rect 13412 6296 13414 6316
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 12898 3032 12954 3088
rect 15290 15544 15346 15600
rect 15198 14728 15254 14784
rect 13542 9696 13598 9752
rect 13726 9016 13782 9072
rect 13818 8336 13874 8392
rect 13726 7792 13782 7848
rect 13634 7148 13636 7168
rect 13636 7148 13688 7168
rect 13688 7148 13690 7168
rect 13634 7112 13690 7148
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 14646 8472 14702 8528
rect 15842 16360 15898 16416
rect 16486 16768 16542 16824
rect 16210 15952 16266 16008
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 15750 13776 15806 13832
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15658 12824 15714 12880
rect 15290 12552 15346 12608
rect 15198 12144 15254 12200
rect 15106 10648 15162 10704
rect 15014 9444 15070 9480
rect 15014 9424 15016 9444
rect 15016 9424 15068 9444
rect 15068 9424 15070 9444
rect 15014 8880 15070 8936
rect 15198 10376 15254 10432
rect 15198 9424 15254 9480
rect 15474 12280 15530 12336
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 16302 14184 16358 14240
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 16210 10240 16266 10296
rect 16118 9424 16174 9480
rect 15566 8064 15622 8120
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15658 5616 15714 5672
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 17406 13368 17462 13424
rect 17774 15136 17830 15192
rect 16578 11192 16634 11248
rect 16762 11192 16818 11248
rect 16578 10260 16634 10296
rect 16578 10240 16580 10260
rect 16580 10240 16632 10260
rect 16632 10240 16634 10260
rect 16486 9560 16542 9616
rect 16854 9968 16910 10024
rect 17130 9968 17186 10024
rect 16854 9152 16910 9208
rect 16762 8880 16818 8936
rect 18142 11736 18198 11792
rect 17406 10512 17462 10568
rect 17774 9152 17830 9208
rect 17682 8200 17738 8256
rect 17866 7384 17922 7440
rect 18142 7792 18198 7848
rect 17590 7284 17592 7304
rect 17592 7284 17644 7304
rect 17644 7284 17646 7304
rect 17590 7248 17646 7284
rect 17130 5652 17132 5672
rect 17132 5652 17184 5672
rect 17184 5652 17186 5672
rect 17130 5616 17186 5652
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 17774 6568 17830 6624
rect 17682 5772 17738 5808
rect 17682 5752 17684 5772
rect 17684 5752 17736 5772
rect 17736 5752 17738 5772
rect 18142 7112 18198 7168
rect 18050 6196 18052 6216
rect 18052 6196 18104 6216
rect 18104 6196 18106 6216
rect 18050 6160 18106 6196
rect 18050 5636 18106 5672
rect 18234 6160 18290 6216
rect 18050 5616 18052 5636
rect 18052 5616 18104 5636
rect 18104 5616 18106 5636
rect 17590 2252 17592 2272
rect 17592 2252 17644 2272
rect 17644 2252 17646 2272
rect 17590 2216 17646 2252
rect 3238 584 3294 640
rect 17774 4800 17830 4856
rect 18602 8744 18658 8800
rect 18326 5208 18382 5264
rect 17866 3576 17922 3632
rect 18050 3168 18106 3224
rect 17774 2624 17830 2680
rect 17774 1808 17830 1864
rect 17866 992 17922 1048
rect 18234 4392 18290 4448
rect 18418 3984 18474 4040
rect 17682 584 17738 640
rect 18970 7012 18972 7032
rect 18972 7012 19024 7032
rect 19024 7012 19026 7032
rect 18970 6976 19026 7012
rect 18510 1400 18566 1456
rect 18234 176 18290 232
<< metal3 >>
rect 0 16826 800 16856
rect 3325 16826 3391 16829
rect 0 16824 3391 16826
rect 0 16768 3330 16824
rect 3386 16768 3391 16824
rect 0 16766 3391 16768
rect 0 16736 800 16766
rect 3325 16763 3391 16766
rect 16481 16826 16547 16829
rect 19200 16826 20000 16856
rect 16481 16824 20000 16826
rect 16481 16768 16486 16824
rect 16542 16768 20000 16824
rect 16481 16766 20000 16768
rect 16481 16763 16547 16766
rect 19200 16736 20000 16766
rect 0 16418 800 16448
rect 2773 16418 2839 16421
rect 0 16416 2839 16418
rect 0 16360 2778 16416
rect 2834 16360 2839 16416
rect 0 16358 2839 16360
rect 0 16328 800 16358
rect 2773 16355 2839 16358
rect 15837 16418 15903 16421
rect 19200 16418 20000 16448
rect 15837 16416 20000 16418
rect 15837 16360 15842 16416
rect 15898 16360 20000 16416
rect 15837 16358 20000 16360
rect 15837 16355 15903 16358
rect 19200 16328 20000 16358
rect 0 16010 800 16040
rect 3049 16010 3115 16013
rect 0 16008 3115 16010
rect 0 15952 3054 16008
rect 3110 15952 3115 16008
rect 0 15950 3115 15952
rect 0 15920 800 15950
rect 3049 15947 3115 15950
rect 16205 16010 16271 16013
rect 19200 16010 20000 16040
rect 16205 16008 20000 16010
rect 16205 15952 16210 16008
rect 16266 15952 20000 16008
rect 16205 15950 20000 15952
rect 16205 15947 16271 15950
rect 19200 15920 20000 15950
rect 0 15602 800 15632
rect 3233 15602 3299 15605
rect 0 15600 3299 15602
rect 0 15544 3238 15600
rect 3294 15544 3299 15600
rect 0 15542 3299 15544
rect 0 15512 800 15542
rect 3233 15539 3299 15542
rect 15285 15602 15351 15605
rect 19200 15602 20000 15632
rect 15285 15600 20000 15602
rect 15285 15544 15290 15600
rect 15346 15544 20000 15600
rect 15285 15542 20000 15544
rect 15285 15539 15351 15542
rect 19200 15512 20000 15542
rect 0 15194 800 15224
rect 3325 15194 3391 15197
rect 0 15192 3391 15194
rect 0 15136 3330 15192
rect 3386 15136 3391 15192
rect 0 15134 3391 15136
rect 0 15104 800 15134
rect 3325 15131 3391 15134
rect 17769 15194 17835 15197
rect 19200 15194 20000 15224
rect 17769 15192 20000 15194
rect 17769 15136 17774 15192
rect 17830 15136 20000 15192
rect 17769 15134 20000 15136
rect 17769 15131 17835 15134
rect 19200 15104 20000 15134
rect 0 14786 800 14816
rect 4061 14786 4127 14789
rect 0 14784 4127 14786
rect 0 14728 4066 14784
rect 4122 14728 4127 14784
rect 0 14726 4127 14728
rect 0 14696 800 14726
rect 4061 14723 4127 14726
rect 15193 14786 15259 14789
rect 19200 14786 20000 14816
rect 15193 14784 20000 14786
rect 15193 14728 15198 14784
rect 15254 14728 20000 14784
rect 15193 14726 20000 14728
rect 15193 14723 15259 14726
rect 6874 14720 7194 14721
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 19200 14696 20000 14726
rect 12805 14655 13125 14656
rect 0 14378 800 14408
rect 4337 14378 4403 14381
rect 0 14376 4403 14378
rect 0 14320 4342 14376
rect 4398 14320 4403 14376
rect 0 14318 4403 14320
rect 0 14288 800 14318
rect 4337 14315 4403 14318
rect 16297 14242 16363 14245
rect 19200 14242 20000 14272
rect 16297 14240 20000 14242
rect 16297 14184 16302 14240
rect 16358 14184 20000 14240
rect 16297 14182 20000 14184
rect 16297 14179 16363 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19200 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13970 800 14000
rect 2865 13970 2931 13973
rect 0 13968 2931 13970
rect 0 13912 2870 13968
rect 2926 13912 2931 13968
rect 0 13910 2931 13912
rect 0 13880 800 13910
rect 2865 13907 2931 13910
rect 15745 13834 15811 13837
rect 19200 13834 20000 13864
rect 15745 13832 20000 13834
rect 15745 13776 15750 13832
rect 15806 13776 20000 13832
rect 15745 13774 20000 13776
rect 15745 13771 15811 13774
rect 19200 13744 20000 13774
rect 6874 13632 7194 13633
rect 0 13562 800 13592
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 3325 13562 3391 13565
rect 0 13560 3391 13562
rect 0 13504 3330 13560
rect 3386 13504 3391 13560
rect 0 13502 3391 13504
rect 0 13472 800 13502
rect 3325 13499 3391 13502
rect 17401 13426 17467 13429
rect 19200 13426 20000 13456
rect 17401 13424 20000 13426
rect 17401 13368 17406 13424
rect 17462 13368 20000 13424
rect 17401 13366 20000 13368
rect 17401 13363 17467 13366
rect 19200 13336 20000 13366
rect 0 13154 800 13184
rect 3325 13154 3391 13157
rect 0 13152 3391 13154
rect 0 13096 3330 13152
rect 3386 13096 3391 13152
rect 0 13094 3391 13096
rect 0 13064 800 13094
rect 3325 13091 3391 13094
rect 3909 13088 4229 13089
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 19200 13018 20000 13048
rect 16208 12958 20000 13018
rect 15653 12882 15719 12885
rect 16208 12882 16268 12958
rect 19200 12928 20000 12958
rect 15653 12880 16268 12882
rect 15653 12824 15658 12880
rect 15714 12824 16268 12880
rect 15653 12822 16268 12824
rect 15653 12819 15719 12822
rect 0 12746 800 12776
rect 2957 12746 3023 12749
rect 0 12744 3023 12746
rect 0 12688 2962 12744
rect 3018 12688 3023 12744
rect 0 12686 3023 12688
rect 0 12656 800 12686
rect 2957 12683 3023 12686
rect 15285 12610 15351 12613
rect 15510 12610 15516 12612
rect 15285 12608 15516 12610
rect 15285 12552 15290 12608
rect 15346 12552 15516 12608
rect 15285 12550 15516 12552
rect 15285 12547 15351 12550
rect 15510 12548 15516 12550
rect 15580 12548 15586 12612
rect 16246 12548 16252 12612
rect 16316 12610 16322 12612
rect 19200 12610 20000 12640
rect 16316 12550 20000 12610
rect 16316 12548 16322 12550
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 19200 12520 20000 12550
rect 12805 12479 13125 12480
rect 0 12338 800 12368
rect 3417 12338 3483 12341
rect 15469 12340 15535 12341
rect 15469 12338 15516 12340
rect 0 12336 3483 12338
rect 0 12280 3422 12336
rect 3478 12280 3483 12336
rect 0 12278 3483 12280
rect 15424 12336 15516 12338
rect 15424 12280 15474 12336
rect 15424 12278 15516 12280
rect 0 12248 800 12278
rect 3417 12275 3483 12278
rect 15469 12276 15516 12278
rect 15580 12276 15586 12340
rect 15469 12275 15535 12276
rect 15193 12202 15259 12205
rect 19200 12202 20000 12232
rect 15193 12200 20000 12202
rect 15193 12144 15198 12200
rect 15254 12144 20000 12200
rect 15193 12142 20000 12144
rect 15193 12139 15259 12142
rect 19200 12112 20000 12142
rect 3909 12000 4229 12001
rect 0 11930 800 11960
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 3693 11930 3759 11933
rect 0 11928 3759 11930
rect 0 11872 3698 11928
rect 3754 11872 3759 11928
rect 0 11870 3759 11872
rect 0 11840 800 11870
rect 3693 11867 3759 11870
rect 9673 11794 9739 11797
rect 18137 11794 18203 11797
rect 19200 11794 20000 11824
rect 9673 11792 20000 11794
rect 9673 11736 9678 11792
rect 9734 11736 18142 11792
rect 18198 11736 20000 11792
rect 9673 11734 20000 11736
rect 9673 11731 9739 11734
rect 18137 11731 18203 11734
rect 19200 11704 20000 11734
rect 6637 11658 6703 11661
rect 9581 11658 9647 11661
rect 6637 11656 9647 11658
rect 6637 11600 6642 11656
rect 6698 11600 9586 11656
rect 9642 11600 9647 11656
rect 6637 11598 9647 11600
rect 6637 11595 6703 11598
rect 9581 11595 9647 11598
rect 6874 11456 7194 11457
rect 0 11386 800 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 1577 11386 1643 11389
rect 0 11384 1643 11386
rect 0 11328 1582 11384
rect 1638 11328 1643 11384
rect 0 11326 1643 11328
rect 0 11296 800 11326
rect 1577 11323 1643 11326
rect 16573 11250 16639 11253
rect 16757 11250 16823 11253
rect 19200 11250 20000 11280
rect 16573 11248 20000 11250
rect 16573 11192 16578 11248
rect 16634 11192 16762 11248
rect 16818 11192 20000 11248
rect 16573 11190 20000 11192
rect 16573 11187 16639 11190
rect 16757 11187 16823 11190
rect 19200 11160 20000 11190
rect 0 10978 800 11008
rect 3509 10978 3575 10981
rect 0 10976 3575 10978
rect 0 10920 3514 10976
rect 3570 10920 3575 10976
rect 0 10918 3575 10920
rect 0 10888 800 10918
rect 3509 10915 3575 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 19200 10842 20000 10872
rect 16254 10782 20000 10842
rect 15101 10706 15167 10709
rect 16254 10706 16314 10782
rect 19200 10752 20000 10782
rect 15101 10704 16314 10706
rect 15101 10648 15106 10704
rect 15162 10648 16314 10704
rect 15101 10646 16314 10648
rect 15101 10643 15167 10646
rect 0 10570 800 10600
rect 4061 10570 4127 10573
rect 0 10568 4127 10570
rect 0 10512 4066 10568
rect 4122 10512 4127 10568
rect 0 10510 4127 10512
rect 0 10480 800 10510
rect 4061 10507 4127 10510
rect 10133 10570 10199 10573
rect 17401 10570 17467 10573
rect 10133 10568 17467 10570
rect 10133 10512 10138 10568
rect 10194 10512 17406 10568
rect 17462 10512 17467 10568
rect 10133 10510 17467 10512
rect 10133 10507 10199 10510
rect 17401 10507 17467 10510
rect 15193 10434 15259 10437
rect 19200 10434 20000 10464
rect 15193 10432 20000 10434
rect 15193 10376 15198 10432
rect 15254 10376 20000 10432
rect 15193 10374 20000 10376
rect 15193 10371 15259 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19200 10344 20000 10374
rect 12805 10303 13125 10304
rect 16205 10298 16271 10301
rect 16573 10298 16639 10301
rect 16205 10296 16639 10298
rect 16205 10240 16210 10296
rect 16266 10240 16578 10296
rect 16634 10240 16639 10296
rect 16205 10238 16639 10240
rect 16205 10235 16271 10238
rect 16573 10235 16639 10238
rect 0 10162 800 10192
rect 4061 10162 4127 10165
rect 0 10160 4127 10162
rect 0 10104 4066 10160
rect 4122 10104 4127 10160
rect 0 10102 4127 10104
rect 0 10072 800 10102
rect 4061 10099 4127 10102
rect 3325 10026 3391 10029
rect 7465 10026 7531 10029
rect 3325 10024 7531 10026
rect 3325 9968 3330 10024
rect 3386 9968 7470 10024
rect 7526 9968 7531 10024
rect 3325 9966 7531 9968
rect 3325 9963 3391 9966
rect 7465 9963 7531 9966
rect 12433 10026 12499 10029
rect 16849 10026 16915 10029
rect 12433 10024 16915 10026
rect 12433 9968 12438 10024
rect 12494 9968 16854 10024
rect 16910 9968 16915 10024
rect 12433 9966 16915 9968
rect 12433 9963 12499 9966
rect 16849 9963 16915 9966
rect 17125 10026 17191 10029
rect 19200 10026 20000 10056
rect 17125 10024 20000 10026
rect 17125 9968 17130 10024
rect 17186 9968 20000 10024
rect 17125 9966 20000 9968
rect 17125 9963 17191 9966
rect 19200 9936 20000 9966
rect 5349 9890 5415 9893
rect 7833 9890 7899 9893
rect 5349 9888 7899 9890
rect 5349 9832 5354 9888
rect 5410 9832 7838 9888
rect 7894 9832 7899 9888
rect 5349 9830 7899 9832
rect 5349 9827 5415 9830
rect 7833 9827 7899 9830
rect 3909 9824 4229 9825
rect 0 9754 800 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 9759 16090 9760
rect 3601 9754 3667 9757
rect 0 9752 3667 9754
rect 0 9696 3606 9752
rect 3662 9696 3667 9752
rect 0 9694 3667 9696
rect 0 9664 800 9694
rect 3601 9691 3667 9694
rect 5257 9754 5323 9757
rect 7833 9754 7899 9757
rect 5257 9752 7899 9754
rect 5257 9696 5262 9752
rect 5318 9696 7838 9752
rect 7894 9696 7899 9752
rect 5257 9694 7899 9696
rect 5257 9691 5323 9694
rect 7833 9691 7899 9694
rect 11605 9754 11671 9757
rect 13537 9754 13603 9757
rect 11605 9752 13603 9754
rect 11605 9696 11610 9752
rect 11666 9696 13542 9752
rect 13598 9696 13603 9752
rect 11605 9694 13603 9696
rect 11605 9691 11671 9694
rect 13537 9691 13603 9694
rect 3693 9618 3759 9621
rect 6453 9618 6519 9621
rect 3693 9616 6519 9618
rect 3693 9560 3698 9616
rect 3754 9560 6458 9616
rect 6514 9560 6519 9616
rect 3693 9558 6519 9560
rect 3693 9555 3759 9558
rect 6453 9555 6519 9558
rect 8017 9618 8083 9621
rect 16481 9618 16547 9621
rect 19200 9618 20000 9648
rect 8017 9616 16547 9618
rect 8017 9560 8022 9616
rect 8078 9560 16486 9616
rect 16542 9560 16547 9616
rect 8017 9558 16547 9560
rect 8017 9555 8083 9558
rect 16481 9555 16547 9558
rect 16622 9558 20000 9618
rect 5441 9482 5507 9485
rect 6729 9482 6795 9485
rect 5441 9480 6795 9482
rect 5441 9424 5446 9480
rect 5502 9424 6734 9480
rect 6790 9424 6795 9480
rect 5441 9422 6795 9424
rect 5441 9419 5507 9422
rect 6729 9419 6795 9422
rect 6913 9482 6979 9485
rect 7281 9482 7347 9485
rect 6913 9480 7347 9482
rect 6913 9424 6918 9480
rect 6974 9424 7286 9480
rect 7342 9424 7347 9480
rect 6913 9422 7347 9424
rect 6913 9419 6979 9422
rect 7281 9419 7347 9422
rect 10593 9482 10659 9485
rect 13077 9482 13143 9485
rect 15009 9482 15075 9485
rect 10593 9480 15075 9482
rect 10593 9424 10598 9480
rect 10654 9424 13082 9480
rect 13138 9424 15014 9480
rect 15070 9424 15075 9480
rect 10593 9422 15075 9424
rect 10593 9419 10659 9422
rect 13077 9419 13143 9422
rect 15009 9419 15075 9422
rect 15193 9482 15259 9485
rect 16113 9482 16179 9485
rect 16622 9482 16682 9558
rect 19200 9528 20000 9558
rect 15193 9480 16682 9482
rect 15193 9424 15198 9480
rect 15254 9424 16118 9480
rect 16174 9424 16682 9480
rect 15193 9422 16682 9424
rect 15193 9419 15259 9422
rect 16113 9419 16179 9422
rect 0 9346 800 9376
rect 5349 9346 5415 9349
rect 0 9344 5415 9346
rect 0 9288 5354 9344
rect 5410 9288 5415 9344
rect 0 9286 5415 9288
rect 0 9256 800 9286
rect 5349 9283 5415 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 6453 9210 6519 9213
rect 6729 9210 6795 9213
rect 16849 9210 16915 9213
rect 6453 9208 6795 9210
rect 6453 9152 6458 9208
rect 6514 9152 6734 9208
rect 6790 9152 6795 9208
rect 6453 9150 6795 9152
rect 6453 9147 6519 9150
rect 6729 9147 6795 9150
rect 16806 9208 16915 9210
rect 16806 9152 16854 9208
rect 16910 9152 16915 9208
rect 16806 9147 16915 9152
rect 17769 9210 17835 9213
rect 19200 9210 20000 9240
rect 17769 9208 20000 9210
rect 17769 9152 17774 9208
rect 17830 9152 20000 9208
rect 17769 9150 20000 9152
rect 17769 9147 17835 9150
rect 5441 9074 5507 9077
rect 9489 9074 9555 9077
rect 5441 9072 9555 9074
rect 5441 9016 5446 9072
rect 5502 9016 9494 9072
rect 9550 9016 9555 9072
rect 5441 9014 9555 9016
rect 5441 9011 5507 9014
rect 9489 9011 9555 9014
rect 9949 9074 10015 9077
rect 10777 9074 10843 9077
rect 13721 9074 13787 9077
rect 9949 9072 13787 9074
rect 9949 9016 9954 9072
rect 10010 9016 10782 9072
rect 10838 9016 13726 9072
rect 13782 9016 13787 9072
rect 9949 9014 13787 9016
rect 9949 9011 10015 9014
rect 10777 9011 10843 9014
rect 13721 9011 13787 9014
rect 0 8938 800 8968
rect 16806 8941 16866 9147
rect 19200 9120 20000 9150
rect 2773 8938 2839 8941
rect 0 8936 2839 8938
rect 0 8880 2778 8936
rect 2834 8880 2839 8936
rect 0 8878 2839 8880
rect 0 8848 800 8878
rect 2773 8875 2839 8878
rect 3969 8938 4035 8941
rect 4981 8938 5047 8941
rect 9121 8938 9187 8941
rect 3969 8936 9187 8938
rect 3969 8880 3974 8936
rect 4030 8880 4986 8936
rect 5042 8880 9126 8936
rect 9182 8880 9187 8936
rect 3969 8878 9187 8880
rect 3969 8875 4035 8878
rect 4981 8875 5047 8878
rect 9121 8875 9187 8878
rect 15009 8938 15075 8941
rect 15009 8936 16314 8938
rect 15009 8880 15014 8936
rect 15070 8880 16314 8936
rect 15009 8878 16314 8880
rect 15009 8875 15075 8878
rect 5809 8802 5875 8805
rect 7005 8802 7071 8805
rect 5809 8800 7071 8802
rect 5809 8744 5814 8800
rect 5870 8744 7010 8800
rect 7066 8744 7071 8800
rect 5809 8742 7071 8744
rect 16254 8802 16314 8878
rect 16757 8936 16866 8941
rect 16757 8880 16762 8936
rect 16818 8880 16866 8936
rect 16757 8878 16866 8880
rect 16757 8875 16823 8878
rect 18597 8802 18663 8805
rect 19200 8802 20000 8832
rect 16254 8800 20000 8802
rect 16254 8744 18602 8800
rect 18658 8744 20000 8800
rect 16254 8742 20000 8744
rect 5809 8739 5875 8742
rect 7005 8739 7071 8742
rect 18597 8739 18663 8742
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 19200 8712 20000 8742
rect 15770 8671 16090 8672
rect 0 8530 800 8560
rect 2221 8530 2287 8533
rect 0 8528 2287 8530
rect 0 8472 2226 8528
rect 2282 8472 2287 8528
rect 0 8470 2287 8472
rect 0 8440 800 8470
rect 2221 8467 2287 8470
rect 10225 8530 10291 8533
rect 11329 8530 11395 8533
rect 10225 8528 11395 8530
rect 10225 8472 10230 8528
rect 10286 8472 11334 8528
rect 11390 8472 11395 8528
rect 10225 8470 11395 8472
rect 10225 8467 10291 8470
rect 11329 8467 11395 8470
rect 14641 8530 14707 8533
rect 14641 8528 15348 8530
rect 14641 8472 14646 8528
rect 14702 8472 15348 8528
rect 14641 8470 15348 8472
rect 14641 8467 14707 8470
rect 6729 8394 6795 8397
rect 8661 8394 8727 8397
rect 6729 8392 8727 8394
rect 6729 8336 6734 8392
rect 6790 8336 8666 8392
rect 8722 8336 8727 8392
rect 6729 8334 8727 8336
rect 6729 8331 6795 8334
rect 8661 8331 8727 8334
rect 9673 8394 9739 8397
rect 12801 8394 12867 8397
rect 13813 8394 13879 8397
rect 9673 8392 13879 8394
rect 9673 8336 9678 8392
rect 9734 8336 12806 8392
rect 12862 8336 13818 8392
rect 13874 8336 13879 8392
rect 9673 8334 13879 8336
rect 9673 8331 9739 8334
rect 12801 8331 12867 8334
rect 13813 8331 13879 8334
rect 7741 8258 7807 8261
rect 8937 8258 9003 8261
rect 7741 8256 9003 8258
rect 7741 8200 7746 8256
rect 7802 8200 8942 8256
rect 8998 8200 9003 8256
rect 7741 8198 9003 8200
rect 7741 8195 7807 8198
rect 8937 8195 9003 8198
rect 6874 8192 7194 8193
rect 0 8122 800 8152
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 8127 13125 8128
rect 1853 8122 1919 8125
rect 0 8120 1919 8122
rect 0 8064 1858 8120
rect 1914 8064 1919 8120
rect 0 8062 1919 8064
rect 15288 8122 15348 8470
rect 17677 8258 17743 8261
rect 19200 8258 20000 8288
rect 17677 8256 20000 8258
rect 17677 8200 17682 8256
rect 17738 8200 20000 8256
rect 17677 8198 20000 8200
rect 17677 8195 17743 8198
rect 19200 8168 20000 8198
rect 15561 8122 15627 8125
rect 15288 8120 15627 8122
rect 15288 8064 15566 8120
rect 15622 8064 15627 8120
rect 15288 8062 15627 8064
rect 0 8032 800 8062
rect 1853 8059 1919 8062
rect 15561 8059 15627 8062
rect 12157 7850 12223 7853
rect 13721 7850 13787 7853
rect 12157 7848 13787 7850
rect 12157 7792 12162 7848
rect 12218 7792 13726 7848
rect 13782 7792 13787 7848
rect 12157 7790 13787 7792
rect 12157 7787 12223 7790
rect 13721 7787 13787 7790
rect 18137 7850 18203 7853
rect 19200 7850 20000 7880
rect 18137 7848 20000 7850
rect 18137 7792 18142 7848
rect 18198 7792 20000 7848
rect 18137 7790 20000 7792
rect 18137 7787 18203 7790
rect 19200 7760 20000 7790
rect 0 7714 800 7744
rect 1853 7714 1919 7717
rect 0 7712 1919 7714
rect 0 7656 1858 7712
rect 1914 7656 1919 7712
rect 0 7654 1919 7656
rect 0 7624 800 7654
rect 1853 7651 1919 7654
rect 3909 7648 4229 7649
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 3049 7578 3115 7581
rect 3049 7576 3250 7578
rect 3049 7520 3054 7576
rect 3110 7520 3250 7576
rect 3049 7518 3250 7520
rect 3049 7515 3115 7518
rect 3190 7442 3250 7518
rect 12801 7442 12867 7445
rect 3190 7440 12867 7442
rect 3190 7384 12806 7440
rect 12862 7384 12867 7440
rect 3190 7382 12867 7384
rect 12801 7379 12867 7382
rect 17861 7442 17927 7445
rect 19200 7442 20000 7472
rect 17861 7440 20000 7442
rect 17861 7384 17866 7440
rect 17922 7384 20000 7440
rect 17861 7382 20000 7384
rect 17861 7379 17927 7382
rect 19200 7352 20000 7382
rect 0 7306 800 7336
rect 2773 7306 2839 7309
rect 0 7304 2839 7306
rect 0 7248 2778 7304
rect 2834 7248 2839 7304
rect 0 7246 2839 7248
rect 0 7216 800 7246
rect 2773 7243 2839 7246
rect 11881 7306 11947 7309
rect 17585 7306 17651 7309
rect 11881 7304 17651 7306
rect 11881 7248 11886 7304
rect 11942 7248 17590 7304
rect 17646 7248 17651 7304
rect 11881 7246 17651 7248
rect 11881 7243 11947 7246
rect 17585 7243 17651 7246
rect 13629 7170 13695 7173
rect 18137 7170 18203 7173
rect 13629 7168 18203 7170
rect 13629 7112 13634 7168
rect 13690 7112 18142 7168
rect 18198 7112 18203 7168
rect 13629 7110 18203 7112
rect 13629 7107 13695 7110
rect 18137 7107 18203 7110
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 18965 7034 19031 7037
rect 19200 7034 20000 7064
rect 18965 7032 20000 7034
rect 18965 6976 18970 7032
rect 19026 6976 20000 7032
rect 18965 6974 20000 6976
rect 18965 6971 19031 6974
rect 19200 6944 20000 6974
rect 0 6898 800 6928
rect 2221 6898 2287 6901
rect 0 6896 2287 6898
rect 0 6840 2226 6896
rect 2282 6840 2287 6896
rect 0 6838 2287 6840
rect 0 6808 800 6838
rect 2221 6835 2287 6838
rect 2405 6898 2471 6901
rect 5349 6898 5415 6901
rect 2405 6896 5415 6898
rect 2405 6840 2410 6896
rect 2466 6840 5354 6896
rect 5410 6840 5415 6896
rect 2405 6838 5415 6840
rect 2405 6835 2471 6838
rect 5349 6835 5415 6838
rect 17769 6626 17835 6629
rect 19200 6626 20000 6656
rect 17769 6624 20000 6626
rect 17769 6568 17774 6624
rect 17830 6568 20000 6624
rect 17769 6566 20000 6568
rect 17769 6563 17835 6566
rect 3909 6560 4229 6561
rect 0 6490 800 6520
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 19200 6536 20000 6566
rect 15770 6495 16090 6496
rect 1853 6490 1919 6493
rect 0 6488 1919 6490
rect 0 6432 1858 6488
rect 1914 6432 1919 6488
rect 0 6430 1919 6432
rect 0 6400 800 6430
rect 1853 6427 1919 6430
rect 12617 6354 12683 6357
rect 13353 6354 13419 6357
rect 16246 6354 16252 6356
rect 12617 6352 16252 6354
rect 12617 6296 12622 6352
rect 12678 6296 13358 6352
rect 13414 6296 16252 6352
rect 12617 6294 16252 6296
rect 12617 6291 12683 6294
rect 13353 6291 13419 6294
rect 16246 6292 16252 6294
rect 16316 6292 16322 6356
rect 8477 6218 8543 6221
rect 18045 6218 18111 6221
rect 8477 6216 18111 6218
rect 8477 6160 8482 6216
rect 8538 6160 18050 6216
rect 18106 6160 18111 6216
rect 8477 6158 18111 6160
rect 8477 6155 8543 6158
rect 18045 6155 18111 6158
rect 18229 6218 18295 6221
rect 19200 6218 20000 6248
rect 18229 6216 20000 6218
rect 18229 6160 18234 6216
rect 18290 6160 20000 6216
rect 18229 6158 20000 6160
rect 18229 6155 18295 6158
rect 19200 6128 20000 6158
rect 0 6082 800 6112
rect 1853 6082 1919 6085
rect 0 6080 1919 6082
rect 0 6024 1858 6080
rect 1914 6024 1919 6080
rect 0 6022 1919 6024
rect 0 5992 800 6022
rect 1853 6019 1919 6022
rect 10869 6082 10935 6085
rect 11973 6082 12039 6085
rect 10869 6080 12039 6082
rect 10869 6024 10874 6080
rect 10930 6024 11978 6080
rect 12034 6024 12039 6080
rect 10869 6022 12039 6024
rect 10869 6019 10935 6022
rect 11973 6019 12039 6022
rect 6874 6016 7194 6017
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 5951 13125 5952
rect 4889 5810 4955 5813
rect 5717 5810 5783 5813
rect 4889 5808 5783 5810
rect 4889 5752 4894 5808
rect 4950 5752 5722 5808
rect 5778 5752 5783 5808
rect 4889 5750 5783 5752
rect 4889 5747 4955 5750
rect 5717 5747 5783 5750
rect 6177 5810 6243 5813
rect 17677 5810 17743 5813
rect 6177 5808 17743 5810
rect 6177 5752 6182 5808
rect 6238 5752 17682 5808
rect 17738 5752 17743 5808
rect 6177 5750 17743 5752
rect 6177 5747 6243 5750
rect 17677 5747 17743 5750
rect 5720 5674 5780 5747
rect 9765 5674 9831 5677
rect 15653 5674 15719 5677
rect 17125 5674 17191 5677
rect 5720 5672 10794 5674
rect 5720 5616 9770 5672
rect 9826 5616 10794 5672
rect 5720 5614 10794 5616
rect 9765 5611 9831 5614
rect 0 5538 800 5568
rect 2221 5538 2287 5541
rect 0 5536 2287 5538
rect 0 5480 2226 5536
rect 2282 5480 2287 5536
rect 0 5478 2287 5480
rect 10734 5538 10794 5614
rect 15653 5672 17191 5674
rect 15653 5616 15658 5672
rect 15714 5616 17130 5672
rect 17186 5616 17191 5672
rect 15653 5614 17191 5616
rect 15653 5611 15719 5614
rect 17125 5611 17191 5614
rect 18045 5674 18111 5677
rect 19200 5674 20000 5704
rect 18045 5672 20000 5674
rect 18045 5616 18050 5672
rect 18106 5616 20000 5672
rect 18045 5614 20000 5616
rect 18045 5611 18111 5614
rect 19200 5584 20000 5614
rect 10869 5538 10935 5541
rect 10734 5536 10935 5538
rect 10734 5480 10874 5536
rect 10930 5480 10935 5536
rect 10734 5478 10935 5480
rect 0 5448 800 5478
rect 2221 5475 2287 5478
rect 10869 5475 10935 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 2589 5266 2655 5269
rect 5901 5266 5967 5269
rect 2589 5264 5967 5266
rect 2589 5208 2594 5264
rect 2650 5208 5906 5264
rect 5962 5208 5967 5264
rect 2589 5206 5967 5208
rect 2589 5203 2655 5206
rect 5901 5203 5967 5206
rect 18321 5266 18387 5269
rect 19200 5266 20000 5296
rect 18321 5264 20000 5266
rect 18321 5208 18326 5264
rect 18382 5208 20000 5264
rect 18321 5206 20000 5208
rect 18321 5203 18387 5206
rect 19200 5176 20000 5206
rect 0 5130 800 5160
rect 1853 5130 1919 5133
rect 0 5128 1919 5130
rect 0 5072 1858 5128
rect 1914 5072 1919 5128
rect 0 5070 1919 5072
rect 0 5040 800 5070
rect 1853 5067 1919 5070
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 17769 4858 17835 4861
rect 19200 4858 20000 4888
rect 17769 4856 20000 4858
rect 17769 4800 17774 4856
rect 17830 4800 20000 4856
rect 17769 4798 20000 4800
rect 17769 4795 17835 4798
rect 19200 4768 20000 4798
rect 0 4722 800 4752
rect 2313 4722 2379 4725
rect 0 4720 2379 4722
rect 0 4664 2318 4720
rect 2374 4664 2379 4720
rect 0 4662 2379 4664
rect 0 4632 800 4662
rect 2313 4659 2379 4662
rect 18229 4450 18295 4453
rect 19200 4450 20000 4480
rect 18229 4448 20000 4450
rect 18229 4392 18234 4448
rect 18290 4392 20000 4448
rect 18229 4390 20000 4392
rect 18229 4387 18295 4390
rect 3909 4384 4229 4385
rect 0 4314 800 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19200 4360 20000 4390
rect 15770 4319 16090 4320
rect 1853 4314 1919 4317
rect 0 4312 1919 4314
rect 0 4256 1858 4312
rect 1914 4256 1919 4312
rect 0 4254 1919 4256
rect 0 4224 800 4254
rect 1853 4251 1919 4254
rect 18413 4042 18479 4045
rect 19200 4042 20000 4072
rect 18413 4040 20000 4042
rect 18413 3984 18418 4040
rect 18474 3984 20000 4040
rect 18413 3982 20000 3984
rect 18413 3979 18479 3982
rect 19200 3952 20000 3982
rect 0 3906 800 3936
rect 2313 3906 2379 3909
rect 0 3904 2379 3906
rect 0 3848 2318 3904
rect 2374 3848 2379 3904
rect 0 3846 2379 3848
rect 0 3816 800 3846
rect 2313 3843 2379 3846
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 17861 3634 17927 3637
rect 19200 3634 20000 3664
rect 17861 3632 20000 3634
rect 17861 3576 17866 3632
rect 17922 3576 20000 3632
rect 17861 3574 20000 3576
rect 17861 3571 17927 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 800 3438
rect 1853 3435 1919 3438
rect 10593 3362 10659 3365
rect 11329 3362 11395 3365
rect 11973 3362 12039 3365
rect 10593 3360 12039 3362
rect 10593 3304 10598 3360
rect 10654 3304 11334 3360
rect 11390 3304 11978 3360
rect 12034 3304 12039 3360
rect 10593 3302 12039 3304
rect 10593 3299 10659 3302
rect 11329 3299 11395 3302
rect 11973 3299 12039 3302
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 18045 3226 18111 3229
rect 19200 3226 20000 3256
rect 18045 3224 20000 3226
rect 18045 3168 18050 3224
rect 18106 3168 20000 3224
rect 18045 3166 20000 3168
rect 18045 3163 18111 3166
rect 19200 3136 20000 3166
rect 0 3090 800 3120
rect 2221 3090 2287 3093
rect 0 3088 2287 3090
rect 0 3032 2226 3088
rect 2282 3032 2287 3088
rect 0 3030 2287 3032
rect 0 3000 800 3030
rect 2221 3027 2287 3030
rect 10869 3090 10935 3093
rect 12893 3090 12959 3093
rect 10869 3088 12959 3090
rect 10869 3032 10874 3088
rect 10930 3032 12898 3088
rect 12954 3032 12959 3088
rect 10869 3030 12959 3032
rect 10869 3027 10935 3030
rect 12893 3027 12959 3030
rect 9949 2954 10015 2957
rect 10317 2954 10383 2957
rect 9949 2952 10383 2954
rect 9949 2896 9954 2952
rect 10010 2896 10322 2952
rect 10378 2896 10383 2952
rect 9949 2894 10383 2896
rect 9949 2891 10015 2894
rect 10317 2891 10383 2894
rect 6874 2752 7194 2753
rect 0 2682 800 2712
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2687 13125 2688
rect 1853 2682 1919 2685
rect 0 2680 1919 2682
rect 0 2624 1858 2680
rect 1914 2624 1919 2680
rect 0 2622 1919 2624
rect 0 2592 800 2622
rect 1853 2619 1919 2622
rect 17769 2682 17835 2685
rect 19200 2682 20000 2712
rect 17769 2680 20000 2682
rect 17769 2624 17774 2680
rect 17830 2624 20000 2680
rect 17769 2622 20000 2624
rect 17769 2619 17835 2622
rect 19200 2592 20000 2622
rect 0 2274 800 2304
rect 2865 2274 2931 2277
rect 0 2272 2931 2274
rect 0 2216 2870 2272
rect 2926 2216 2931 2272
rect 0 2214 2931 2216
rect 0 2184 800 2214
rect 2865 2211 2931 2214
rect 17585 2274 17651 2277
rect 19200 2274 20000 2304
rect 17585 2272 20000 2274
rect 17585 2216 17590 2272
rect 17646 2216 20000 2272
rect 17585 2214 20000 2216
rect 17585 2211 17651 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 19200 2184 20000 2214
rect 15770 2143 16090 2144
rect 0 1866 800 1896
rect 3325 1866 3391 1869
rect 0 1864 3391 1866
rect 0 1808 3330 1864
rect 3386 1808 3391 1864
rect 0 1806 3391 1808
rect 0 1776 800 1806
rect 3325 1803 3391 1806
rect 17769 1866 17835 1869
rect 19200 1866 20000 1896
rect 17769 1864 20000 1866
rect 17769 1808 17774 1864
rect 17830 1808 20000 1864
rect 17769 1806 20000 1808
rect 17769 1803 17835 1806
rect 19200 1776 20000 1806
rect 0 1458 800 1488
rect 2957 1458 3023 1461
rect 0 1456 3023 1458
rect 0 1400 2962 1456
rect 3018 1400 3023 1456
rect 0 1398 3023 1400
rect 0 1368 800 1398
rect 2957 1395 3023 1398
rect 18505 1458 18571 1461
rect 19200 1458 20000 1488
rect 18505 1456 20000 1458
rect 18505 1400 18510 1456
rect 18566 1400 20000 1456
rect 18505 1398 20000 1400
rect 18505 1395 18571 1398
rect 19200 1368 20000 1398
rect 0 1050 800 1080
rect 1761 1050 1827 1053
rect 0 1048 1827 1050
rect 0 992 1766 1048
rect 1822 992 1827 1048
rect 0 990 1827 992
rect 0 960 800 990
rect 1761 987 1827 990
rect 17861 1050 17927 1053
rect 19200 1050 20000 1080
rect 17861 1048 20000 1050
rect 17861 992 17866 1048
rect 17922 992 20000 1048
rect 17861 990 20000 992
rect 17861 987 17927 990
rect 19200 960 20000 990
rect 0 642 800 672
rect 3233 642 3299 645
rect 0 640 3299 642
rect 0 584 3238 640
rect 3294 584 3299 640
rect 0 582 3299 584
rect 0 552 800 582
rect 3233 579 3299 582
rect 17677 642 17743 645
rect 19200 642 20000 672
rect 17677 640 20000 642
rect 17677 584 17682 640
rect 17738 584 20000 640
rect 17677 582 20000 584
rect 17677 579 17743 582
rect 19200 552 20000 582
rect 0 234 800 264
rect 3049 234 3115 237
rect 0 232 3115 234
rect 0 176 3054 232
rect 3110 176 3115 232
rect 0 174 3115 176
rect 0 144 800 174
rect 3049 171 3115 174
rect 18229 234 18295 237
rect 19200 234 20000 264
rect 18229 232 20000 234
rect 18229 176 18234 232
rect 18290 176 20000 232
rect 18229 174 20000 176
rect 18229 171 18295 174
rect 19200 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 15516 12548 15580 12612
rect 16252 12548 16316 12612
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 15516 12336 15580 12340
rect 15516 12280 15530 12336
rect 15530 12280 15580 12336
rect 15516 12276 15580 12280
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 16252 6292 16316 6356
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 15770 14176 16091 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16091 14176
rect 15770 13088 16091 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16091 13088
rect 15515 12612 15581 12613
rect 15515 12548 15516 12612
rect 15580 12548 15581 12612
rect 15515 12547 15581 12548
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 15518 12341 15578 12547
rect 15515 12340 15581 12341
rect 15515 12276 15516 12340
rect 15580 12276 15581 12340
rect 15515 12275 15581 12276
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 15770 12000 16091 13024
rect 16251 12612 16317 12613
rect 16251 12548 16252 12612
rect 16316 12548 16317 12612
rect 16251 12547 16317 12548
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16091 12000
rect 15770 10912 16091 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16091 10912
rect 15770 9824 16091 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16091 9824
rect 15770 8736 16091 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16091 8736
rect 15770 7648 16091 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16091 7648
rect 15770 6560 16091 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16091 6560
rect 15770 5472 16091 6496
rect 16254 6357 16314 12547
rect 16251 6356 16317 6357
rect 16251 6292 16252 6356
rect 16316 6292 16317 6356
rect 16251 6291 16317 6292
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16091 5472
rect 15770 4384 16091 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16091 4384
rect 15770 3296 16091 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16091 3296
rect 15770 2208 16091 3232
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16091 2208
rect 15770 2128 16091 2144
use sky130_fd_sc_hd__decap_3  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1564 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _18_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1656 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2116 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1608910539
transform 1 0 2024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2668 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1608910539
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1608910539
transform 1 0 2392 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1608910539
transform 1 0 2760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_34 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4232 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_22
timestamp 1608910539
transform 1 0 3128 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4600 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30
timestamp 1608910539
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1608910539
transform 1 0 3128 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 3312 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_62
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1608910539
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_46
timestamp 1608910539
transform 1 0 5336 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5888 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 5336 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608910539
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 6900 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608910539
transform 1 0 7084 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608910539
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_81
timestamp 1608910539
transform 1 0 8556 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1608910539
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608910539
transform 1 0 8464 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608910539
transform 1 0 8096 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8648 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1608910539
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87
timestamp 1608910539
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608910539
transform 1 0 10304 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 9844 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8832 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608910539
transform 1 0 9936 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608910539
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1608910539
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 12604 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 11040 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608910539
transform 1 0 11132 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_1_138
timestamp 1608910539
transform 1 0 13800 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 13892 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608910539
transform 1 0 13800 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_1_156
timestamp 1608910539
transform 1 0 15456 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1608910539
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 15916 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608910539
transform 1 0 14996 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608910539
transform 1 0 15548 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608910539
transform 1 0 15088 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608910539
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_174
timestamp 1608910539
transform 1 0 17112 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608910539
transform 1 0 17204 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608910539
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608910539
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608910539
transform 1 0 17388 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608910539
transform 1 0 17756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1608910539
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1608910539
transform 1 0 18492 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1608910539
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_14
timestamp 1608910539
transform 1 0 2392 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1608910539
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1608910539
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1608910539
transform 1 0 1656 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1608910539
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_26 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6624 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5152 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608910539
transform 1 0 8096 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1608910539
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10396 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608910539
transform 1 0 9844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608910539
transform 1 0 8924 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608910539
transform 1 0 12512 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608910539
transform 1 0 12236 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608910539
transform 1 0 11868 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_142
timestamp 1608910539
transform 1 0 14168 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_135
timestamp 1608910539
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_129
timestamp 1608910539
transform 1 0 12972 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_148
timestamp 1608910539
transform 1 0 14720 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608910539
transform 1 0 15548 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_164
timestamp 1608910539
transform 1 0 16192 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 16008 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_167
timestamp 1608910539
transform 1 0 16468 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1608910539
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1608910539
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608910539
transform 1 0 17296 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608910539
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608910539
transform 1 0 16928 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608910539
transform 1 0 17848 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1608910539
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1608910539
transform 1 0 1564 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1608910539
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1608910539
transform 1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_23
timestamp 1608910539
transform 1 0 3220 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1608910539
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 3956 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1608910539
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5428 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_64
timestamp 1608910539
transform 1 0 6992 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7084 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608910539
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1608910539
transform 1 0 10212 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608910539
transform 1 0 10304 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608910539
transform 1 0 9384 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608910539
transform 1 0 11132 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608910539
transform 1 0 12512 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_140
timestamp 1608910539
transform 1 0 13984 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608910539
transform 1 0 14076 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608910539
transform 1 0 12788 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 15272 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1608910539
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1608910539
transform 1 0 17664 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 16468 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1608910539
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_14
timestamp 1608910539
transform 1 0 2392 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1608910539
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1608910539
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1608910539
transform 1 0 1656 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1608910539
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_26
timestamp 1608910539
transform 1 0 3496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4324 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4508 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_61
timestamp 1608910539
transform 1 0 6716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5336 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_73
timestamp 1608910539
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8004 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_95
timestamp 1608910539
transform 1 0 9844 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1608910539
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10212 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_4_115
timestamp 1608910539
transform 1 0 11684 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 12144 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_4_145
timestamp 1608910539
transform 1 0 14444 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_136
timestamp 1608910539
transform 1 0 13616 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608910539
transform 1 0 14168 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608910539
transform 1 0 13340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_4_181
timestamp 1608910539
transform 1 0 17756 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_167
timestamp 1608910539
transform 1 0 16468 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_2_
timestamp 1608910539
transform 1 0 16560 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608910539
transform 1 0 17388 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608910539
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608910539
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1608910539
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2668 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1564 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1608910539
transform 1 0 2116 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_41
timestamp 1608910539
transform 1 0 4876 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 3220 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4048 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5244 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_78
timestamp 1608910539
transform 1 0 8280 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_104
timestamp 1608910539
transform 1 0 10672 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_86
timestamp 1608910539
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9200 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_5_125
timestamp 1608910539
transform 1 0 12604 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_108
timestamp 1608910539
transform 1 0 11040 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 11132 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608910539
transform 1 0 13156 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_5_162
timestamp 1608910539
transform 1 0 16008 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_158
timestamp 1608910539
transform 1 0 15640 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_146
timestamp 1608910539
transform 1 0 14536 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_178
timestamp 1608910539
transform 1 0 17480 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16652 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1608910539
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1608910539
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_10
timestamp 1608910539
transform 1 0 2024 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1608910539
transform 1 0 1472 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1608910539
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1608910539
transform 1 0 2024 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1608910539
transform 1 0 1656 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1608910539
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1608910539
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1608910539
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 2944 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2116 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_6_32
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4140 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 3588 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_47
timestamp 1608910539
transform 1 0 5428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_43
timestamp 1608910539
transform 1 0 5060 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 4968 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 5704 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_54
timestamp 1608910539
transform 1 0 6072 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_62
timestamp 1608910539
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _09_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_73
timestamp 1608910539
transform 1 0 7820 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_65
timestamp 1608910539
transform 1 0 7084 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_75
timestamp 1608910539
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1608910539
transform 1 0 8096 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608910539
transform 1 0 6992 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_87
timestamp 1608910539
transform 1 0 9108 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1608910539
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1608910539
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 9476 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_101
timestamp 1608910539
transform 1 0 10396 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_97
timestamp 1608910539
transform 1 0 10028 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 10120 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_105
timestamp 1608910539
transform 1 0 10764 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_120
timestamp 1608910539
transform 1 0 12144 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1608910539
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 10856 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_138
timestamp 1608910539
transform 1 0 13800 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_134
timestamp 1608910539
transform 1 0 13432 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_143
timestamp 1608910539
transform 1 0 14260 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_126
timestamp 1608910539
transform 1 0 12696 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13892 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12788 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_159
timestamp 1608910539
transform 1 0 15732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_155
timestamp 1608910539
transform 1 0 15364 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608910539
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16008 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15824 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16836 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16652 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1608910539
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17664 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1608910539
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1608910539
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1608910539
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1608910539
transform 1 0 17848 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1608910539
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1608910539
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1608910539
transform 1 0 1472 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1608910539
transform 1 0 2760 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1608910539
transform 1 0 2392 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1608910539
transform 1 0 2024 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1608910539
transform 1 0 1656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1608910539
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1608910539
transform 1 0 3588 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1608910539
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 3680 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4232 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _10_
timestamp 1608910539
transform 1 0 3312 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5888 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_73
timestamp 1608910539
transform 1 0 7820 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_65
timestamp 1608910539
transform 1 0 7084 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1608910539
transform 1 0 8096 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp 1608910539
transform 1 0 10396 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_93
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608910539
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10488 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _13_
timestamp 1608910539
transform 1 0 8924 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_140
timestamp 1608910539
transform 1 0 13984 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1608910539
transform 1 0 14352 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12972 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1608910539
transform 1 0 17572 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1608910539
transform 1 0 16744 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1608910539
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1608910539
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1932 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1608910539
transform 1 0 2944 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1608910539
transform 1 0 1564 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_29
timestamp 1608910539
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3864 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5520 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1608910539
transform 1 0 7636 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 8464 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 9936 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_112
timestamp 1608910539
transform 1 0 11408 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_137
timestamp 1608910539
transform 1 0 13708 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 13800 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _14_
timestamp 1608910539
transform 1 0 13248 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_160
timestamp 1608910539
transform 1 0 15824 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_154
timestamp 1608910539
transform 1 0 15272 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1608910539
transform 1 0 16468 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608910539
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _15_
timestamp 1608910539
transform 1 0 17296 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1608910539
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1608910539
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1608910539
transform 1 0 2208 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1608910539
transform 1 0 1656 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1608910539
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1608910539
transform 1 0 3036 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4876 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5704 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_66
timestamp 1608910539
transform 1 0 7176 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7452 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8280 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1608910539
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1608910539
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10212 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 11684 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12144 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_140
timestamp 1608910539
transform 1 0 13984 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12972 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1608910539
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_181
timestamp 1608910539
transform 1 0 17756 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1608910539
transform 1 0 17572 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16744 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608910539
transform 1 0 18216 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608910539
transform 1 0 17848 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1472 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_22
timestamp 1608910539
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 3496 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1608910539
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_42
timestamp 1608910539
transform 1 0 4968 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 6348 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5520 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_64
timestamp 1608910539
transform 1 0 6992 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8372 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7544 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10212 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1608910539
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_140
timestamp 1608910539
transform 1 0 13984 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12972 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_162
timestamp 1608910539
transform 1 0 16008 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14536 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1608910539
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16744 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608910539
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1608910539
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1608910539
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1840 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1608910539
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_24
timestamp 1608910539
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3680 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 4324 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_43
timestamp 1608910539
transform 1 0 5060 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_82
timestamp 1608910539
transform 1 0 8648 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_64
timestamp 1608910539
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8740 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7176 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_123
timestamp 1608910539
transform 1 0 12420 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_106
timestamp 1608910539
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 12512 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10948 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_12_140
timestamp 1608910539
transform 1 0 13984 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12972 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_160
timestamp 1608910539
transform 1 0 15824 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_154
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1608910539
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 15916 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1608910539
transform 1 0 16468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1608910539
transform 1 0 17572 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16744 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1608910539
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_5
timestamp 1608910539
transform 1 0 1564 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1608910539
transform 1 0 1472 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1608910539
transform 1 0 1656 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_13
timestamp 1608910539
transform 1 0 2300 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_16
timestamp 1608910539
transform 1 0 2576 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1608910539
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1608910539
transform 1 0 2024 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1608910539
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1608910539
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1608910539
transform 1 0 4600 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1608910539
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 5336 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6256 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5428 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5796 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_83
timestamp 1608910539
transform 1 0 8740 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_73
timestamp 1608910539
transform 1 0 7820 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7544 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _12_
timestamp 1608910539
transform 1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_86
timestamp 1608910539
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_102
timestamp 1608910539
transform 1 0 10488 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1608910539
transform 1 0 9660 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1608910539
transform 1 0 9752 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1608910539
transform 1 0 10580 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_110
timestamp 1608910539
transform 1 0 11224 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_106
timestamp 1608910539
transform 1 0 10856 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1608910539
transform 1 0 10948 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_118
timestamp 1608910539
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_123
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1608910539
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12144 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12512 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_135
timestamp 1608910539
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_129
timestamp 1608910539
transform 1 0 12972 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13524 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12696 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 13708 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_148
timestamp 1608910539
transform 1 0 14720 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1608910539
transform 1 0 14812 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15640 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_176
timestamp 1608910539
transform 1 0 17296 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1608910539
transform 1 0 16928 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16468 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1608910539
transform 1 0 17756 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1608910539
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 1472 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2300 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_37
timestamp 1608910539
transform 1 0 4508 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_29
timestamp 1608910539
transform 1 0 3772 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4600 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1608910539
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5428 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 7360 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_100
timestamp 1608910539
transform 1 0 10304 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1608910539
transform 1 0 10580 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 8832 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_112
timestamp 1608910539
transform 1 0 11408 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11500 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12604 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_136
timestamp 1608910539
transform 1 0 13616 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13708 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_153
timestamp 1608910539
transform 1 0 15180 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1608910539
transform 1 0 16284 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1608910539
transform 1 0 17112 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1608910539
transform 1 0 17480 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1608910539
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 1840 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1608910539
transform 1 0 2668 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_28
timestamp 1608910539
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_61
timestamp 1608910539
transform 1 0 6716 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_47
timestamp 1608910539
transform 1 0 5428 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_44
timestamp 1608910539
transform 1 0 5152 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1608910539
transform 1 0 5704 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6808 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_78
timestamp 1608910539
transform 1 0 8280 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_99
timestamp 1608910539
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_93
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10304 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_116
timestamp 1608910539
transform 1 0 11776 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12512 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_140
timestamp 1608910539
transform 1 0 13984 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1608910539
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1608910539
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1608910539
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1472 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1608910539
transform 1 0 2300 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_24
timestamp 1608910539
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 3496 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_58
timestamp 1608910539
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4968 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1608910539
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7728 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1608910539
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1608910539
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1608910539
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1608910539
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1608910539
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1608910539
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1608910539
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1608910539
transform 1 0 1656 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2484 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_50
timestamp 1608910539
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_44
timestamp 1608910539
transform 1 0 5152 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5796 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_79
timestamp 1608910539
transform 1 0 8372 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_67
timestamp 1608910539
transform 1 0 7268 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1608910539
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1608910539
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1608910539
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1608910539
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1608910539
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1608910539
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1608910539
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1608910539
transform 1 0 1932 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1608910539
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_12
timestamp 1608910539
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1608910539
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1608910539
transform 1 0 2300 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_16
timestamp 1608910539
transform 1 0 2576 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1608910539
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1608910539
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1608910539
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1608910539
transform 1 0 3128 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1608910539
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1608910539
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608910539
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608910539
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1608910539
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1608910539
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1608910539
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1608910539
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1608910539
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1608910539
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1608910539
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1608910539
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1608910539
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1608910539
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1608910539
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1608910539
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1608910539
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1608910539
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1608910539
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1608910539
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1608910539
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1608910539
transform 1 0 2392 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1608910539
transform 1 0 2024 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1608910539
transform 1 0 1656 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1608910539
transform 1 0 4048 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1608910539
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1608910539
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1608910539
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1608910539
transform 1 0 3128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_52
timestamp 1608910539
transform 1 0 5888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_44
timestamp 1608910539
transform 1 0 5152 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1608910539
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1608910539
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_78
timestamp 1608910539
transform 1 0 8280 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_66
timestamp 1608910539
transform 1 0 7176 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1608910539
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_102
timestamp 1608910539
transform 1 0 10488 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_90
timestamp 1608910539
transform 1 0 9384 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1608910539
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_144
timestamp 1608910539
transform 1 0 14352 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1608910539
transform 1 0 13984 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1608910539
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608910539
transform 1 0 14444 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608910539
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_161
timestamp 1608910539
transform 1 0 15916 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1608910539
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608910539
transform 1 0 15548 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608910539
transform 1 0 15180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_184
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1608910539
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_173
timestamp 1608910539
transform 1 0 17020 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1608910539
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608910539
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1608910539
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1608910539
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1608910539
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1608910539
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1608910539
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1608910539
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1608910539
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1608910539
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1608910539
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1608910539
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1608910539
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1608910539
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1608910539
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_180
timestamp 1608910539
transform 1 0 17664 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1608910539
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 7378 16400 7434 17200 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 SC_IN_BOT
port 1 nsew signal input
rlabel metal2 s 6090 16400 6146 17200 6 SC_IN_TOP
port 2 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 SC_OUT_BOT
port 3 nsew signal tristate
rlabel metal2 s 6734 16400 6790 17200 6 SC_OUT_TOP
port 4 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 bottom_grid_pin_0_
port 5 nsew signal tristate
rlabel metal2 s 2686 0 2742 800 6 bottom_grid_pin_10_
port 6 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 bottom_grid_pin_12_
port 7 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 bottom_grid_pin_14_
port 8 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 bottom_grid_pin_16_
port 9 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 bottom_grid_pin_2_
port 10 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 bottom_grid_pin_4_
port 11 nsew signal tristate
rlabel metal2 s 1674 0 1730 800 6 bottom_grid_pin_6_
port 12 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 bottom_grid_pin_8_
port 13 nsew signal tristate
rlabel metal2 s 4618 0 4674 800 6 ccff_head
port 14 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 ccff_tail
port 15 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[0]
port 16 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[10]
port 17 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_in[11]
port 18 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 chanx_left_in[12]
port 19 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 chanx_left_in[13]
port 20 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 chanx_left_in[14]
port 21 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 chanx_left_in[15]
port 22 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 chanx_left_in[16]
port 23 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 chanx_left_in[17]
port 24 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 chanx_left_in[18]
port 25 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 chanx_left_in[19]
port 26 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[1]
port 27 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[2]
port 28 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[3]
port 29 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[4]
port 30 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[5]
port 31 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[6]
port 32 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[7]
port 33 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[8]
port 34 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[9]
port 35 nsew signal input
rlabel metal3 s 0 552 800 672 6 chanx_left_out[0]
port 36 nsew signal tristate
rlabel metal3 s 0 4632 800 4752 6 chanx_left_out[10]
port 37 nsew signal tristate
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[11]
port 38 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 chanx_left_out[12]
port 39 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 chanx_left_out[13]
port 40 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[14]
port 41 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 chanx_left_out[15]
port 42 nsew signal tristate
rlabel metal3 s 0 7216 800 7336 6 chanx_left_out[16]
port 43 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 chanx_left_out[17]
port 44 nsew signal tristate
rlabel metal3 s 0 8032 800 8152 6 chanx_left_out[18]
port 45 nsew signal tristate
rlabel metal3 s 0 8440 800 8560 6 chanx_left_out[19]
port 46 nsew signal tristate
rlabel metal3 s 0 960 800 1080 6 chanx_left_out[1]
port 47 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 chanx_left_out[2]
port 48 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[3]
port 49 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 chanx_left_out[4]
port 50 nsew signal tristate
rlabel metal3 s 0 2592 800 2712 6 chanx_left_out[5]
port 51 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 chanx_left_out[6]
port 52 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[7]
port 53 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_out[8]
port 54 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 chanx_left_out[9]
port 55 nsew signal tristate
rlabel metal3 s 19200 8712 20000 8832 6 chanx_right_in[0]
port 56 nsew signal input
rlabel metal3 s 19200 12928 20000 13048 6 chanx_right_in[10]
port 57 nsew signal input
rlabel metal3 s 19200 13336 20000 13456 6 chanx_right_in[11]
port 58 nsew signal input
rlabel metal3 s 19200 13744 20000 13864 6 chanx_right_in[12]
port 59 nsew signal input
rlabel metal3 s 19200 14152 20000 14272 6 chanx_right_in[13]
port 60 nsew signal input
rlabel metal3 s 19200 14696 20000 14816 6 chanx_right_in[14]
port 61 nsew signal input
rlabel metal3 s 19200 15104 20000 15224 6 chanx_right_in[15]
port 62 nsew signal input
rlabel metal3 s 19200 15512 20000 15632 6 chanx_right_in[16]
port 63 nsew signal input
rlabel metal3 s 19200 15920 20000 16040 6 chanx_right_in[17]
port 64 nsew signal input
rlabel metal3 s 19200 16328 20000 16448 6 chanx_right_in[18]
port 65 nsew signal input
rlabel metal3 s 19200 16736 20000 16856 6 chanx_right_in[19]
port 66 nsew signal input
rlabel metal3 s 19200 9120 20000 9240 6 chanx_right_in[1]
port 67 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 chanx_right_in[2]
port 68 nsew signal input
rlabel metal3 s 19200 9936 20000 10056 6 chanx_right_in[3]
port 69 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[4]
port 70 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[5]
port 71 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[6]
port 72 nsew signal input
rlabel metal3 s 19200 11704 20000 11824 6 chanx_right_in[7]
port 73 nsew signal input
rlabel metal3 s 19200 12112 20000 12232 6 chanx_right_in[8]
port 74 nsew signal input
rlabel metal3 s 19200 12520 20000 12640 6 chanx_right_in[9]
port 75 nsew signal input
rlabel metal3 s 19200 144 20000 264 6 chanx_right_out[0]
port 76 nsew signal tristate
rlabel metal3 s 19200 4360 20000 4480 6 chanx_right_out[10]
port 77 nsew signal tristate
rlabel metal3 s 19200 4768 20000 4888 6 chanx_right_out[11]
port 78 nsew signal tristate
rlabel metal3 s 19200 5176 20000 5296 6 chanx_right_out[12]
port 79 nsew signal tristate
rlabel metal3 s 19200 5584 20000 5704 6 chanx_right_out[13]
port 80 nsew signal tristate
rlabel metal3 s 19200 6128 20000 6248 6 chanx_right_out[14]
port 81 nsew signal tristate
rlabel metal3 s 19200 6536 20000 6656 6 chanx_right_out[15]
port 82 nsew signal tristate
rlabel metal3 s 19200 6944 20000 7064 6 chanx_right_out[16]
port 83 nsew signal tristate
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[17]
port 84 nsew signal tristate
rlabel metal3 s 19200 7760 20000 7880 6 chanx_right_out[18]
port 85 nsew signal tristate
rlabel metal3 s 19200 8168 20000 8288 6 chanx_right_out[19]
port 86 nsew signal tristate
rlabel metal3 s 19200 552 20000 672 6 chanx_right_out[1]
port 87 nsew signal tristate
rlabel metal3 s 19200 960 20000 1080 6 chanx_right_out[2]
port 88 nsew signal tristate
rlabel metal3 s 19200 1368 20000 1488 6 chanx_right_out[3]
port 89 nsew signal tristate
rlabel metal3 s 19200 1776 20000 1896 6 chanx_right_out[4]
port 90 nsew signal tristate
rlabel metal3 s 19200 2184 20000 2304 6 chanx_right_out[5]
port 91 nsew signal tristate
rlabel metal3 s 19200 2592 20000 2712 6 chanx_right_out[6]
port 92 nsew signal tristate
rlabel metal3 s 19200 3136 20000 3256 6 chanx_right_out[7]
port 93 nsew signal tristate
rlabel metal3 s 19200 3544 20000 3664 6 chanx_right_out[8]
port 94 nsew signal tristate
rlabel metal3 s 19200 3952 20000 4072 6 chanx_right_out[9]
port 95 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 96 nsew signal tristate
rlabel metal2 s 7102 0 7158 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 97 nsew signal tristate
rlabel metal2 s 7654 0 7710 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 98 nsew signal tristate
rlabel metal2 s 8114 0 8170 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 99 nsew signal tristate
rlabel metal2 s 8666 0 8722 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 100 nsew signal tristate
rlabel metal2 s 9126 0 9182 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 101 nsew signal tristate
rlabel metal2 s 9678 0 9734 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 102 nsew signal tristate
rlabel metal2 s 10138 0 10194 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 103 nsew signal tristate
rlabel metal2 s 10598 0 10654 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 104 nsew signal tristate
rlabel metal2 s 11150 0 11206 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 105 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 106 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 107 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 108 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 109 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 110 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 111 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 112 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 113 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 114 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 115 nsew signal tristate
rlabel metal2 s 16670 0 16726 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 116 nsew signal tristate
rlabel metal2 s 17130 0 17186 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 117 nsew signal tristate
rlabel metal2 s 17590 0 17646 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 118 nsew signal tristate
rlabel metal2 s 18142 0 18198 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 119 nsew signal tristate
rlabel metal2 s 18602 0 18658 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 120 nsew signal tristate
rlabel metal2 s 19154 0 19210 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 121 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 122 nsew signal tristate
rlabel metal2 s 8022 16400 8078 17200 6 prog_clk_0_N_in
port 123 nsew signal input
rlabel metal3 s 0 144 800 264 6 prog_clk_0_W_out
port 124 nsew signal tristate
rlabel metal2 s 8666 16400 8722 17200 6 top_width_0_height_0__pin_0_
port 125 nsew signal input
rlabel metal2 s 11886 16400 11942 17200 6 top_width_0_height_0__pin_10_
port 126 nsew signal input
rlabel metal2 s 14462 16400 14518 17200 6 top_width_0_height_0__pin_11_lower
port 127 nsew signal tristate
rlabel metal2 s 3514 16400 3570 17200 6 top_width_0_height_0__pin_11_upper
port 128 nsew signal tristate
rlabel metal2 s 12530 16400 12586 17200 6 top_width_0_height_0__pin_12_
port 129 nsew signal input
rlabel metal2 s 15106 16400 15162 17200 6 top_width_0_height_0__pin_13_lower
port 130 nsew signal tristate
rlabel metal2 s 4158 16400 4214 17200 6 top_width_0_height_0__pin_13_upper
port 131 nsew signal tristate
rlabel metal2 s 13174 16400 13230 17200 6 top_width_0_height_0__pin_14_
port 132 nsew signal input
rlabel metal2 s 15750 16400 15806 17200 6 top_width_0_height_0__pin_15_lower
port 133 nsew signal tristate
rlabel metal2 s 4802 16400 4858 17200 6 top_width_0_height_0__pin_15_upper
port 134 nsew signal tristate
rlabel metal2 s 13818 16400 13874 17200 6 top_width_0_height_0__pin_16_
port 135 nsew signal input
rlabel metal2 s 16394 16400 16450 17200 6 top_width_0_height_0__pin_17_lower
port 136 nsew signal tristate
rlabel metal2 s 5446 16400 5502 17200 6 top_width_0_height_0__pin_17_upper
port 137 nsew signal tristate
rlabel metal2 s 17038 16400 17094 17200 6 top_width_0_height_0__pin_1_lower
port 138 nsew signal tristate
rlabel metal2 s 294 16400 350 17200 6 top_width_0_height_0__pin_1_upper
port 139 nsew signal tristate
rlabel metal2 s 9310 16400 9366 17200 6 top_width_0_height_0__pin_2_
port 140 nsew signal input
rlabel metal2 s 17682 16400 17738 17200 6 top_width_0_height_0__pin_3_lower
port 141 nsew signal tristate
rlabel metal2 s 938 16400 994 17200 6 top_width_0_height_0__pin_3_upper
port 142 nsew signal tristate
rlabel metal2 s 9954 16400 10010 17200 6 top_width_0_height_0__pin_4_
port 143 nsew signal input
rlabel metal2 s 18326 16400 18382 17200 6 top_width_0_height_0__pin_5_lower
port 144 nsew signal tristate
rlabel metal2 s 1582 16400 1638 17200 6 top_width_0_height_0__pin_5_upper
port 145 nsew signal tristate
rlabel metal2 s 10598 16400 10654 17200 6 top_width_0_height_0__pin_6_
port 146 nsew signal input
rlabel metal2 s 18970 16400 19026 17200 6 top_width_0_height_0__pin_7_lower
port 147 nsew signal tristate
rlabel metal2 s 2226 16400 2282 17200 6 top_width_0_height_0__pin_7_upper
port 148 nsew signal tristate
rlabel metal2 s 11242 16400 11298 17200 6 top_width_0_height_0__pin_8_
port 149 nsew signal input
rlabel metal2 s 19614 16400 19670 17200 6 top_width_0_height_0__pin_9_lower
port 150 nsew signal tristate
rlabel metal2 s 2870 16400 2926 17200 6 top_width_0_height_0__pin_9_upper
port 151 nsew signal tristate
rlabel metal4 s 15771 2128 16091 14736 6 VPWR
port 152 nsew power bidirectional
rlabel metal4 s 9840 2128 10160 14736 6 VPWR
port 153 nsew power bidirectional
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 154 nsew power bidirectional
rlabel metal4 s 12805 2128 13125 14736 6 VGND
port 155 nsew ground bidirectional
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 156 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
