VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.000 BY 110.000 ;
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 2.400 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 107.600 105.250 110.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.400 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 107.600 108.470 110.000 ;
    END
  END SC_OUT_TOP
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.400 ;
    END
  END Test_en
  PIN bottom_width_0_height_0__pin_50_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END bottom_width_0_height_0__pin_50_
  PIN bottom_width_0_height_0__pin_51_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.400 ;
    END
  END bottom_width_0_height_0__pin_51_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 27.920 110.000 28.520 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 2.400 ;
    END
  END clk
  PIN left_width_0_height_0__pin_52_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 2.400 92.440 ;
    END
  END left_width_0_height_0__pin_52_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.400 19.000 ;
    END
  END prog_clk
  PIN right_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 31.320 110.000 31.920 ;
    END
  END right_width_0_height_0__pin_16_
  PIN right_width_0_height_0__pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 34.720 110.000 35.320 ;
    END
  END right_width_0_height_0__pin_17_
  PIN right_width_0_height_0__pin_18_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 38.120 110.000 38.720 ;
    END
  END right_width_0_height_0__pin_18_
  PIN right_width_0_height_0__pin_19_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 40.840 110.000 41.440 ;
    END
  END right_width_0_height_0__pin_19_
  PIN right_width_0_height_0__pin_20_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 44.240 110.000 44.840 ;
    END
  END right_width_0_height_0__pin_20_
  PIN right_width_0_height_0__pin_21_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 47.640 110.000 48.240 ;
    END
  END right_width_0_height_0__pin_21_
  PIN right_width_0_height_0__pin_22_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 51.040 110.000 51.640 ;
    END
  END right_width_0_height_0__pin_22_
  PIN right_width_0_height_0__pin_23_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 54.440 110.000 55.040 ;
    END
  END right_width_0_height_0__pin_23_
  PIN right_width_0_height_0__pin_24_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 57.840 110.000 58.440 ;
    END
  END right_width_0_height_0__pin_24_
  PIN right_width_0_height_0__pin_25_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 61.240 110.000 61.840 ;
    END
  END right_width_0_height_0__pin_25_
  PIN right_width_0_height_0__pin_26_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 64.640 110.000 65.240 ;
    END
  END right_width_0_height_0__pin_26_
  PIN right_width_0_height_0__pin_27_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 68.040 110.000 68.640 ;
    END
  END right_width_0_height_0__pin_27_
  PIN right_width_0_height_0__pin_28_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 71.440 110.000 72.040 ;
    END
  END right_width_0_height_0__pin_28_
  PIN right_width_0_height_0__pin_29_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 74.840 110.000 75.440 ;
    END
  END right_width_0_height_0__pin_29_
  PIN right_width_0_height_0__pin_30_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 77.560 110.000 78.160 ;
    END
  END right_width_0_height_0__pin_30_
  PIN right_width_0_height_0__pin_31_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 80.960 110.000 81.560 ;
    END
  END right_width_0_height_0__pin_31_
  PIN right_width_0_height_0__pin_42_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 1.400 110.000 2.000 ;
    END
  END right_width_0_height_0__pin_42_lower
  PIN right_width_0_height_0__pin_42_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 84.360 110.000 84.960 ;
    END
  END right_width_0_height_0__pin_42_upper
  PIN right_width_0_height_0__pin_43_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 4.120 110.000 4.720 ;
    END
  END right_width_0_height_0__pin_43_lower
  PIN right_width_0_height_0__pin_43_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 87.760 110.000 88.360 ;
    END
  END right_width_0_height_0__pin_43_upper
  PIN right_width_0_height_0__pin_44_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 7.520 110.000 8.120 ;
    END
  END right_width_0_height_0__pin_44_lower
  PIN right_width_0_height_0__pin_44_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 91.160 110.000 91.760 ;
    END
  END right_width_0_height_0__pin_44_upper
  PIN right_width_0_height_0__pin_45_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 10.920 110.000 11.520 ;
    END
  END right_width_0_height_0__pin_45_lower
  PIN right_width_0_height_0__pin_45_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 94.560 110.000 95.160 ;
    END
  END right_width_0_height_0__pin_45_upper
  PIN right_width_0_height_0__pin_46_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 14.320 110.000 14.920 ;
    END
  END right_width_0_height_0__pin_46_lower
  PIN right_width_0_height_0__pin_46_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 97.960 110.000 98.560 ;
    END
  END right_width_0_height_0__pin_46_upper
  PIN right_width_0_height_0__pin_47_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 17.720 110.000 18.320 ;
    END
  END right_width_0_height_0__pin_47_lower
  PIN right_width_0_height_0__pin_47_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 101.360 110.000 101.960 ;
    END
  END right_width_0_height_0__pin_47_upper
  PIN right_width_0_height_0__pin_48_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 21.120 110.000 21.720 ;
    END
  END right_width_0_height_0__pin_48_lower
  PIN right_width_0_height_0__pin_48_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 104.760 110.000 105.360 ;
    END
  END right_width_0_height_0__pin_48_upper
  PIN right_width_0_height_0__pin_49_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 24.520 110.000 25.120 ;
    END
  END right_width_0_height_0__pin_49_lower
  PIN right_width_0_height_0__pin_49_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 108.160 110.000 108.760 ;
    END
  END right_width_0_height_0__pin_49_upper
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 107.600 26.130 110.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 107.600 56.490 110.000 ;
    END
  END top_width_0_height_0__pin_10_
  PIN top_width_0_height_0__pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 107.600 59.710 110.000 ;
    END
  END top_width_0_height_0__pin_11_
  PIN top_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 107.600 62.470 110.000 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 107.600 65.690 110.000 ;
    END
  END top_width_0_height_0__pin_13_
  PIN top_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 107.600 68.910 110.000 ;
    END
  END top_width_0_height_0__pin_14_
  PIN top_width_0_height_0__pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.390 107.600 71.670 110.000 ;
    END
  END top_width_0_height_0__pin_15_
  PIN top_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 107.600 28.890 110.000 ;
    END
  END top_width_0_height_0__pin_1_
  PIN top_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 107.600 32.110 110.000 ;
    END
  END top_width_0_height_0__pin_2_
  PIN top_width_0_height_0__pin_32_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 107.600 74.890 110.000 ;
    END
  END top_width_0_height_0__pin_32_
  PIN top_width_0_height_0__pin_33_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 107.600 77.650 110.000 ;
    END
  END top_width_0_height_0__pin_33_
  PIN top_width_0_height_0__pin_34_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.590 107.600 80.870 110.000 ;
    END
  END top_width_0_height_0__pin_34_lower
  PIN top_width_0_height_0__pin_34_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.470 107.600 1.750 110.000 ;
    END
  END top_width_0_height_0__pin_34_upper
  PIN top_width_0_height_0__pin_35_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 107.600 84.090 110.000 ;
    END
  END top_width_0_height_0__pin_35_lower
  PIN top_width_0_height_0__pin_35_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.230 107.600 4.510 110.000 ;
    END
  END top_width_0_height_0__pin_35_upper
  PIN top_width_0_height_0__pin_36_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 107.600 86.850 110.000 ;
    END
  END top_width_0_height_0__pin_36_lower
  PIN top_width_0_height_0__pin_36_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 107.600 7.730 110.000 ;
    END
  END top_width_0_height_0__pin_36_upper
  PIN top_width_0_height_0__pin_37_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 107.600 90.070 110.000 ;
    END
  END top_width_0_height_0__pin_37_lower
  PIN top_width_0_height_0__pin_37_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.210 107.600 10.490 110.000 ;
    END
  END top_width_0_height_0__pin_37_upper
  PIN top_width_0_height_0__pin_38_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 107.600 93.290 110.000 ;
    END
  END top_width_0_height_0__pin_38_lower
  PIN top_width_0_height_0__pin_38_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.430 107.600 13.710 110.000 ;
    END
  END top_width_0_height_0__pin_38_upper
  PIN top_width_0_height_0__pin_39_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 107.600 96.050 110.000 ;
    END
  END top_width_0_height_0__pin_39_lower
  PIN top_width_0_height_0__pin_39_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.650 107.600 16.930 110.000 ;
    END
  END top_width_0_height_0__pin_39_upper
  PIN top_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 107.600 35.330 110.000 ;
    END
  END top_width_0_height_0__pin_3_
  PIN top_width_0_height_0__pin_40_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 107.600 99.270 110.000 ;
    END
  END top_width_0_height_0__pin_40_lower
  PIN top_width_0_height_0__pin_40_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 107.600 19.690 110.000 ;
    END
  END top_width_0_height_0__pin_40_upper
  PIN top_width_0_height_0__pin_41_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 107.600 102.490 110.000 ;
    END
  END top_width_0_height_0__pin_41_lower
  PIN top_width_0_height_0__pin_41_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.630 107.600 22.910 110.000 ;
    END
  END top_width_0_height_0__pin_41_upper
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 107.600 38.090 110.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 107.600 41.310 110.000 ;
    END
  END top_width_0_height_0__pin_5_
  PIN top_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 107.600 44.070 110.000 ;
    END
  END top_width_0_height_0__pin_6_
  PIN top_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 107.600 47.290 110.000 ;
    END
  END top_width_0_height_0__pin_7_
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 107.600 50.510 110.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN top_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 107.600 53.270 110.000 ;
    END
  END top_width_0_height_0__pin_9_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.215 10.640 22.815 98.160 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 37.705 10.640 39.305 98.160 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 105.195 98.005 ;
      LAYER met1 ;
        RECT 1.450 6.160 108.490 98.560 ;
      LAYER met2 ;
        RECT 2.030 107.320 3.950 108.645 ;
        RECT 4.790 107.320 7.170 108.645 ;
        RECT 8.010 107.320 9.930 108.645 ;
        RECT 10.770 107.320 13.150 108.645 ;
        RECT 13.990 107.320 16.370 108.645 ;
        RECT 17.210 107.320 19.130 108.645 ;
        RECT 19.970 107.320 22.350 108.645 ;
        RECT 23.190 107.320 25.570 108.645 ;
        RECT 26.410 107.320 28.330 108.645 ;
        RECT 29.170 107.320 31.550 108.645 ;
        RECT 32.390 107.320 34.770 108.645 ;
        RECT 35.610 107.320 37.530 108.645 ;
        RECT 38.370 107.320 40.750 108.645 ;
        RECT 41.590 107.320 43.510 108.645 ;
        RECT 44.350 107.320 46.730 108.645 ;
        RECT 47.570 107.320 49.950 108.645 ;
        RECT 50.790 107.320 52.710 108.645 ;
        RECT 53.550 107.320 55.930 108.645 ;
        RECT 56.770 107.320 59.150 108.645 ;
        RECT 59.990 107.320 61.910 108.645 ;
        RECT 62.750 107.320 65.130 108.645 ;
        RECT 65.970 107.320 68.350 108.645 ;
        RECT 69.190 107.320 71.110 108.645 ;
        RECT 71.950 107.320 74.330 108.645 ;
        RECT 75.170 107.320 77.090 108.645 ;
        RECT 77.930 107.320 80.310 108.645 ;
        RECT 81.150 107.320 83.530 108.645 ;
        RECT 84.370 107.320 86.290 108.645 ;
        RECT 87.130 107.320 89.510 108.645 ;
        RECT 90.350 107.320 92.730 108.645 ;
        RECT 93.570 107.320 95.490 108.645 ;
        RECT 96.330 107.320 98.710 108.645 ;
        RECT 99.550 107.320 101.930 108.645 ;
        RECT 102.770 107.320 104.690 108.645 ;
        RECT 105.530 107.320 107.910 108.645 ;
        RECT 1.480 2.680 108.460 107.320 ;
        RECT 1.480 1.515 8.550 2.680 ;
        RECT 9.390 1.515 26.490 2.680 ;
        RECT 27.330 1.515 44.890 2.680 ;
        RECT 45.730 1.515 63.290 2.680 ;
        RECT 64.130 1.515 81.690 2.680 ;
        RECT 82.530 1.515 100.090 2.680 ;
        RECT 100.930 1.515 108.460 2.680 ;
      LAYER met3 ;
        RECT 2.400 107.760 107.200 108.625 ;
        RECT 2.400 105.760 107.600 107.760 ;
        RECT 2.400 104.360 107.200 105.760 ;
        RECT 2.400 102.360 107.600 104.360 ;
        RECT 2.400 100.960 107.200 102.360 ;
        RECT 2.400 98.960 107.600 100.960 ;
        RECT 2.400 97.560 107.200 98.960 ;
        RECT 2.400 95.560 107.600 97.560 ;
        RECT 2.400 94.160 107.200 95.560 ;
        RECT 2.400 92.840 107.600 94.160 ;
        RECT 2.800 92.160 107.600 92.840 ;
        RECT 2.800 91.440 107.200 92.160 ;
        RECT 2.400 90.760 107.200 91.440 ;
        RECT 2.400 88.760 107.600 90.760 ;
        RECT 2.400 87.360 107.200 88.760 ;
        RECT 2.400 85.360 107.600 87.360 ;
        RECT 2.400 83.960 107.200 85.360 ;
        RECT 2.400 81.960 107.600 83.960 ;
        RECT 2.400 80.560 107.200 81.960 ;
        RECT 2.400 78.560 107.600 80.560 ;
        RECT 2.400 77.160 107.200 78.560 ;
        RECT 2.400 75.840 107.600 77.160 ;
        RECT 2.400 74.440 107.200 75.840 ;
        RECT 2.400 72.440 107.600 74.440 ;
        RECT 2.400 71.040 107.200 72.440 ;
        RECT 2.400 69.040 107.600 71.040 ;
        RECT 2.400 67.640 107.200 69.040 ;
        RECT 2.400 65.640 107.600 67.640 ;
        RECT 2.400 64.240 107.200 65.640 ;
        RECT 2.400 62.240 107.600 64.240 ;
        RECT 2.400 60.840 107.200 62.240 ;
        RECT 2.400 58.840 107.600 60.840 ;
        RECT 2.400 57.440 107.200 58.840 ;
        RECT 2.400 56.120 107.600 57.440 ;
        RECT 2.800 55.440 107.600 56.120 ;
        RECT 2.800 54.720 107.200 55.440 ;
        RECT 2.400 54.040 107.200 54.720 ;
        RECT 2.400 52.040 107.600 54.040 ;
        RECT 2.400 50.640 107.200 52.040 ;
        RECT 2.400 48.640 107.600 50.640 ;
        RECT 2.400 47.240 107.200 48.640 ;
        RECT 2.400 45.240 107.600 47.240 ;
        RECT 2.400 43.840 107.200 45.240 ;
        RECT 2.400 41.840 107.600 43.840 ;
        RECT 2.400 40.440 107.200 41.840 ;
        RECT 2.400 39.120 107.600 40.440 ;
        RECT 2.400 37.720 107.200 39.120 ;
        RECT 2.400 35.720 107.600 37.720 ;
        RECT 2.400 34.320 107.200 35.720 ;
        RECT 2.400 32.320 107.600 34.320 ;
        RECT 2.400 30.920 107.200 32.320 ;
        RECT 2.400 28.920 107.600 30.920 ;
        RECT 2.400 27.520 107.200 28.920 ;
        RECT 2.400 25.520 107.600 27.520 ;
        RECT 2.400 24.120 107.200 25.520 ;
        RECT 2.400 22.120 107.600 24.120 ;
        RECT 2.400 20.720 107.200 22.120 ;
        RECT 2.400 19.400 107.600 20.720 ;
        RECT 2.800 18.720 107.600 19.400 ;
        RECT 2.800 18.000 107.200 18.720 ;
        RECT 2.400 17.320 107.200 18.000 ;
        RECT 2.400 15.320 107.600 17.320 ;
        RECT 2.400 13.920 107.200 15.320 ;
        RECT 2.400 11.920 107.600 13.920 ;
        RECT 2.400 10.520 107.200 11.920 ;
        RECT 2.400 8.520 107.600 10.520 ;
        RECT 2.400 7.120 107.200 8.520 ;
        RECT 2.400 5.120 107.600 7.120 ;
        RECT 2.400 3.720 107.200 5.120 ;
        RECT 2.400 2.400 107.600 3.720 ;
        RECT 2.400 1.535 107.200 2.400 ;
      LAYER met4 ;
        RECT 23.215 10.640 37.305 98.160 ;
        RECT 39.705 10.640 88.785 98.160 ;
  END
END grid_clb
END LIBRARY

