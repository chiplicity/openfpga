VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decoder6to61
  CLASS BLOCK ;
  FOREIGN decoder6to61 ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 117.600 3.130 120.000 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 117.600 9.110 120.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 2.760 120.000 3.360 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 8.200 120.000 8.800 ;
    END
  END address[5]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 14.320 120.000 14.920 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 32.680 120.000 33.280 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 117.600 27.970 120.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 2.400 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 38.120 120.000 38.720 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 44.240 120.000 44.840 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.130 117.600 34.410 120.000 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.570 117.600 40.850 120.000 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.010 117.600 47.290 120.000 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 2.400 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 50.360 120.000 50.960 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 2.400 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 56.480 120.000 57.080 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 2.400 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 62.600 120.000 63.200 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.990 117.600 53.270 120.000 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 68.040 120.000 68.640 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.430 117.600 59.710 120.000 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 117.600 66.150 120.000 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 2.400 29.880 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 74.160 120.000 74.760 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 2.400 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.310 117.600 72.590 120.000 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 2.400 46.880 ;
    END
  END data_out[31]
  PIN data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END data_out[32]
  PIN data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 80.280 120.000 80.880 ;
    END
  END data_out[33]
  PIN data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END data_out[34]
  PIN data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 117.600 78.570 120.000 ;
    END
  END data_out[35]
  PIN data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 2.400 72.720 ;
    END
  END data_out[36]
  PIN data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 86.400 120.000 87.000 ;
    END
  END data_out[37]
  PIN data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 2.400 81.560 ;
    END
  END data_out[38]
  PIN data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.400 ;
    END
  END data_out[39]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.400 ;
    END
  END data_out[3]
  PIN data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 2.400 89.720 ;
    END
  END data_out[40]
  PIN data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 2.400 98.560 ;
    END
  END data_out[41]
  PIN data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 92.520 120.000 93.120 ;
    END
  END data_out[42]
  PIN data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 97.960 120.000 98.560 ;
    END
  END data_out[43]
  PIN data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 104.080 120.000 104.680 ;
    END
  END data_out[44]
  PIN data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 2.400 ;
    END
  END data_out[45]
  PIN data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 117.600 85.010 120.000 ;
    END
  END data_out[46]
  PIN data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 117.600 91.450 120.000 ;
    END
  END data_out[47]
  PIN data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 117.600 97.890 120.000 ;
    END
  END data_out[48]
  PIN data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.400 106.720 ;
    END
  END data_out[49]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 20.440 120.000 21.040 ;
    END
  END data_out[4]
  PIN data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 117.600 103.870 120.000 ;
    END
  END data_out[50]
  PIN data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.400 ;
    END
  END data_out[51]
  PIN data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 2.400 ;
    END
  END data_out[52]
  PIN data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 2.400 ;
    END
  END data_out[53]
  PIN data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.030 117.600 110.310 120.000 ;
    END
  END data_out[54]
  PIN data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 2.400 ;
    END
  END data_out[55]
  PIN data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 110.200 120.000 110.800 ;
    END
  END data_out[56]
  PIN data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 116.320 120.000 116.920 ;
    END
  END data_out[57]
  PIN data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 2.400 115.560 ;
    END
  END data_out[58]
  PIN data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.470 117.600 116.750 120.000 ;
    END
  END data_out[59]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END data_out[5]
  PIN data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 2.400 ;
    END
  END data_out[60]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.270 117.600 15.550 120.000 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 26.560 120.000 27.160 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 21.710 117.600 21.990 120.000 ;
    END
  END data_out[9]
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 2.400 ;
    END
  END enable
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 24.720 10.640 26.320 109.040 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 44.720 10.640 46.320 109.040 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 114.080 108.885 ;
      LAYER met1 ;
        RECT 0.530 10.640 118.150 116.240 ;
      LAYER met2 ;
        RECT 0.550 117.320 2.570 118.050 ;
        RECT 3.410 117.320 8.550 118.050 ;
        RECT 9.390 117.320 14.990 118.050 ;
        RECT 15.830 117.320 21.430 118.050 ;
        RECT 22.270 117.320 27.410 118.050 ;
        RECT 28.250 117.320 33.850 118.050 ;
        RECT 34.690 117.320 40.290 118.050 ;
        RECT 41.130 117.320 46.730 118.050 ;
        RECT 47.570 117.320 52.710 118.050 ;
        RECT 53.550 117.320 59.150 118.050 ;
        RECT 59.990 117.320 65.590 118.050 ;
        RECT 66.430 117.320 72.030 118.050 ;
        RECT 72.870 117.320 78.010 118.050 ;
        RECT 78.850 117.320 84.450 118.050 ;
        RECT 85.290 117.320 90.890 118.050 ;
        RECT 91.730 117.320 97.330 118.050 ;
        RECT 98.170 117.320 103.310 118.050 ;
        RECT 104.150 117.320 109.750 118.050 ;
        RECT 110.590 117.320 116.190 118.050 ;
        RECT 117.030 117.320 118.590 118.050 ;
        RECT 0.550 2.680 118.590 117.320 ;
        RECT 0.550 0.270 3.490 2.680 ;
        RECT 4.330 0.270 11.310 2.680 ;
        RECT 12.150 0.270 19.130 2.680 ;
        RECT 19.970 0.270 27.410 2.680 ;
        RECT 28.250 0.270 35.230 2.680 ;
        RECT 36.070 0.270 43.510 2.680 ;
        RECT 44.350 0.270 51.330 2.680 ;
        RECT 52.170 0.270 59.150 2.680 ;
        RECT 59.990 0.270 67.430 2.680 ;
        RECT 68.270 0.270 75.250 2.680 ;
        RECT 76.090 0.270 83.530 2.680 ;
        RECT 84.370 0.270 91.350 2.680 ;
        RECT 92.190 0.270 99.170 2.680 ;
        RECT 100.010 0.270 107.450 2.680 ;
        RECT 108.290 0.270 115.270 2.680 ;
        RECT 116.110 0.270 118.590 2.680 ;
      LAYER met3 ;
        RECT 0.310 115.960 117.200 116.320 ;
        RECT 2.800 115.920 117.200 115.960 ;
        RECT 2.800 114.560 118.370 115.920 ;
        RECT 0.310 111.200 118.370 114.560 ;
        RECT 0.310 109.800 117.200 111.200 ;
        RECT 0.310 107.120 118.370 109.800 ;
        RECT 2.800 105.720 118.370 107.120 ;
        RECT 0.310 105.080 118.370 105.720 ;
        RECT 0.310 103.680 117.200 105.080 ;
        RECT 0.310 98.960 118.370 103.680 ;
        RECT 2.800 97.560 117.200 98.960 ;
        RECT 0.310 93.520 118.370 97.560 ;
        RECT 0.310 92.120 117.200 93.520 ;
        RECT 0.310 90.120 118.370 92.120 ;
        RECT 2.800 88.720 118.370 90.120 ;
        RECT 0.310 87.400 118.370 88.720 ;
        RECT 0.310 86.000 117.200 87.400 ;
        RECT 0.310 81.960 118.370 86.000 ;
        RECT 2.800 81.280 118.370 81.960 ;
        RECT 2.800 80.560 117.200 81.280 ;
        RECT 0.310 79.880 117.200 80.560 ;
        RECT 0.310 75.160 118.370 79.880 ;
        RECT 0.310 73.760 117.200 75.160 ;
        RECT 0.310 73.120 118.370 73.760 ;
        RECT 2.800 71.720 118.370 73.120 ;
        RECT 0.310 69.040 118.370 71.720 ;
        RECT 0.310 67.640 117.200 69.040 ;
        RECT 0.310 64.960 118.370 67.640 ;
        RECT 2.800 63.600 118.370 64.960 ;
        RECT 2.800 63.560 117.200 63.600 ;
        RECT 0.310 62.200 117.200 63.560 ;
        RECT 0.310 57.480 118.370 62.200 ;
        RECT 0.310 56.120 117.200 57.480 ;
        RECT 2.800 56.080 117.200 56.120 ;
        RECT 2.800 54.720 118.370 56.080 ;
        RECT 0.310 51.360 118.370 54.720 ;
        RECT 0.310 49.960 117.200 51.360 ;
        RECT 0.310 47.280 118.370 49.960 ;
        RECT 2.800 45.880 118.370 47.280 ;
        RECT 0.310 45.240 118.370 45.880 ;
        RECT 0.310 43.840 117.200 45.240 ;
        RECT 0.310 39.120 118.370 43.840 ;
        RECT 2.800 37.720 117.200 39.120 ;
        RECT 0.310 33.680 118.370 37.720 ;
        RECT 0.310 32.280 117.200 33.680 ;
        RECT 0.310 30.280 118.370 32.280 ;
        RECT 2.800 28.880 118.370 30.280 ;
        RECT 0.310 27.560 118.370 28.880 ;
        RECT 0.310 26.160 117.200 27.560 ;
        RECT 0.310 22.120 118.370 26.160 ;
        RECT 2.800 21.440 118.370 22.120 ;
        RECT 2.800 20.720 117.200 21.440 ;
        RECT 0.310 20.040 117.200 20.720 ;
        RECT 0.310 15.320 118.370 20.040 ;
        RECT 0.310 13.920 117.200 15.320 ;
        RECT 0.310 13.280 118.370 13.920 ;
        RECT 2.800 11.880 118.370 13.280 ;
        RECT 0.310 9.200 118.370 11.880 ;
        RECT 0.310 7.800 117.200 9.200 ;
        RECT 0.310 5.120 118.370 7.800 ;
        RECT 2.800 3.760 118.370 5.120 ;
        RECT 2.800 3.720 117.200 3.760 ;
        RECT 0.310 3.360 117.200 3.720 ;
      LAYER met4 ;
        RECT 64.720 10.640 106.320 109.040 ;
  END
END decoder6to61
END LIBRARY

