VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__2_
  CLASS BLOCK ;
  FOREIGN cbx_1__2_ ;
  ORIGIN 0.000 -0.005 ;
  SIZE 150.000 BY 119.845 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 117.450 56.030 119.850 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 117.450 93.750 119.850 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.090 2.400 61.690 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.010 2.400 91.610 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.730 2.400 94.330 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.450 2.400 97.050 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.850 2.400 100.450 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.570 2.400 103.170 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.970 2.400 106.570 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.690 2.400 109.290 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.410 2.400 112.010 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.810 2.400 115.410 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.530 2.400 118.130 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.810 2.400 64.410 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.530 2.400 67.130 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.930 2.400 70.530 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.650 2.400 73.250 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.050 2.400 76.650 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.770 2.400 79.370 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.490 2.400 82.090 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.890 2.400 85.490 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.610 2.400 88.210 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.250 2.400 1.850 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.170 2.400 31.770 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.890 2.400 34.490 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.610 2.400 37.210 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.010 2.400 40.610 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.730 2.400 43.330 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.130 2.400 46.730 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.850 2.400 49.450 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.570 2.400 52.170 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.970 2.400 55.570 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.690 2.400 58.290 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.970 2.400 4.570 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.690 2.400 7.290 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.090 2.400 10.690 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.810 2.400 13.410 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.210 2.400 16.810 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.930 2.400 19.530 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.650 2.400 22.250 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.050 2.400 25.650 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.770 2.400 28.370 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 61.090 150.000 61.690 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 91.010 150.000 91.610 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 93.730 150.000 94.330 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 96.450 150.000 97.050 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 99.850 150.000 100.450 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 102.570 150.000 103.170 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 105.970 150.000 106.570 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 108.690 150.000 109.290 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 111.410 150.000 112.010 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 114.810 150.000 115.410 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 117.530 150.000 118.130 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 63.810 150.000 64.410 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 66.530 150.000 67.130 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 69.930 150.000 70.530 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 72.650 150.000 73.250 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 76.050 150.000 76.650 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 78.770 150.000 79.370 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 81.490 150.000 82.090 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 84.890 150.000 85.490 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 87.610 150.000 88.210 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 1.250 150.000 1.850 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 31.170 150.000 31.770 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 33.890 150.000 34.490 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 36.610 150.000 37.210 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 40.010 150.000 40.610 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 42.730 150.000 43.330 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 46.130 150.000 46.730 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 48.850 150.000 49.450 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 51.570 150.000 52.170 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 54.970 150.000 55.570 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 57.690 150.000 58.290 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 3.970 150.000 4.570 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 6.690 150.000 7.290 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 10.090 150.000 10.690 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 12.810 150.000 13.410 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 16.210 150.000 16.810 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 18.930 150.000 19.530 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 21.650 150.000 22.250 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 25.050 150.000 25.650 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 27.770 150.000 28.370 ;
    END
  END chanx_right_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 117.450 18.770 119.850 ;
    END
  END prog_clk
  PIN top_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 117.450 131.010 119.850 ;
    END
  END top_grid_pin_0_
  PIN vpwr
    USE POWER ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 29.720 10.490 31.320 108.890 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 54.720 10.490 56.320 108.890 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.645 144.440 108.735 ;
      LAYER met1 ;
        RECT 5.520 10.490 144.440 108.890 ;
      LAYER met2 ;
        RECT 6.530 117.170 18.210 118.015 ;
        RECT 19.050 117.170 55.470 118.015 ;
        RECT 56.310 117.170 93.190 118.015 ;
        RECT 94.030 117.170 130.450 118.015 ;
        RECT 6.530 0.005 131.260 117.170 ;
      LAYER met3 ;
        RECT 2.800 117.130 147.200 117.995 ;
        RECT 2.400 115.810 147.600 117.130 ;
        RECT 2.800 114.410 147.200 115.810 ;
        RECT 2.400 112.410 147.600 114.410 ;
        RECT 2.800 111.010 147.200 112.410 ;
        RECT 2.400 109.690 147.600 111.010 ;
        RECT 2.800 108.290 147.200 109.690 ;
        RECT 2.400 106.970 147.600 108.290 ;
        RECT 2.800 105.570 147.200 106.970 ;
        RECT 2.400 103.570 147.600 105.570 ;
        RECT 2.800 102.170 147.200 103.570 ;
        RECT 2.400 100.850 147.600 102.170 ;
        RECT 2.800 99.450 147.200 100.850 ;
        RECT 2.400 97.450 147.600 99.450 ;
        RECT 2.800 96.050 147.200 97.450 ;
        RECT 2.400 94.730 147.600 96.050 ;
        RECT 2.800 93.330 147.200 94.730 ;
        RECT 2.400 92.010 147.600 93.330 ;
        RECT 2.800 90.610 147.200 92.010 ;
        RECT 2.400 88.610 147.600 90.610 ;
        RECT 2.800 87.210 147.200 88.610 ;
        RECT 2.400 85.890 147.600 87.210 ;
        RECT 2.800 84.490 147.200 85.890 ;
        RECT 2.400 82.490 147.600 84.490 ;
        RECT 2.800 81.090 147.200 82.490 ;
        RECT 2.400 79.770 147.600 81.090 ;
        RECT 2.800 78.370 147.200 79.770 ;
        RECT 2.400 77.050 147.600 78.370 ;
        RECT 2.800 75.650 147.200 77.050 ;
        RECT 2.400 73.650 147.600 75.650 ;
        RECT 2.800 72.250 147.200 73.650 ;
        RECT 2.400 70.930 147.600 72.250 ;
        RECT 2.800 69.530 147.200 70.930 ;
        RECT 2.400 67.530 147.600 69.530 ;
        RECT 2.800 66.130 147.200 67.530 ;
        RECT 2.400 64.810 147.600 66.130 ;
        RECT 2.800 63.410 147.200 64.810 ;
        RECT 2.400 62.090 147.600 63.410 ;
        RECT 2.800 60.690 147.200 62.090 ;
        RECT 2.400 58.690 147.600 60.690 ;
        RECT 2.800 57.290 147.200 58.690 ;
        RECT 2.400 55.970 147.600 57.290 ;
        RECT 2.800 54.570 147.200 55.970 ;
        RECT 2.400 52.570 147.600 54.570 ;
        RECT 2.800 51.170 147.200 52.570 ;
        RECT 2.400 49.850 147.600 51.170 ;
        RECT 2.800 48.450 147.200 49.850 ;
        RECT 2.400 47.130 147.600 48.450 ;
        RECT 2.800 45.730 147.200 47.130 ;
        RECT 2.400 43.730 147.600 45.730 ;
        RECT 2.800 42.330 147.200 43.730 ;
        RECT 2.400 41.010 147.600 42.330 ;
        RECT 2.800 39.610 147.200 41.010 ;
        RECT 2.400 37.610 147.600 39.610 ;
        RECT 2.800 36.210 147.200 37.610 ;
        RECT 2.400 34.890 147.600 36.210 ;
        RECT 2.800 33.490 147.200 34.890 ;
        RECT 2.400 32.170 147.600 33.490 ;
        RECT 2.800 30.770 147.200 32.170 ;
        RECT 2.400 28.770 147.600 30.770 ;
        RECT 2.800 27.370 147.200 28.770 ;
        RECT 2.400 26.050 147.600 27.370 ;
        RECT 2.800 24.650 147.200 26.050 ;
        RECT 2.400 22.650 147.600 24.650 ;
        RECT 2.800 21.250 147.200 22.650 ;
        RECT 2.400 19.930 147.600 21.250 ;
        RECT 2.800 18.530 147.200 19.930 ;
        RECT 2.400 17.210 147.600 18.530 ;
        RECT 2.800 15.810 147.200 17.210 ;
        RECT 2.400 13.810 147.600 15.810 ;
        RECT 2.800 12.410 147.200 13.810 ;
        RECT 2.400 11.090 147.600 12.410 ;
        RECT 2.800 9.690 147.200 11.090 ;
        RECT 2.400 7.690 147.600 9.690 ;
        RECT 2.800 6.290 147.200 7.690 ;
        RECT 2.400 4.970 147.600 6.290 ;
        RECT 2.800 3.570 147.200 4.970 ;
        RECT 2.400 2.250 147.600 3.570 ;
        RECT 2.800 0.850 147.200 2.250 ;
        RECT 2.400 0.025 147.600 0.850 ;
      LAYER met4 ;
        RECT 16.430 10.090 29.320 108.890 ;
        RECT 31.720 10.090 54.320 108.890 ;
        RECT 56.720 10.090 131.320 108.890 ;
        RECT 16.430 0.025 131.320 10.090 ;
      LAYER met5 ;
        RECT 16.220 58.550 125.460 60.150 ;
  END
END cbx_1__2_
END LIBRARY

