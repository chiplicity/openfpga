magic
tech sky130A
magscale 1 2
timestamp 1605203969
<< locali >>
rect 6561 6715 6595 6817
<< viali >>
rect 8769 13481 8803 13515
rect 11529 13481 11563 13515
rect 7389 13413 7423 13447
rect 2145 13345 2179 13379
rect 4077 13345 4111 13379
rect 5181 13345 5215 13379
rect 7481 13345 7515 13379
rect 8585 13345 8619 13379
rect 10149 13345 10183 13379
rect 11345 13345 11379 13379
rect 7573 13277 7607 13311
rect 10241 13277 10275 13311
rect 10333 13277 10367 13311
rect 7021 13209 7055 13243
rect 2329 13141 2363 13175
rect 4261 13141 4295 13175
rect 5365 13141 5399 13175
rect 9781 13141 9815 13175
rect 4537 12937 4571 12971
rect 7021 12937 7055 12971
rect 8585 12937 8619 12971
rect 3433 12869 3467 12903
rect 11437 12869 11471 12903
rect 12633 12869 12667 12903
rect 2145 12733 2179 12767
rect 3249 12733 3283 12767
rect 4353 12733 4387 12767
rect 5457 12733 5491 12767
rect 6837 12733 6871 12767
rect 8401 12733 8435 12767
rect 10149 12733 10183 12767
rect 11253 12733 11287 12767
rect 12449 12733 12483 12767
rect 13553 12665 13587 12699
rect 2329 12597 2363 12631
rect 5641 12597 5675 12631
rect 10333 12597 10367 12631
rect 6929 12393 6963 12427
rect 7297 12393 7331 12427
rect 9873 12393 9907 12427
rect 13645 12393 13679 12427
rect 2145 12257 2179 12291
rect 4077 12257 4111 12291
rect 5181 12257 5215 12291
rect 8493 12257 8527 12291
rect 9695 12257 9729 12291
rect 11253 12257 11287 12291
rect 12357 12257 12391 12291
rect 13461 12257 13495 12291
rect 7389 12189 7423 12223
rect 7573 12189 7607 12223
rect 8677 12121 8711 12155
rect 12541 12121 12575 12155
rect 2329 12053 2363 12087
rect 4261 12053 4295 12087
rect 5365 12053 5399 12087
rect 11437 12053 11471 12087
rect 5917 11849 5951 11883
rect 8401 11849 8435 11883
rect 10793 11781 10827 11815
rect 3617 11713 3651 11747
rect 7481 11713 7515 11747
rect 9045 11713 9079 11747
rect 11437 11713 11471 11747
rect 13001 11713 13035 11747
rect 1961 11645 1995 11679
rect 4629 11645 4663 11679
rect 7205 11645 7239 11679
rect 8861 11645 8895 11679
rect 11161 11645 11195 11679
rect 12909 11645 12943 11679
rect 3433 11577 3467 11611
rect 12817 11577 12851 11611
rect 2145 11509 2179 11543
rect 3065 11509 3099 11543
rect 3525 11509 3559 11543
rect 4813 11509 4847 11543
rect 6837 11509 6871 11543
rect 7297 11509 7331 11543
rect 8769 11509 8803 11543
rect 11253 11509 11287 11543
rect 12449 11509 12483 11543
rect 2145 11305 2179 11339
rect 4445 11305 4479 11339
rect 8401 11305 8435 11339
rect 4537 11237 4571 11271
rect 2513 11169 2547 11203
rect 5641 11169 5675 11203
rect 9945 11169 9979 11203
rect 13369 11169 13403 11203
rect 2605 11101 2639 11135
rect 2697 11101 2731 11135
rect 4721 11101 4755 11135
rect 7021 11101 7055 11135
rect 8493 11101 8527 11135
rect 8585 11101 8619 11135
rect 9689 11101 9723 11135
rect 11897 11101 11931 11135
rect 4077 11033 4111 11067
rect 5825 11033 5859 11067
rect 8033 11033 8067 11067
rect 11069 11033 11103 11067
rect 13553 11033 13587 11067
rect 8493 10761 8527 10795
rect 12817 10761 12851 10795
rect 11437 10693 11471 10727
rect 7481 10625 7515 10659
rect 8953 10625 8987 10659
rect 9045 10625 9079 10659
rect 13369 10625 13403 10659
rect 1777 10557 1811 10591
rect 2881 10557 2915 10591
rect 3148 10557 3182 10591
rect 5089 10557 5123 10591
rect 10057 10557 10091 10591
rect 11253 10557 11287 10591
rect 7389 10489 7423 10523
rect 13277 10489 13311 10523
rect 1961 10421 1995 10455
rect 4261 10421 4295 10455
rect 5273 10421 5307 10455
rect 6929 10421 6963 10455
rect 7297 10421 7331 10455
rect 8861 10421 8895 10455
rect 10241 10421 10275 10455
rect 13185 10421 13219 10455
rect 3157 10217 3191 10251
rect 8585 10217 8619 10251
rect 4966 10149 5000 10183
rect 1777 10081 1811 10115
rect 2044 10081 2078 10115
rect 7472 10081 7506 10115
rect 9965 10081 9999 10115
rect 11069 10081 11103 10115
rect 11336 10081 11370 10115
rect 13369 10081 13403 10115
rect 4721 10013 4755 10047
rect 7205 10013 7239 10047
rect 6101 9945 6135 9979
rect 13553 9945 13587 9979
rect 10149 9877 10183 9911
rect 12449 9877 12483 9911
rect 2237 9605 2271 9639
rect 9321 9605 9355 9639
rect 2789 9537 2823 9571
rect 7941 9537 7975 9571
rect 10149 9537 10183 9571
rect 12909 9537 12943 9571
rect 13001 9537 13035 9571
rect 2605 9469 2639 9503
rect 2697 9469 2731 9503
rect 3893 9469 3927 9503
rect 6837 9469 6871 9503
rect 8208 9469 8242 9503
rect 12817 9469 12851 9503
rect 4138 9401 4172 9435
rect 10416 9401 10450 9435
rect 5273 9333 5307 9367
rect 7021 9333 7055 9367
rect 11529 9333 11563 9367
rect 12449 9333 12483 9367
rect 2881 9129 2915 9163
rect 4077 9129 4111 9163
rect 4537 9129 4571 9163
rect 5641 9129 5675 9163
rect 6009 9129 6043 9163
rect 7665 9129 7699 9163
rect 12725 9129 12759 9163
rect 10416 9061 10450 9095
rect 2789 8993 2823 9027
rect 4445 8993 4479 9027
rect 6101 8993 6135 9027
rect 7573 8993 7607 9027
rect 8953 8993 8987 9027
rect 10149 8993 10183 9027
rect 1409 8925 1443 8959
rect 3065 8925 3099 8959
rect 4629 8925 4663 8959
rect 6193 8925 6227 8959
rect 7757 8925 7791 8959
rect 12817 8925 12851 8959
rect 12909 8925 12943 8959
rect 11529 8857 11563 8891
rect 2421 8789 2455 8823
rect 7205 8789 7239 8823
rect 8769 8789 8803 8823
rect 12357 8789 12391 8823
rect 2145 8585 2179 8619
rect 3801 8585 3835 8619
rect 10793 8585 10827 8619
rect 12449 8585 12483 8619
rect 5365 8517 5399 8551
rect 5825 8517 5859 8551
rect 6837 8517 6871 8551
rect 2697 8449 2731 8483
rect 4353 8449 4387 8483
rect 7481 8449 7515 8483
rect 8953 8449 8987 8483
rect 11345 8449 11379 8483
rect 12909 8449 12943 8483
rect 13001 8449 13035 8483
rect 2513 8381 2547 8415
rect 2605 8381 2639 8415
rect 5549 8381 5583 8415
rect 5641 8381 5675 8415
rect 7205 8381 7239 8415
rect 10149 8381 10183 8415
rect 12817 8381 12851 8415
rect 8769 8313 8803 8347
rect 8861 8313 8895 8347
rect 11161 8313 11195 8347
rect 11253 8313 11287 8347
rect 4169 8245 4203 8279
rect 4261 8245 4295 8279
rect 7297 8245 7331 8279
rect 8401 8245 8435 8279
rect 9965 8245 9999 8279
rect 5457 8041 5491 8075
rect 7297 8041 7331 8075
rect 2789 7973 2823 8007
rect 11428 7973 11462 8007
rect 4333 7905 4367 7939
rect 8493 7905 8527 7939
rect 10057 7905 10091 7939
rect 11161 7905 11195 7939
rect 13369 7905 13403 7939
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 4077 7837 4111 7871
rect 7389 7837 7423 7871
rect 7573 7837 7607 7871
rect 8677 7769 8711 7803
rect 2421 7701 2455 7735
rect 6929 7701 6963 7735
rect 10241 7701 10275 7735
rect 12541 7701 12575 7735
rect 13553 7701 13587 7735
rect 3709 7497 3743 7531
rect 4537 7497 4571 7531
rect 7665 7497 7699 7531
rect 12449 7497 12483 7531
rect 4997 7361 5031 7395
rect 5181 7361 5215 7395
rect 8217 7361 8251 7395
rect 10885 7361 10919 7395
rect 13093 7361 13127 7395
rect 2329 7293 2363 7327
rect 8033 7293 8067 7327
rect 9229 7293 9263 7327
rect 10701 7293 10735 7327
rect 2596 7225 2630 7259
rect 10793 7225 10827 7259
rect 12817 7225 12851 7259
rect 4905 7157 4939 7191
rect 8125 7157 8159 7191
rect 9413 7157 9447 7191
rect 10333 7157 10367 7191
rect 12909 7157 12943 7191
rect 8861 6953 8895 6987
rect 13553 6953 13587 6987
rect 2789 6885 2823 6919
rect 8217 6885 8251 6919
rect 12440 6885 12474 6919
rect 1409 6817 1443 6851
rect 4077 6817 4111 6851
rect 5365 6817 5399 6851
rect 6561 6817 6595 6851
rect 6653 6817 6687 6851
rect 10232 6817 10266 6851
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 9965 6749 9999 6783
rect 12173 6749 12207 6783
rect 6561 6681 6595 6715
rect 11345 6681 11379 6715
rect 2421 6613 2455 6647
rect 4261 6613 4295 6647
rect 5181 6613 5215 6647
rect 8493 6613 8527 6647
rect 3801 6409 3835 6443
rect 6653 6409 6687 6443
rect 10885 6409 10919 6443
rect 12633 6409 12667 6443
rect 4445 6341 4479 6375
rect 2421 6273 2455 6307
rect 4997 6273 5031 6307
rect 5273 6273 5307 6307
rect 9505 6273 9539 6307
rect 13185 6273 13219 6307
rect 4905 6205 4939 6239
rect 7297 6205 7331 6239
rect 13093 6205 13127 6239
rect 2688 6137 2722 6171
rect 5540 6137 5574 6171
rect 7564 6137 7598 6171
rect 9772 6137 9806 6171
rect 13001 6137 13035 6171
rect 1409 6069 1443 6103
rect 4813 6069 4847 6103
rect 8677 6069 8711 6103
rect 8401 5865 8435 5899
rect 11069 5865 11103 5899
rect 12633 5865 12667 5899
rect 2789 5797 2823 5831
rect 5632 5797 5666 5831
rect 8493 5797 8527 5831
rect 13001 5797 13035 5831
rect 1409 5729 1443 5763
rect 1777 5729 1811 5763
rect 4077 5729 4111 5763
rect 9956 5729 9990 5763
rect 2881 5661 2915 5695
rect 2973 5661 3007 5695
rect 5365 5661 5399 5695
rect 8677 5661 8711 5695
rect 9689 5661 9723 5695
rect 13093 5661 13127 5695
rect 13185 5661 13219 5695
rect 1961 5593 1995 5627
rect 2329 5593 2363 5627
rect 1593 5525 1627 5559
rect 2421 5525 2455 5559
rect 4261 5525 4295 5559
rect 6745 5525 6779 5559
rect 8033 5525 8067 5559
rect 1409 5321 1443 5355
rect 3341 5321 3375 5355
rect 4905 5321 4939 5355
rect 6469 5321 6503 5355
rect 9597 5321 9631 5355
rect 9965 5321 9999 5355
rect 7113 5253 7147 5287
rect 1961 5185 1995 5219
rect 2881 5185 2915 5219
rect 3801 5185 3835 5219
rect 3985 5185 4019 5219
rect 5457 5185 5491 5219
rect 8493 5185 8527 5219
rect 8677 5185 8711 5219
rect 10609 5185 10643 5219
rect 13185 5185 13219 5219
rect 1777 5117 1811 5151
rect 5273 5117 5307 5151
rect 6653 5117 6687 5151
rect 6929 5117 6963 5151
rect 9781 5117 9815 5151
rect 10425 5117 10459 5151
rect 12909 5117 12943 5151
rect 3709 5049 3743 5083
rect 8401 5049 8435 5083
rect 13001 5049 13035 5083
rect 1869 4981 1903 5015
rect 2237 4981 2271 5015
rect 2605 4981 2639 5015
rect 2697 4981 2731 5015
rect 5365 4981 5399 5015
rect 8033 4981 8067 5015
rect 10333 4981 10367 5015
rect 12541 4981 12575 5015
rect 1409 4777 1443 4811
rect 2789 4777 2823 4811
rect 5457 4777 5491 4811
rect 7757 4777 7791 4811
rect 7849 4777 7883 4811
rect 10333 4777 10367 4811
rect 10701 4777 10735 4811
rect 12081 4777 12115 4811
rect 12541 4777 12575 4811
rect 4322 4709 4356 4743
rect 1777 4641 1811 4675
rect 1869 4641 1903 4675
rect 3249 4641 3283 4675
rect 6285 4641 6319 4675
rect 12449 4641 12483 4675
rect 2053 4573 2087 4607
rect 2881 4573 2915 4607
rect 3065 4573 3099 4607
rect 3433 4573 3467 4607
rect 4077 4573 4111 4607
rect 7941 4573 7975 4607
rect 10793 4573 10827 4607
rect 10977 4573 11011 4607
rect 12633 4573 12667 4607
rect 6469 4505 6503 4539
rect 2421 4437 2455 4471
rect 7389 4437 7423 4471
rect 13553 4233 13587 4267
rect 2237 4165 2271 4199
rect 1961 4097 1995 4131
rect 2697 4097 2731 4131
rect 2789 4097 2823 4131
rect 4261 4097 4295 4131
rect 7297 4097 7331 4131
rect 7481 4097 7515 4131
rect 8401 4097 8435 4131
rect 3065 4029 3099 4063
rect 4169 4029 4203 4063
rect 4537 4029 4571 4063
rect 5457 4029 5491 4063
rect 8668 4029 8702 4063
rect 11253 4029 11287 4063
rect 13369 4029 13403 4063
rect 1777 3961 1811 3995
rect 3341 3961 3375 3995
rect 5733 3961 5767 3995
rect 7205 3961 7239 3995
rect 1409 3893 1443 3927
rect 1869 3893 1903 3927
rect 2605 3893 2639 3927
rect 3709 3893 3743 3927
rect 4077 3893 4111 3927
rect 4721 3893 4755 3927
rect 6837 3893 6871 3927
rect 9781 3893 9815 3927
rect 11437 3893 11471 3927
rect 2881 3689 2915 3723
rect 3249 3689 3283 3723
rect 5457 3689 5491 3723
rect 12449 3689 12483 3723
rect 13553 3689 13587 3723
rect 1676 3621 1710 3655
rect 4445 3621 4479 3655
rect 4537 3621 4571 3655
rect 7012 3621 7046 3655
rect 9965 3621 9999 3655
rect 3341 3553 3375 3587
rect 4905 3553 4939 3587
rect 5273 3553 5307 3587
rect 5641 3553 5675 3587
rect 6745 3553 6779 3587
rect 9689 3553 9723 3587
rect 11161 3553 11195 3587
rect 12265 3553 12299 3587
rect 13369 3553 13403 3587
rect 3525 3485 3559 3519
rect 4629 3485 4663 3519
rect 2789 3417 2823 3451
rect 4077 3417 4111 3451
rect 5089 3349 5123 3383
rect 5825 3349 5859 3383
rect 8125 3349 8159 3383
rect 11345 3349 11379 3383
rect 13553 3145 13587 3179
rect 4353 3077 4387 3111
rect 9229 3077 9263 3111
rect 4905 3009 4939 3043
rect 1676 2941 1710 2975
rect 2881 2941 2915 2975
rect 5181 2941 5215 2975
rect 5733 2941 5767 2975
rect 6837 2941 6871 2975
rect 7941 2941 7975 2975
rect 9045 2941 9079 2975
rect 10149 2941 10183 2975
rect 11253 2941 11287 2975
rect 13369 2941 13403 2975
rect 3148 2873 3182 2907
rect 4813 2873 4847 2907
rect 5457 2873 5491 2907
rect 2789 2805 2823 2839
rect 4261 2805 4295 2839
rect 4721 2805 4755 2839
rect 5917 2805 5951 2839
rect 7021 2805 7055 2839
rect 8125 2805 8159 2839
rect 10333 2805 10367 2839
rect 11437 2805 11471 2839
rect 8309 2601 8343 2635
rect 13553 2601 13587 2635
rect 1676 2533 1710 2567
rect 4353 2533 4387 2567
rect 7196 2533 7230 2567
rect 1409 2465 1443 2499
rect 3249 2465 3283 2499
rect 4077 2465 4111 2499
rect 4885 2465 4919 2499
rect 6101 2465 6135 2499
rect 6469 2465 6503 2499
rect 6929 2465 6963 2499
rect 9781 2465 9815 2499
rect 11437 2465 11471 2499
rect 13369 2465 13403 2499
rect 3341 2397 3375 2431
rect 3525 2397 3559 2431
rect 4629 2397 4663 2431
rect 2789 2329 2823 2363
rect 6009 2329 6043 2363
rect 2881 2261 2915 2295
rect 6285 2261 6319 2295
rect 6653 2261 6687 2295
rect 9965 2261 9999 2295
rect 11621 2261 11655 2295
<< metal1 >>
rect 3326 15036 3332 15088
rect 3384 15076 3390 15088
rect 6822 15076 6828 15088
rect 3384 15048 6828 15076
rect 3384 15036 3390 15048
rect 6822 15036 6828 15048
rect 6880 15036 6886 15088
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 7282 14260 7288 14272
rect 2832 14232 7288 14260
rect 2832 14220 2838 14232
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 4062 14152 4068 14204
rect 4120 14192 4126 14204
rect 6914 14192 6920 14204
rect 4120 14164 6920 14192
rect 4120 14152 4126 14164
rect 6914 14152 6920 14164
rect 6972 14152 6978 14204
rect 4338 14016 4344 14068
rect 4396 14056 4402 14068
rect 8478 14056 8484 14068
rect 4396 14028 8484 14056
rect 4396 14016 4402 14028
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 5074 13948 5080 14000
rect 5132 13988 5138 14000
rect 11238 13988 11244 14000
rect 5132 13960 11244 13988
rect 5132 13948 5138 13960
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 5258 13880 5264 13932
rect 5316 13920 5322 13932
rect 11054 13920 11060 13932
rect 5316 13892 11060 13920
rect 5316 13880 5322 13892
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 5442 13852 5448 13864
rect 4120 13824 5448 13852
rect 4120 13812 4126 13824
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 7742 13852 7748 13864
rect 7116 13824 7748 13852
rect 4798 13744 4804 13796
rect 4856 13784 4862 13796
rect 7116 13784 7144 13824
rect 7742 13812 7748 13824
rect 7800 13852 7806 13864
rect 11146 13852 11152 13864
rect 7800 13824 11152 13852
rect 7800 13812 7806 13824
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 4856 13756 7144 13784
rect 4856 13744 4862 13756
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 6178 13716 6184 13728
rect 2004 13688 6184 13716
rect 2004 13676 2010 13688
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 1104 13626 14812 13648
rect 1104 13574 5579 13626
rect 5631 13574 5643 13626
rect 5695 13574 5707 13626
rect 5759 13574 5771 13626
rect 5823 13574 10176 13626
rect 10228 13574 10240 13626
rect 10292 13574 10304 13626
rect 10356 13574 10368 13626
rect 10420 13574 14812 13626
rect 1104 13552 14812 13574
rect 1118 13472 1124 13524
rect 1176 13512 1182 13524
rect 8757 13515 8815 13521
rect 8757 13512 8769 13515
rect 1176 13484 8769 13512
rect 1176 13472 1182 13484
rect 8757 13481 8769 13484
rect 8803 13481 8815 13515
rect 11514 13512 11520 13524
rect 11475 13484 11520 13512
rect 8757 13475 8815 13481
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 3050 13404 3056 13456
rect 3108 13444 3114 13456
rect 7377 13447 7435 13453
rect 7377 13444 7389 13447
rect 3108 13416 7389 13444
rect 3108 13404 3114 13416
rect 7377 13413 7389 13416
rect 7423 13444 7435 13447
rect 8202 13444 8208 13456
rect 7423 13416 8208 13444
rect 7423 13413 7435 13416
rect 7377 13407 7435 13413
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 10594 13444 10600 13456
rect 8588 13416 10600 13444
rect 2133 13379 2191 13385
rect 2133 13345 2145 13379
rect 2179 13345 2191 13379
rect 2133 13339 2191 13345
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 4798 13376 4804 13388
rect 4111 13348 4804 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 2148 13240 2176 13339
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 4890 13336 4896 13388
rect 4948 13376 4954 13388
rect 5169 13379 5227 13385
rect 5169 13376 5181 13379
rect 4948 13348 5181 13376
rect 4948 13336 4954 13348
rect 5169 13345 5181 13348
rect 5215 13376 5227 13379
rect 5258 13376 5264 13388
rect 5215 13348 5264 13376
rect 5215 13345 5227 13348
rect 5169 13339 5227 13345
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 8588 13385 8616 13416
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7156 13348 7481 13376
rect 7156 13336 7162 13348
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 8573 13379 8631 13385
rect 8573 13345 8585 13379
rect 8619 13345 8631 13379
rect 8573 13339 8631 13345
rect 9122 13336 9128 13388
rect 9180 13376 9186 13388
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 9180 13348 10149 13376
rect 9180 13336 9186 13348
rect 10137 13345 10149 13348
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 10560 13348 11345 13376
rect 10560 13336 10566 13348
rect 11333 13345 11345 13348
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 7558 13308 7564 13320
rect 7519 13280 7564 13308
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 9272 13280 10241 13308
rect 9272 13268 9278 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 7009 13243 7067 13249
rect 2148 13212 6960 13240
rect 1670 13132 1676 13184
rect 1728 13172 1734 13184
rect 2317 13175 2375 13181
rect 2317 13172 2329 13175
rect 1728 13144 2329 13172
rect 1728 13132 1734 13144
rect 2317 13141 2329 13144
rect 2363 13141 2375 13175
rect 2317 13135 2375 13141
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 4212 13144 4261 13172
rect 4212 13132 4218 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 5350 13172 5356 13184
rect 5311 13144 5356 13172
rect 4249 13135 4307 13141
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 6932 13172 6960 13212
rect 7009 13209 7021 13243
rect 7055 13240 7067 13243
rect 8846 13240 8852 13252
rect 7055 13212 8852 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 8846 13200 8852 13212
rect 8904 13200 8910 13252
rect 10042 13200 10048 13252
rect 10100 13240 10106 13252
rect 10336 13240 10364 13271
rect 10100 13212 10364 13240
rect 10100 13200 10106 13212
rect 7374 13172 7380 13184
rect 6932 13144 7380 13172
rect 7374 13132 7380 13144
rect 7432 13172 7438 13184
rect 9306 13172 9312 13184
rect 7432 13144 9312 13172
rect 7432 13132 7438 13144
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 9766 13172 9772 13184
rect 9727 13144 9772 13172
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 1104 13082 14812 13104
rect 1104 13030 3280 13082
rect 3332 13030 3344 13082
rect 3396 13030 3408 13082
rect 3460 13030 3472 13082
rect 3524 13030 7878 13082
rect 7930 13030 7942 13082
rect 7994 13030 8006 13082
rect 8058 13030 8070 13082
rect 8122 13030 12475 13082
rect 12527 13030 12539 13082
rect 12591 13030 12603 13082
rect 12655 13030 12667 13082
rect 12719 13030 14812 13082
rect 1104 13008 14812 13030
rect 2038 12928 2044 12980
rect 2096 12968 2102 12980
rect 4525 12971 4583 12977
rect 4525 12968 4537 12971
rect 2096 12940 4537 12968
rect 2096 12928 2102 12940
rect 4525 12937 4537 12940
rect 4571 12937 4583 12971
rect 4525 12931 4583 12937
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 7009 12971 7067 12977
rect 7009 12968 7021 12971
rect 5224 12940 7021 12968
rect 5224 12928 5230 12940
rect 7009 12937 7021 12940
rect 7055 12937 7067 12971
rect 7009 12931 7067 12937
rect 8573 12971 8631 12977
rect 8573 12937 8585 12971
rect 8619 12968 8631 12971
rect 13538 12968 13544 12980
rect 8619 12940 13544 12968
rect 8619 12937 8631 12940
rect 8573 12931 8631 12937
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 2498 12860 2504 12912
rect 2556 12900 2562 12912
rect 3421 12903 3479 12909
rect 3421 12900 3433 12903
rect 2556 12872 3433 12900
rect 2556 12860 2562 12872
rect 3421 12869 3433 12872
rect 3467 12869 3479 12903
rect 3421 12863 3479 12869
rect 4356 12872 6040 12900
rect 2130 12764 2136 12776
rect 2091 12736 2136 12764
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 3234 12764 3240 12776
rect 3195 12736 3240 12764
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 3694 12724 3700 12776
rect 3752 12764 3758 12776
rect 4356 12773 4384 12872
rect 4341 12767 4399 12773
rect 3752 12736 4292 12764
rect 3752 12724 3758 12736
rect 4264 12696 4292 12736
rect 4341 12733 4353 12767
rect 4387 12733 4399 12767
rect 4341 12727 4399 12733
rect 5445 12767 5503 12773
rect 5445 12733 5457 12767
rect 5491 12733 5503 12767
rect 6012 12764 6040 12872
rect 7282 12860 7288 12912
rect 7340 12900 7346 12912
rect 11425 12903 11483 12909
rect 11425 12900 11437 12903
rect 7340 12872 11437 12900
rect 7340 12860 7346 12872
rect 11425 12869 11437 12872
rect 11471 12869 11483 12903
rect 11425 12863 11483 12869
rect 12621 12903 12679 12909
rect 12621 12869 12633 12903
rect 12667 12869 12679 12903
rect 12621 12863 12679 12869
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 11054 12832 11060 12844
rect 6144 12804 11060 12832
rect 6144 12792 6150 12804
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 12636 12832 12664 12863
rect 11164 12804 12664 12832
rect 6825 12767 6883 12773
rect 6012 12736 6684 12764
rect 5445 12727 5503 12733
rect 4264 12668 4936 12696
rect 2317 12631 2375 12637
rect 2317 12597 2329 12631
rect 2363 12628 2375 12631
rect 2866 12628 2872 12640
rect 2363 12600 2872 12628
rect 2363 12597 2375 12600
rect 2317 12591 2375 12597
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 4430 12628 4436 12640
rect 3568 12600 4436 12628
rect 3568 12588 3574 12600
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 4908 12628 4936 12668
rect 5074 12628 5080 12640
rect 4908 12600 5080 12628
rect 5074 12588 5080 12600
rect 5132 12628 5138 12640
rect 5460 12628 5488 12727
rect 6656 12696 6684 12736
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 7006 12764 7012 12776
rect 6871 12736 7012 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 7708 12736 8401 12764
rect 7708 12724 7714 12736
rect 8389 12733 8401 12736
rect 8435 12733 8447 12767
rect 8389 12727 8447 12733
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 9732 12736 10149 12764
rect 9732 12724 9738 12736
rect 10137 12733 10149 12736
rect 10183 12733 10195 12767
rect 11164 12764 11192 12804
rect 10137 12727 10195 12733
rect 10244 12736 11192 12764
rect 11241 12767 11299 12773
rect 9858 12696 9864 12708
rect 6656 12668 9864 12696
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 5132 12600 5488 12628
rect 5629 12631 5687 12637
rect 5132 12588 5138 12600
rect 5629 12597 5641 12631
rect 5675 12628 5687 12631
rect 5994 12628 6000 12640
rect 5675 12600 6000 12628
rect 5675 12597 5687 12600
rect 5629 12591 5687 12597
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10244 12628 10272 12736
rect 11241 12733 11253 12767
rect 11287 12764 11299 12767
rect 11330 12764 11336 12776
rect 11287 12736 11336 12764
rect 11287 12733 11299 12736
rect 11241 12727 11299 12733
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 13078 12764 13084 12776
rect 12483 12736 13084 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 11146 12656 11152 12708
rect 11204 12696 11210 12708
rect 13541 12699 13599 12705
rect 13541 12696 13553 12699
rect 11204 12668 13553 12696
rect 11204 12656 11210 12668
rect 13541 12665 13553 12668
rect 13587 12665 13599 12699
rect 13541 12659 13599 12665
rect 9824 12600 10272 12628
rect 10321 12631 10379 12637
rect 9824 12588 9830 12600
rect 10321 12597 10333 12631
rect 10367 12628 10379 12631
rect 10962 12628 10968 12640
rect 10367 12600 10968 12628
rect 10367 12597 10379 12600
rect 10321 12591 10379 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 1104 12538 14812 12560
rect 1104 12486 5579 12538
rect 5631 12486 5643 12538
rect 5695 12486 5707 12538
rect 5759 12486 5771 12538
rect 5823 12486 10176 12538
rect 10228 12486 10240 12538
rect 10292 12486 10304 12538
rect 10356 12486 10368 12538
rect 10420 12486 14812 12538
rect 1104 12464 14812 12486
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 6638 12424 6644 12436
rect 3292 12396 6644 12424
rect 3292 12384 3298 12396
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 6917 12427 6975 12433
rect 6917 12393 6929 12427
rect 6963 12424 6975 12427
rect 7098 12424 7104 12436
rect 6963 12396 7104 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7285 12427 7343 12433
rect 7285 12424 7297 12427
rect 7208 12396 7297 12424
rect 7208 12368 7236 12396
rect 7285 12393 7297 12396
rect 7331 12393 7343 12427
rect 7285 12387 7343 12393
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 9766 12424 9772 12436
rect 8536 12396 9772 12424
rect 8536 12384 8542 12396
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 9861 12427 9919 12433
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 13633 12427 13691 12433
rect 9907 12396 13400 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 4982 12316 4988 12368
rect 5040 12356 5046 12368
rect 7006 12356 7012 12368
rect 5040 12328 7012 12356
rect 5040 12316 5046 12328
rect 7006 12316 7012 12328
rect 7064 12316 7070 12368
rect 7190 12316 7196 12368
rect 7248 12316 7254 12368
rect 8386 12316 8392 12368
rect 8444 12356 8450 12368
rect 8444 12328 9720 12356
rect 8444 12316 8450 12328
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2682 12288 2688 12300
rect 2179 12260 2688 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12288 4123 12291
rect 4246 12288 4252 12300
rect 4111 12260 4252 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 5166 12288 5172 12300
rect 5127 12260 5172 12288
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 8481 12291 8539 12297
rect 8481 12257 8493 12291
rect 8527 12288 8539 12291
rect 9030 12288 9036 12300
rect 8527 12260 9036 12288
rect 8527 12257 8539 12260
rect 8481 12251 8539 12257
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 9692 12297 9720 12328
rect 10686 12316 10692 12368
rect 10744 12356 10750 12368
rect 11422 12356 11428 12368
rect 10744 12328 11428 12356
rect 10744 12316 10750 12328
rect 11422 12316 11428 12328
rect 11480 12316 11486 12368
rect 11790 12316 11796 12368
rect 11848 12356 11854 12368
rect 11974 12356 11980 12368
rect 11848 12328 11980 12356
rect 11848 12316 11854 12328
rect 11974 12316 11980 12328
rect 12032 12316 12038 12368
rect 13372 12356 13400 12396
rect 13633 12393 13645 12427
rect 13679 12424 13691 12427
rect 14734 12424 14740 12436
rect 13679 12396 14740 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 14090 12356 14096 12368
rect 13372 12328 14096 12356
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 9683 12291 9741 12297
rect 9683 12257 9695 12291
rect 9729 12257 9741 12291
rect 9683 12251 9741 12257
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12257 11299 12291
rect 11241 12251 11299 12257
rect 382 12180 388 12232
rect 440 12220 446 12232
rect 440 12192 5764 12220
rect 440 12180 446 12192
rect 5736 12152 5764 12192
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 7156 12192 7389 12220
rect 7156 12180 7162 12192
rect 7377 12189 7389 12192
rect 7423 12189 7435 12223
rect 7558 12220 7564 12232
rect 7519 12192 7564 12220
rect 7377 12183 7435 12189
rect 7558 12180 7564 12192
rect 7616 12180 7622 12232
rect 11256 12220 11284 12251
rect 11330 12248 11336 12300
rect 11388 12288 11394 12300
rect 12345 12291 12403 12297
rect 12345 12288 12357 12291
rect 11388 12260 12357 12288
rect 11388 12248 11394 12260
rect 12345 12257 12357 12260
rect 12391 12257 12403 12291
rect 12345 12251 12403 12257
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 8772 12192 11284 12220
rect 8665 12155 8723 12161
rect 8665 12152 8677 12155
rect 5736 12124 8677 12152
rect 8665 12121 8677 12124
rect 8711 12121 8723 12155
rect 8665 12115 8723 12121
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 2317 12087 2375 12093
rect 2317 12084 2329 12087
rect 2096 12056 2329 12084
rect 2096 12044 2102 12056
rect 2317 12053 2329 12056
rect 2363 12053 2375 12087
rect 2317 12047 2375 12053
rect 2406 12044 2412 12096
rect 2464 12084 2470 12096
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 2464 12056 4261 12084
rect 2464 12044 2470 12056
rect 4249 12053 4261 12056
rect 4295 12053 4307 12087
rect 4249 12047 4307 12053
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5353 12087 5411 12093
rect 5353 12084 5365 12087
rect 4856 12056 5365 12084
rect 4856 12044 4862 12056
rect 5353 12053 5365 12056
rect 5399 12053 5411 12087
rect 5353 12047 5411 12053
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 8772 12084 8800 12192
rect 11974 12180 11980 12232
rect 12032 12220 12038 12232
rect 13464 12220 13492 12251
rect 12032 12192 13492 12220
rect 12032 12180 12038 12192
rect 8938 12112 8944 12164
rect 8996 12152 9002 12164
rect 9674 12152 9680 12164
rect 8996 12124 9680 12152
rect 8996 12112 9002 12124
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 12529 12155 12587 12161
rect 12529 12121 12541 12155
rect 12575 12152 12587 12155
rect 13906 12152 13912 12164
rect 12575 12124 13912 12152
rect 12575 12121 12587 12124
rect 12529 12115 12587 12121
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 6788 12056 8800 12084
rect 6788 12044 6794 12056
rect 9030 12044 9036 12096
rect 9088 12084 9094 12096
rect 10502 12084 10508 12096
rect 9088 12056 10508 12084
rect 9088 12044 9094 12056
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 11425 12087 11483 12093
rect 11425 12053 11437 12087
rect 11471 12084 11483 12087
rect 13446 12084 13452 12096
rect 11471 12056 13452 12084
rect 11471 12053 11483 12056
rect 11425 12047 11483 12053
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 1104 11994 14812 12016
rect 1104 11942 3280 11994
rect 3332 11942 3344 11994
rect 3396 11942 3408 11994
rect 3460 11942 3472 11994
rect 3524 11942 7878 11994
rect 7930 11942 7942 11994
rect 7994 11942 8006 11994
rect 8058 11942 8070 11994
rect 8122 11942 12475 11994
rect 12527 11942 12539 11994
rect 12591 11942 12603 11994
rect 12655 11942 12667 11994
rect 12719 11942 14812 11994
rect 1104 11920 14812 11942
rect 3602 11840 3608 11892
rect 3660 11880 3666 11892
rect 4522 11880 4528 11892
rect 3660 11852 4528 11880
rect 3660 11840 3666 11852
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 5902 11880 5908 11892
rect 5863 11852 5908 11880
rect 5902 11840 5908 11852
rect 5960 11840 5966 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 7466 11880 7472 11892
rect 7248 11852 7472 11880
rect 7248 11840 7254 11852
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 8389 11883 8447 11889
rect 8389 11849 8401 11883
rect 8435 11880 8447 11883
rect 9214 11880 9220 11892
rect 8435 11852 9220 11880
rect 8435 11849 8447 11852
rect 8389 11843 8447 11849
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 12250 11880 12256 11892
rect 9916 11852 12256 11880
rect 9916 11840 9922 11852
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 1946 11772 1952 11824
rect 2004 11812 2010 11824
rect 2004 11784 3464 11812
rect 2004 11772 2010 11784
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11676 2007 11679
rect 2774 11676 2780 11688
rect 1995 11648 2780 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 3436 11676 3464 11784
rect 3510 11772 3516 11824
rect 3568 11812 3574 11824
rect 4246 11812 4252 11824
rect 3568 11784 4252 11812
rect 3568 11772 3574 11784
rect 4246 11772 4252 11784
rect 4304 11772 4310 11824
rect 6178 11772 6184 11824
rect 6236 11812 6242 11824
rect 9674 11812 9680 11824
rect 6236 11784 9680 11812
rect 6236 11772 6242 11784
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 9766 11772 9772 11824
rect 9824 11812 9830 11824
rect 10042 11812 10048 11824
rect 9824 11784 10048 11812
rect 9824 11772 9830 11784
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 10781 11815 10839 11821
rect 10781 11781 10793 11815
rect 10827 11812 10839 11815
rect 12802 11812 12808 11824
rect 10827 11784 12808 11812
rect 10827 11781 10839 11784
rect 10781 11775 10839 11781
rect 12802 11772 12808 11784
rect 12860 11772 12866 11824
rect 3602 11744 3608 11756
rect 3563 11716 3608 11744
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 5074 11704 5080 11756
rect 5132 11744 5138 11756
rect 6546 11744 6552 11756
rect 5132 11716 6552 11744
rect 5132 11704 5138 11716
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 7469 11747 7527 11753
rect 6696 11716 7328 11744
rect 6696 11704 6702 11716
rect 4617 11679 4675 11685
rect 4617 11676 4629 11679
rect 3436 11648 4629 11676
rect 4617 11645 4629 11648
rect 4663 11645 4675 11679
rect 4617 11639 4675 11645
rect 3421 11611 3479 11617
rect 3421 11577 3433 11611
rect 3467 11608 3479 11611
rect 4062 11608 4068 11620
rect 3467 11580 4068 11608
rect 3467 11577 3479 11580
rect 3421 11571 3479 11577
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 4632 11608 4660 11639
rect 5902 11636 5908 11688
rect 5960 11676 5966 11688
rect 7006 11676 7012 11688
rect 5960 11648 7012 11676
rect 5960 11636 5966 11648
rect 7006 11636 7012 11648
rect 7064 11676 7070 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 7064 11648 7205 11676
rect 7064 11636 7070 11648
rect 7193 11645 7205 11648
rect 7239 11645 7251 11679
rect 7300 11676 7328 11716
rect 7469 11713 7481 11747
rect 7515 11744 7527 11747
rect 7558 11744 7564 11756
rect 7515 11716 7564 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 9030 11744 9036 11756
rect 8991 11716 9036 11744
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 11054 11744 11060 11756
rect 9364 11716 11060 11744
rect 9364 11704 9370 11716
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 11425 11747 11483 11753
rect 11425 11713 11437 11747
rect 11471 11744 11483 11747
rect 11514 11744 11520 11756
rect 11471 11716 11520 11744
rect 11471 11713 11483 11716
rect 11425 11707 11483 11713
rect 11514 11704 11520 11716
rect 11572 11744 11578 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 11572 11716 13001 11744
rect 11572 11704 11578 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 8846 11676 8852 11688
rect 7300 11648 8524 11676
rect 8807 11648 8852 11676
rect 7193 11639 7251 11645
rect 8386 11608 8392 11620
rect 4632 11580 8392 11608
rect 8386 11568 8392 11580
rect 8444 11568 8450 11620
rect 8496 11608 8524 11648
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 9214 11636 9220 11688
rect 9272 11676 9278 11688
rect 11146 11676 11152 11688
rect 9272 11648 11008 11676
rect 11107 11648 11152 11676
rect 9272 11636 9278 11648
rect 10870 11608 10876 11620
rect 8496 11580 10876 11608
rect 10870 11568 10876 11580
rect 10928 11568 10934 11620
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 2133 11543 2191 11549
rect 2133 11540 2145 11543
rect 1636 11512 2145 11540
rect 1636 11500 1642 11512
rect 2133 11509 2145 11512
rect 2179 11509 2191 11543
rect 3050 11540 3056 11552
rect 3011 11512 3056 11540
rect 2133 11503 2191 11509
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 3513 11543 3571 11549
rect 3513 11509 3525 11543
rect 3559 11540 3571 11543
rect 3786 11540 3792 11552
rect 3559 11512 3792 11540
rect 3559 11509 3571 11512
rect 3513 11503 3571 11509
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4801 11543 4859 11549
rect 4801 11540 4813 11543
rect 4396 11512 4813 11540
rect 4396 11500 4402 11512
rect 4801 11509 4813 11512
rect 4847 11509 4859 11543
rect 4801 11503 4859 11509
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6696 11512 6837 11540
rect 6696 11500 6702 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 7285 11543 7343 11549
rect 7285 11509 7297 11543
rect 7331 11540 7343 11543
rect 7466 11540 7472 11552
rect 7331 11512 7472 11540
rect 7331 11509 7343 11512
rect 7285 11503 7343 11509
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 8757 11543 8815 11549
rect 8757 11509 8769 11543
rect 8803 11540 8815 11543
rect 8938 11540 8944 11552
rect 8803 11512 8944 11540
rect 8803 11509 8815 11512
rect 8757 11503 8815 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 10778 11540 10784 11552
rect 9456 11512 10784 11540
rect 9456 11500 9462 11512
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 10980 11540 11008 11648
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 12894 11676 12900 11688
rect 12855 11648 12900 11676
rect 12894 11636 12900 11648
rect 12952 11636 12958 11688
rect 12805 11611 12863 11617
rect 12805 11608 12817 11611
rect 11164 11580 12817 11608
rect 11164 11540 11192 11580
rect 12805 11577 12817 11580
rect 12851 11577 12863 11611
rect 12805 11571 12863 11577
rect 13538 11568 13544 11620
rect 13596 11608 13602 11620
rect 15562 11608 15568 11620
rect 13596 11580 15568 11608
rect 13596 11568 13602 11580
rect 15562 11568 15568 11580
rect 15620 11568 15626 11620
rect 10980 11512 11192 11540
rect 11241 11543 11299 11549
rect 11241 11509 11253 11543
rect 11287 11540 11299 11543
rect 11606 11540 11612 11552
rect 11287 11512 11612 11540
rect 11287 11509 11299 11512
rect 11241 11503 11299 11509
rect 11606 11500 11612 11512
rect 11664 11500 11670 11552
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 12894 11540 12900 11552
rect 12483 11512 12900 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 1104 11450 14812 11472
rect 1104 11398 5579 11450
rect 5631 11398 5643 11450
rect 5695 11398 5707 11450
rect 5759 11398 5771 11450
rect 5823 11398 10176 11450
rect 10228 11398 10240 11450
rect 10292 11398 10304 11450
rect 10356 11398 10368 11450
rect 10420 11398 14812 11450
rect 1104 11376 14812 11398
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 4433 11339 4491 11345
rect 4433 11336 4445 11339
rect 2179 11308 4445 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 4433 11305 4445 11308
rect 4479 11305 4491 11339
rect 4433 11299 4491 11305
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 8389 11339 8447 11345
rect 8389 11336 8401 11339
rect 6512 11308 8401 11336
rect 6512 11296 6518 11308
rect 8389 11305 8401 11308
rect 8435 11336 8447 11339
rect 8435 11308 13400 11336
rect 8435 11305 8447 11308
rect 8389 11299 8447 11305
rect 3050 11228 3056 11280
rect 3108 11268 3114 11280
rect 4525 11271 4583 11277
rect 4525 11268 4537 11271
rect 3108 11240 4537 11268
rect 3108 11228 3114 11240
rect 4525 11237 4537 11240
rect 4571 11237 4583 11271
rect 10134 11268 10140 11280
rect 4525 11231 4583 11237
rect 5644 11240 10140 11268
rect 2130 11160 2136 11212
rect 2188 11200 2194 11212
rect 5644 11209 5672 11240
rect 10134 11228 10140 11240
rect 10192 11268 10198 11280
rect 10192 11240 10456 11268
rect 10192 11228 10198 11240
rect 2501 11203 2559 11209
rect 2501 11200 2513 11203
rect 2188 11172 2513 11200
rect 2188 11160 2194 11172
rect 2501 11169 2513 11172
rect 2547 11169 2559 11203
rect 2501 11163 2559 11169
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11169 5687 11203
rect 5629 11163 5687 11169
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 9214 11200 9220 11212
rect 6880 11172 9220 11200
rect 6880 11160 6886 11172
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 9933 11203 9991 11209
rect 9933 11200 9945 11203
rect 9824 11172 9945 11200
rect 9824 11160 9830 11172
rect 9933 11169 9945 11172
rect 9979 11169 9991 11203
rect 10428 11200 10456 11240
rect 11054 11200 11060 11212
rect 10428 11172 11060 11200
rect 9933 11163 9991 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 13372 11209 13400 11308
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11169 13415 11203
rect 13357 11163 13415 11169
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2593 11135 2651 11141
rect 2593 11132 2605 11135
rect 2280 11104 2605 11132
rect 2280 11092 2286 11104
rect 2593 11101 2605 11104
rect 2639 11101 2651 11135
rect 2593 11095 2651 11101
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 3142 11132 3148 11144
rect 2731 11104 3148 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 3142 11092 3148 11104
rect 3200 11132 3206 11144
rect 3602 11132 3608 11144
rect 3200 11104 3608 11132
rect 3200 11092 3206 11104
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7650 11132 7656 11144
rect 7055 11104 7656 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 1394 11024 1400 11076
rect 1452 11064 1458 11076
rect 2406 11064 2412 11076
rect 1452 11036 2412 11064
rect 1452 11024 1458 11036
rect 2406 11024 2412 11036
rect 2464 11024 2470 11076
rect 3878 11024 3884 11076
rect 3936 11064 3942 11076
rect 4065 11067 4123 11073
rect 4065 11064 4077 11067
rect 3936 11036 4077 11064
rect 3936 11024 3942 11036
rect 4065 11033 4077 11036
rect 4111 11033 4123 11067
rect 4065 11027 4123 11033
rect 4246 11024 4252 11076
rect 4304 11064 4310 11076
rect 4724 11064 4752 11095
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 8478 11132 8484 11144
rect 7944 11104 8484 11132
rect 4304 11036 4752 11064
rect 5813 11067 5871 11073
rect 4304 11024 4310 11036
rect 5813 11033 5825 11067
rect 5859 11064 5871 11067
rect 6362 11064 6368 11076
rect 5859 11036 6368 11064
rect 5859 11033 5871 11036
rect 5813 11027 5871 11033
rect 6362 11024 6368 11036
rect 6420 11024 6426 11076
rect 6730 11024 6736 11076
rect 6788 11064 6794 11076
rect 7944 11064 7972 11104
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 9677 11135 9735 11141
rect 8628 11104 8673 11132
rect 8628 11092 8634 11104
rect 9677 11101 9689 11135
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 6788 11036 7972 11064
rect 8021 11067 8079 11073
rect 6788 11024 6794 11036
rect 8021 11033 8033 11067
rect 8067 11064 8079 11067
rect 8938 11064 8944 11076
rect 8067 11036 8944 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 9306 10996 9312 11008
rect 4028 10968 9312 10996
rect 4028 10956 4034 10968
rect 9306 10956 9312 10968
rect 9364 10956 9370 11008
rect 9692 10996 9720 11095
rect 10686 11092 10692 11144
rect 10744 11132 10750 11144
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 10744 11104 11897 11132
rect 10744 11092 10750 11104
rect 11885 11101 11897 11104
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 11057 11067 11115 11073
rect 11057 11033 11069 11067
rect 11103 11064 11115 11067
rect 12066 11064 12072 11076
rect 11103 11036 12072 11064
rect 11103 11033 11115 11036
rect 11057 11027 11115 11033
rect 12066 11024 12072 11036
rect 12124 11024 12130 11076
rect 12342 11024 12348 11076
rect 12400 11064 12406 11076
rect 13541 11067 13599 11073
rect 13541 11064 13553 11067
rect 12400 11036 13553 11064
rect 12400 11024 12406 11036
rect 13541 11033 13553 11036
rect 13587 11033 13599 11067
rect 13541 11027 13599 11033
rect 10962 10996 10968 11008
rect 9692 10968 10968 10996
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 1104 10906 14812 10928
rect 1104 10854 3280 10906
rect 3332 10854 3344 10906
rect 3396 10854 3408 10906
rect 3460 10854 3472 10906
rect 3524 10854 7878 10906
rect 7930 10854 7942 10906
rect 7994 10854 8006 10906
rect 8058 10854 8070 10906
rect 8122 10854 12475 10906
rect 12527 10854 12539 10906
rect 12591 10854 12603 10906
rect 12655 10854 12667 10906
rect 12719 10854 14812 10906
rect 1104 10832 14812 10854
rect 8481 10795 8539 10801
rect 8481 10761 8493 10795
rect 8527 10792 8539 10795
rect 9122 10792 9128 10804
rect 8527 10764 9128 10792
rect 8527 10761 8539 10764
rect 8481 10755 8539 10761
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 12805 10795 12863 10801
rect 12805 10792 12817 10795
rect 9232 10764 12817 10792
rect 5810 10724 5816 10736
rect 3988 10696 5816 10724
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 1780 10520 1808 10551
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 3142 10597 3148 10600
rect 2869 10591 2927 10597
rect 2869 10588 2881 10591
rect 2556 10560 2881 10588
rect 2556 10548 2562 10560
rect 2869 10557 2881 10560
rect 2915 10557 2927 10591
rect 3136 10588 3148 10597
rect 3103 10560 3148 10588
rect 2869 10551 2927 10557
rect 3136 10551 3148 10560
rect 3142 10548 3148 10551
rect 3200 10548 3206 10600
rect 2958 10520 2964 10532
rect 1780 10492 2964 10520
rect 2958 10480 2964 10492
rect 3016 10520 3022 10532
rect 3988 10520 4016 10696
rect 5810 10684 5816 10696
rect 5868 10684 5874 10736
rect 5994 10684 6000 10736
rect 6052 10724 6058 10736
rect 9232 10724 9260 10764
rect 12805 10761 12817 10764
rect 12851 10761 12863 10795
rect 12805 10755 12863 10761
rect 6052 10696 9260 10724
rect 6052 10684 6058 10696
rect 9490 10684 9496 10736
rect 9548 10724 9554 10736
rect 11425 10727 11483 10733
rect 9548 10696 11376 10724
rect 9548 10684 9554 10696
rect 6178 10616 6184 10668
rect 6236 10656 6242 10668
rect 7469 10659 7527 10665
rect 7469 10656 7481 10659
rect 6236 10628 7481 10656
rect 6236 10616 6242 10628
rect 7469 10625 7481 10628
rect 7515 10656 7527 10659
rect 7558 10656 7564 10668
rect 7515 10628 7564 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 8018 10616 8024 10668
rect 8076 10656 8082 10668
rect 8570 10656 8576 10668
rect 8076 10628 8576 10656
rect 8076 10616 8082 10628
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8938 10656 8944 10668
rect 8899 10628 8944 10656
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 11054 10656 11060 10668
rect 9088 10628 9133 10656
rect 9232 10628 11060 10656
rect 9088 10616 9094 10628
rect 5077 10591 5135 10597
rect 5077 10557 5089 10591
rect 5123 10588 5135 10591
rect 5123 10560 7503 10588
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 3016 10492 4016 10520
rect 3016 10480 3022 10492
rect 6086 10480 6092 10532
rect 6144 10520 6150 10532
rect 7377 10523 7435 10529
rect 7377 10520 7389 10523
rect 6144 10492 7389 10520
rect 6144 10480 6150 10492
rect 7377 10489 7389 10492
rect 7423 10489 7435 10523
rect 7475 10520 7503 10560
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 9232 10588 9260 10628
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11348 10656 11376 10696
rect 11425 10693 11437 10727
rect 11471 10724 11483 10727
rect 13538 10724 13544 10736
rect 11471 10696 13544 10724
rect 11471 10693 11483 10696
rect 11425 10687 11483 10693
rect 13538 10684 13544 10696
rect 13596 10684 13602 10736
rect 11698 10656 11704 10668
rect 11348 10628 11704 10656
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 13357 10659 13415 10665
rect 13357 10656 13369 10659
rect 12124 10628 13369 10656
rect 12124 10616 12130 10628
rect 13357 10625 13369 10628
rect 13403 10625 13415 10659
rect 13357 10619 13415 10625
rect 8444 10560 9260 10588
rect 8444 10548 8450 10560
rect 9306 10548 9312 10600
rect 9364 10588 9370 10600
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9364 10560 10057 10588
rect 9364 10548 9370 10560
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11241 10591 11299 10597
rect 11241 10588 11253 10591
rect 11204 10560 11253 10588
rect 11204 10548 11210 10560
rect 11241 10557 11253 10560
rect 11287 10557 11299 10591
rect 11241 10551 11299 10557
rect 7475 10492 11284 10520
rect 7377 10483 7435 10489
rect 1949 10455 2007 10461
rect 1949 10421 1961 10455
rect 1995 10452 2007 10455
rect 2314 10452 2320 10464
rect 1995 10424 2320 10452
rect 1995 10421 2007 10424
rect 1949 10415 2007 10421
rect 2314 10412 2320 10424
rect 2372 10412 2378 10464
rect 4246 10452 4252 10464
rect 4207 10424 4252 10452
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 5258 10452 5264 10464
rect 5219 10424 5264 10452
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 6917 10455 6975 10461
rect 6917 10421 6929 10455
rect 6963 10452 6975 10455
rect 7098 10452 7104 10464
rect 6963 10424 7104 10452
rect 6963 10421 6975 10424
rect 6917 10415 6975 10421
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7285 10455 7343 10461
rect 7285 10421 7297 10455
rect 7331 10452 7343 10455
rect 7558 10452 7564 10464
rect 7331 10424 7564 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 8754 10412 8760 10464
rect 8812 10452 8818 10464
rect 8849 10455 8907 10461
rect 8849 10452 8861 10455
rect 8812 10424 8861 10452
rect 8812 10412 8818 10424
rect 8849 10421 8861 10424
rect 8895 10421 8907 10455
rect 8849 10415 8907 10421
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 9732 10424 10241 10452
rect 9732 10412 9738 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 11256 10452 11284 10492
rect 11698 10480 11704 10532
rect 11756 10520 11762 10532
rect 13265 10523 13323 10529
rect 13265 10520 13277 10523
rect 11756 10492 13277 10520
rect 11756 10480 11762 10492
rect 13265 10489 13277 10492
rect 13311 10489 13323 10523
rect 13265 10483 13323 10489
rect 11606 10452 11612 10464
rect 11256 10424 11612 10452
rect 10229 10415 10287 10421
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 13170 10452 13176 10464
rect 13131 10424 13176 10452
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 1104 10362 14812 10384
rect 1104 10310 5579 10362
rect 5631 10310 5643 10362
rect 5695 10310 5707 10362
rect 5759 10310 5771 10362
rect 5823 10310 10176 10362
rect 10228 10310 10240 10362
rect 10292 10310 10304 10362
rect 10356 10310 10368 10362
rect 10420 10310 14812 10362
rect 1104 10288 14812 10310
rect 2498 10208 2504 10260
rect 2556 10208 2562 10260
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 4172 10220 6224 10248
rect 2516 10180 2544 10208
rect 1780 10152 2636 10180
rect 1780 10121 1808 10152
rect 1765 10115 1823 10121
rect 1765 10081 1777 10115
rect 1811 10081 1823 10115
rect 1765 10075 1823 10081
rect 2032 10115 2090 10121
rect 2032 10081 2044 10115
rect 2078 10112 2090 10115
rect 2498 10112 2504 10124
rect 2078 10084 2504 10112
rect 2078 10081 2090 10084
rect 2032 10075 2090 10081
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 2608 10112 2636 10152
rect 2682 10140 2688 10192
rect 2740 10180 2746 10192
rect 4172 10180 4200 10220
rect 2740 10152 4200 10180
rect 2740 10140 2746 10152
rect 4246 10140 4252 10192
rect 4304 10180 4310 10192
rect 4954 10183 5012 10189
rect 4954 10180 4966 10183
rect 4304 10152 4966 10180
rect 4304 10140 4310 10152
rect 4954 10149 4966 10152
rect 5000 10149 5012 10183
rect 4954 10143 5012 10149
rect 2608 10084 4660 10112
rect 4632 10056 4660 10084
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 4709 10047 4767 10053
rect 4709 10044 4721 10047
rect 4672 10016 4721 10044
rect 4672 10004 4678 10016
rect 4709 10013 4721 10016
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 3970 9936 3976 9988
rect 4028 9976 4034 9988
rect 4246 9976 4252 9988
rect 4028 9948 4252 9976
rect 4028 9936 4034 9948
rect 4246 9936 4252 9948
rect 4304 9936 4310 9988
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 6089 9979 6147 9985
rect 6089 9976 6101 9979
rect 5868 9948 6101 9976
rect 5868 9936 5874 9948
rect 6089 9945 6101 9948
rect 6135 9945 6147 9979
rect 6089 9939 6147 9945
rect 2406 9868 2412 9920
rect 2464 9908 2470 9920
rect 5994 9908 6000 9920
rect 2464 9880 6000 9908
rect 2464 9868 2470 9880
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 6196 9908 6224 10220
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7466 10248 7472 10260
rect 7248 10220 7472 10248
rect 7248 10208 7254 10220
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 8570 10248 8576 10260
rect 8483 10220 8576 10248
rect 8570 10208 8576 10220
rect 8628 10248 8634 10260
rect 9030 10248 9036 10260
rect 8628 10220 9036 10248
rect 8628 10208 8634 10220
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9122 10208 9128 10260
rect 9180 10248 9186 10260
rect 12250 10248 12256 10260
rect 9180 10220 12256 10248
rect 9180 10208 9186 10220
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 7006 10140 7012 10192
rect 7064 10180 7070 10192
rect 10042 10180 10048 10192
rect 7064 10152 9812 10180
rect 7064 10140 7070 10152
rect 7466 10121 7472 10124
rect 7460 10112 7472 10121
rect 7427 10084 7472 10112
rect 7460 10075 7472 10084
rect 7524 10112 7530 10124
rect 8018 10112 8024 10124
rect 7524 10084 8024 10112
rect 7466 10072 7472 10075
rect 7524 10072 7530 10084
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 9306 10112 9312 10124
rect 8260 10084 9312 10112
rect 8260 10072 8266 10084
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 9784 10112 9812 10152
rect 9876 10152 10048 10180
rect 9876 10112 9904 10152
rect 10042 10140 10048 10152
rect 10100 10140 10106 10192
rect 9784 10084 9904 10112
rect 9953 10115 10011 10121
rect 9953 10081 9965 10115
rect 9999 10081 10011 10115
rect 9953 10075 10011 10081
rect 7190 10044 7196 10056
rect 7151 10016 7196 10044
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 9968 9908 9996 10075
rect 10962 10072 10968 10124
rect 11020 10112 11026 10124
rect 11057 10115 11115 10121
rect 11057 10112 11069 10115
rect 11020 10084 11069 10112
rect 11020 10072 11026 10084
rect 11057 10081 11069 10084
rect 11103 10081 11115 10115
rect 11057 10075 11115 10081
rect 11324 10115 11382 10121
rect 11324 10081 11336 10115
rect 11370 10112 11382 10115
rect 11606 10112 11612 10124
rect 11370 10084 11612 10112
rect 11370 10081 11382 10084
rect 11324 10075 11382 10081
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 11698 10072 11704 10124
rect 11756 10112 11762 10124
rect 13357 10115 13415 10121
rect 13357 10112 13369 10115
rect 11756 10084 13369 10112
rect 11756 10072 11762 10084
rect 13357 10081 13369 10084
rect 13403 10081 13415 10115
rect 13357 10075 13415 10081
rect 12158 9936 12164 9988
rect 12216 9976 12222 9988
rect 13541 9979 13599 9985
rect 13541 9976 13553 9979
rect 12216 9948 13553 9976
rect 12216 9936 12222 9948
rect 13541 9945 13553 9948
rect 13587 9945 13599 9979
rect 13541 9939 13599 9945
rect 6196 9880 9996 9908
rect 10137 9911 10195 9917
rect 10137 9877 10149 9911
rect 10183 9908 10195 9911
rect 10594 9908 10600 9920
rect 10183 9880 10600 9908
rect 10183 9877 10195 9880
rect 10137 9871 10195 9877
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 12437 9911 12495 9917
rect 12437 9877 12449 9911
rect 12483 9908 12495 9911
rect 12986 9908 12992 9920
rect 12483 9880 12992 9908
rect 12483 9877 12495 9880
rect 12437 9871 12495 9877
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 1104 9818 14812 9840
rect 1104 9766 3280 9818
rect 3332 9766 3344 9818
rect 3396 9766 3408 9818
rect 3460 9766 3472 9818
rect 3524 9766 7878 9818
rect 7930 9766 7942 9818
rect 7994 9766 8006 9818
rect 8058 9766 8070 9818
rect 8122 9766 12475 9818
rect 12527 9766 12539 9818
rect 12591 9766 12603 9818
rect 12655 9766 12667 9818
rect 12719 9766 14812 9818
rect 1104 9744 14812 9766
rect 1486 9664 1492 9716
rect 1544 9704 1550 9716
rect 2866 9704 2872 9716
rect 1544 9676 2872 9704
rect 1544 9664 1550 9676
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4304 9676 5580 9704
rect 4304 9664 4310 9676
rect 2222 9636 2228 9648
rect 2183 9608 2228 9636
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 5552 9636 5580 9676
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 6178 9704 6184 9716
rect 5868 9676 6184 9704
rect 5868 9664 5874 9676
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 7944 9676 10180 9704
rect 6270 9636 6276 9648
rect 5552 9608 6276 9636
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 7374 9636 7380 9648
rect 7116 9608 7380 9636
rect 2498 9528 2504 9580
rect 2556 9568 2562 9580
rect 2777 9571 2835 9577
rect 2777 9568 2789 9571
rect 2556 9540 2789 9568
rect 2556 9528 2562 9540
rect 2777 9537 2789 9540
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 5074 9528 5080 9580
rect 5132 9568 5138 9580
rect 7116 9568 7144 9608
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 5132 9540 7144 9568
rect 5132 9528 5138 9540
rect 7190 9528 7196 9580
rect 7248 9568 7254 9580
rect 7944 9577 7972 9676
rect 9309 9639 9367 9645
rect 9309 9605 9321 9639
rect 9355 9636 9367 9639
rect 9766 9636 9772 9648
rect 9355 9608 9772 9636
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 7929 9571 7987 9577
rect 7929 9568 7941 9571
rect 7248 9540 7941 9568
rect 7248 9528 7254 9540
rect 7929 9537 7941 9540
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 10042 9528 10048 9580
rect 10100 9568 10106 9580
rect 10152 9577 10180 9676
rect 11146 9664 11152 9716
rect 11204 9704 11210 9716
rect 13078 9704 13084 9716
rect 11204 9676 13084 9704
rect 11204 9664 11210 9676
rect 13078 9664 13084 9676
rect 13136 9704 13142 9716
rect 13354 9704 13360 9716
rect 13136 9676 13360 9704
rect 13136 9664 13142 9676
rect 13354 9664 13360 9676
rect 13412 9664 13418 9716
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 10100 9540 10149 9568
rect 10100 9528 10106 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 12894 9568 12900 9580
rect 12855 9540 12900 9568
rect 10137 9531 10195 9537
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 12986 9528 12992 9580
rect 13044 9568 13050 9580
rect 13044 9540 13089 9568
rect 13044 9528 13050 9540
rect 1026 9460 1032 9512
rect 1084 9500 1090 9512
rect 1670 9500 1676 9512
rect 1084 9472 1676 9500
rect 1084 9460 1090 9472
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 2590 9500 2596 9512
rect 2551 9472 2596 9500
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 2685 9503 2743 9509
rect 2685 9469 2697 9503
rect 2731 9500 2743 9503
rect 3602 9500 3608 9512
rect 2731 9472 3608 9500
rect 2731 9469 2743 9472
rect 2685 9463 2743 9469
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 3970 9500 3976 9512
rect 3927 9472 3976 9500
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 3970 9460 3976 9472
rect 4028 9500 4034 9512
rect 4614 9500 4620 9512
rect 4028 9472 4620 9500
rect 4028 9460 4034 9472
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 5442 9500 5448 9512
rect 5224 9472 5448 9500
rect 5224 9460 5230 9472
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 7006 9500 7012 9512
rect 6871 9472 7012 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 7006 9460 7012 9472
rect 7064 9500 7070 9512
rect 7558 9500 7564 9512
rect 7064 9472 7564 9500
rect 7064 9460 7070 9472
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 8196 9503 8254 9509
rect 8196 9469 8208 9503
rect 8242 9500 8254 9503
rect 8570 9500 8576 9512
rect 8242 9472 8576 9500
rect 8242 9469 8254 9472
rect 8196 9463 8254 9469
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 12802 9500 12808 9512
rect 12763 9472 12808 9500
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 3326 9392 3332 9444
rect 3384 9432 3390 9444
rect 4154 9441 4160 9444
rect 4126 9435 4160 9441
rect 4126 9432 4138 9435
rect 3384 9404 4138 9432
rect 3384 9392 3390 9404
rect 4126 9401 4138 9404
rect 4212 9432 4218 9444
rect 10404 9435 10462 9441
rect 4212 9404 4274 9432
rect 4540 9404 9904 9432
rect 4126 9395 4160 9401
rect 4154 9392 4160 9395
rect 4212 9392 4218 9404
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 4540 9364 4568 9404
rect 1728 9336 4568 9364
rect 1728 9324 1734 9336
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 4672 9336 5273 9364
rect 4672 9324 4678 9336
rect 5261 9333 5273 9336
rect 5307 9333 5319 9367
rect 5261 9327 5319 9333
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9364 7067 9367
rect 7282 9364 7288 9376
rect 7055 9336 7288 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 9876 9364 9904 9404
rect 10404 9401 10416 9435
rect 10450 9432 10462 9435
rect 12066 9432 12072 9444
rect 10450 9404 12072 9432
rect 10450 9401 10462 9404
rect 10404 9395 10462 9401
rect 12066 9392 12072 9404
rect 12124 9392 12130 9444
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 9876 9336 11529 9364
rect 11517 9333 11529 9336
rect 11563 9364 11575 9367
rect 11606 9364 11612 9376
rect 11563 9336 11612 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12710 9364 12716 9376
rect 12483 9336 12716 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 1104 9274 14812 9296
rect 1104 9222 5579 9274
rect 5631 9222 5643 9274
rect 5695 9222 5707 9274
rect 5759 9222 5771 9274
rect 5823 9222 10176 9274
rect 10228 9222 10240 9274
rect 10292 9222 10304 9274
rect 10356 9222 10368 9274
rect 10420 9222 14812 9274
rect 1104 9200 14812 9222
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 2869 9163 2927 9169
rect 2869 9160 2881 9163
rect 2740 9132 2881 9160
rect 2740 9120 2746 9132
rect 2869 9129 2881 9132
rect 2915 9129 2927 9163
rect 4062 9160 4068 9172
rect 4023 9132 4068 9160
rect 2869 9123 2927 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 4571 9132 5641 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 5629 9123 5687 9129
rect 5997 9163 6055 9169
rect 5997 9129 6009 9163
rect 6043 9160 6055 9163
rect 7006 9160 7012 9172
rect 6043 9132 7012 9160
rect 6043 9129 6055 9132
rect 5997 9123 6055 9129
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 7742 9160 7748 9172
rect 7699 9132 7748 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 11054 9160 11060 9172
rect 8628 9132 11060 9160
rect 8628 9120 8634 9132
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 12710 9160 12716 9172
rect 12671 9132 12716 9160
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 13814 9160 13820 9172
rect 13320 9132 13820 9160
rect 13320 9120 13326 9132
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 5442 9092 5448 9104
rect 4212 9064 5448 9092
rect 4212 9052 4218 9064
rect 5442 9052 5448 9064
rect 5500 9092 5506 9104
rect 5810 9092 5816 9104
rect 5500 9064 5816 9092
rect 5500 9052 5506 9064
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 10404 9095 10462 9101
rect 6012 9064 10272 9092
rect 2774 9024 2780 9036
rect 2735 8996 2780 9024
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 4430 9024 4436 9036
rect 4343 8996 4436 9024
rect 4430 8984 4436 8996
rect 4488 9024 4494 9036
rect 6012 9024 6040 9064
rect 4488 8996 6040 9024
rect 6089 9027 6147 9033
rect 4488 8984 4494 8996
rect 6089 8993 6101 9027
rect 6135 9024 6147 9027
rect 6270 9024 6276 9036
rect 6135 8996 6276 9024
rect 6135 8993 6147 8996
rect 6089 8987 6147 8993
rect 6270 8984 6276 8996
rect 6328 9024 6334 9036
rect 6328 8996 6960 9024
rect 6328 8984 6334 8996
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 2498 8956 2504 8968
rect 1443 8928 2504 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3326 8956 3332 8968
rect 3099 8928 3332 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 4614 8956 4620 8968
rect 4575 8928 4620 8956
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 5810 8916 5816 8968
rect 5868 8956 5874 8968
rect 6181 8959 6239 8965
rect 6181 8956 6193 8959
rect 5868 8928 6193 8956
rect 5868 8916 5874 8928
rect 6181 8925 6193 8928
rect 6227 8925 6239 8959
rect 6932 8956 6960 8996
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 7064 8996 7573 9024
rect 7064 8984 7070 8996
rect 7561 8993 7573 8996
rect 7607 8993 7619 9027
rect 7561 8987 7619 8993
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 8941 9027 8999 9033
rect 8941 9024 8953 9027
rect 8260 8996 8953 9024
rect 8260 8984 8266 8996
rect 8941 8993 8953 8996
rect 8987 8993 8999 9027
rect 8941 8987 8999 8993
rect 10042 8984 10048 9036
rect 10100 9024 10106 9036
rect 10137 9027 10195 9033
rect 10137 9024 10149 9027
rect 10100 8996 10149 9024
rect 10100 8984 10106 8996
rect 10137 8993 10149 8996
rect 10183 8993 10195 9027
rect 10244 9024 10272 9064
rect 10404 9061 10416 9095
rect 10450 9092 10462 9095
rect 12986 9092 12992 9104
rect 10450 9064 12992 9092
rect 10450 9061 10462 9064
rect 10404 9055 10462 9061
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 13262 9024 13268 9036
rect 10244 8996 13268 9024
rect 10137 8987 10195 8993
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 6932 8928 7420 8956
rect 6181 8919 6239 8925
rect 842 8848 848 8900
rect 900 8888 906 8900
rect 5902 8888 5908 8900
rect 900 8860 5908 8888
rect 900 8848 906 8860
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 7392 8888 7420 8928
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7708 8928 7757 8956
rect 7708 8916 7714 8928
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 12802 8956 12808 8968
rect 12763 8928 12808 8956
rect 7745 8919 7803 8925
rect 12802 8916 12808 8928
rect 12860 8916 12866 8968
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8925 12955 8959
rect 12897 8919 12955 8925
rect 8294 8888 8300 8900
rect 7392 8860 8300 8888
rect 8294 8848 8300 8860
rect 8352 8848 8358 8900
rect 9214 8848 9220 8900
rect 9272 8888 9278 8900
rect 11514 8888 11520 8900
rect 9272 8860 9904 8888
rect 11427 8860 11520 8888
rect 9272 8848 9278 8860
rect 2409 8823 2467 8829
rect 2409 8789 2421 8823
rect 2455 8820 2467 8823
rect 4062 8820 4068 8832
rect 2455 8792 4068 8820
rect 2455 8789 2467 8792
rect 2409 8783 2467 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 7193 8823 7251 8829
rect 7193 8789 7205 8823
rect 7239 8820 7251 8823
rect 8478 8820 8484 8832
rect 7239 8792 8484 8820
rect 7239 8789 7251 8792
rect 7193 8783 7251 8789
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 8757 8823 8815 8829
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 9766 8820 9772 8832
rect 8803 8792 9772 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 9876 8820 9904 8860
rect 11514 8848 11520 8860
rect 11572 8888 11578 8900
rect 12912 8888 12940 8919
rect 11572 8860 12940 8888
rect 11572 8848 11578 8860
rect 10778 8820 10784 8832
rect 9876 8792 10784 8820
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 11698 8780 11704 8832
rect 11756 8820 11762 8832
rect 12345 8823 12403 8829
rect 12345 8820 12357 8823
rect 11756 8792 12357 8820
rect 11756 8780 11762 8792
rect 12345 8789 12357 8792
rect 12391 8789 12403 8823
rect 12345 8783 12403 8789
rect 1104 8730 14812 8752
rect 1104 8678 3280 8730
rect 3332 8678 3344 8730
rect 3396 8678 3408 8730
rect 3460 8678 3472 8730
rect 3524 8678 7878 8730
rect 7930 8678 7942 8730
rect 7994 8678 8006 8730
rect 8058 8678 8070 8730
rect 8122 8678 12475 8730
rect 12527 8678 12539 8730
rect 12591 8678 12603 8730
rect 12655 8678 12667 8730
rect 12719 8678 14812 8730
rect 1104 8656 14812 8678
rect 2130 8616 2136 8628
rect 2091 8588 2136 8616
rect 2130 8576 2136 8588
rect 2188 8576 2194 8628
rect 3786 8616 3792 8628
rect 2240 8588 2719 8616
rect 3747 8588 3792 8616
rect 1394 8508 1400 8560
rect 1452 8548 1458 8560
rect 2240 8548 2268 8588
rect 1452 8520 2268 8548
rect 1452 8508 1458 8520
rect 2590 8508 2596 8560
rect 2648 8508 2654 8560
rect 2691 8548 2719 8588
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 10410 8616 10416 8628
rect 3896 8588 10416 8616
rect 3896 8548 3924 8588
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10778 8616 10784 8628
rect 10739 8588 10784 8616
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 12437 8619 12495 8625
rect 12437 8585 12449 8619
rect 12483 8616 12495 8619
rect 12802 8616 12808 8628
rect 12483 8588 12808 8616
rect 12483 8585 12495 8588
rect 12437 8579 12495 8585
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 2691 8520 3924 8548
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 5353 8551 5411 8557
rect 5353 8548 5365 8551
rect 4028 8520 5365 8548
rect 4028 8508 4034 8520
rect 5353 8517 5365 8520
rect 5399 8517 5411 8551
rect 5353 8511 5411 8517
rect 5813 8551 5871 8557
rect 5813 8517 5825 8551
rect 5859 8548 5871 8551
rect 6825 8551 6883 8557
rect 5859 8520 6776 8548
rect 5859 8517 5871 8520
rect 5813 8511 5871 8517
rect 2608 8480 2636 8508
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2608 8452 2697 8480
rect 2685 8449 2697 8452
rect 2731 8480 2743 8483
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 2731 8452 4353 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 4341 8449 4353 8452
rect 4387 8480 4399 8483
rect 4614 8480 4620 8492
rect 4387 8452 4620 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 5902 8480 5908 8492
rect 5552 8452 5908 8480
rect 2498 8412 2504 8424
rect 2459 8384 2504 8412
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 4890 8412 4896 8424
rect 2639 8384 4896 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 5552 8421 5580 8452
rect 5902 8440 5908 8452
rect 5960 8440 5966 8492
rect 6748 8480 6776 8520
rect 6825 8517 6837 8551
rect 6871 8548 6883 8551
rect 9030 8548 9036 8560
rect 6871 8520 9036 8548
rect 6871 8517 6883 8520
rect 6825 8511 6883 8517
rect 9030 8508 9036 8520
rect 9088 8508 9094 8560
rect 10612 8520 12940 8548
rect 7469 8483 7527 8489
rect 6748 8452 7420 8480
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8412 5687 8415
rect 6822 8412 6828 8424
rect 5675 8384 6828 8412
rect 5675 8381 5687 8384
rect 5629 8375 5687 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7193 8415 7251 8421
rect 7193 8412 7205 8415
rect 6972 8384 7205 8412
rect 6972 8372 6978 8384
rect 7193 8381 7205 8384
rect 7239 8381 7251 8415
rect 7392 8412 7420 8452
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7650 8480 7656 8492
rect 7515 8452 7656 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 8938 8480 8944 8492
rect 8899 8452 8944 8480
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 10612 8480 10640 8520
rect 11330 8480 11336 8492
rect 9180 8452 10640 8480
rect 11291 8452 11336 8480
rect 9180 8440 9186 8452
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 12912 8489 12940 8520
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13044 8452 13089 8480
rect 13044 8440 13050 8452
rect 7392 8384 9720 8412
rect 7193 8375 7251 8381
rect 2222 8304 2228 8356
rect 2280 8344 2286 8356
rect 2280 8316 8432 8344
rect 2280 8304 2286 8316
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4157 8279 4215 8285
rect 4157 8276 4169 8279
rect 4120 8248 4169 8276
rect 4120 8236 4126 8248
rect 4157 8245 4169 8248
rect 4203 8245 4215 8279
rect 4157 8239 4215 8245
rect 4249 8279 4307 8285
rect 4249 8245 4261 8279
rect 4295 8276 4307 8279
rect 4614 8276 4620 8288
rect 4295 8248 4620 8276
rect 4295 8245 4307 8248
rect 4249 8239 4307 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 7285 8279 7343 8285
rect 7285 8245 7297 8279
rect 7331 8276 7343 8279
rect 7374 8276 7380 8288
rect 7331 8248 7380 8276
rect 7331 8245 7343 8248
rect 7285 8239 7343 8245
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 8404 8285 8432 8316
rect 8478 8304 8484 8356
rect 8536 8344 8542 8356
rect 8757 8347 8815 8353
rect 8757 8344 8769 8347
rect 8536 8316 8769 8344
rect 8536 8304 8542 8316
rect 8757 8313 8769 8316
rect 8803 8313 8815 8347
rect 8757 8307 8815 8313
rect 8849 8347 8907 8353
rect 8849 8313 8861 8347
rect 8895 8344 8907 8347
rect 9030 8344 9036 8356
rect 8895 8316 9036 8344
rect 8895 8313 8907 8316
rect 8849 8307 8907 8313
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 9692 8344 9720 8384
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 10137 8415 10195 8421
rect 10137 8412 10149 8415
rect 9824 8384 10149 8412
rect 9824 8372 9830 8384
rect 10137 8381 10149 8384
rect 10183 8381 10195 8415
rect 10137 8375 10195 8381
rect 10410 8372 10416 8424
rect 10468 8412 10474 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 10468 8384 12817 8412
rect 10468 8372 10474 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 11146 8344 11152 8356
rect 9692 8316 11008 8344
rect 11107 8316 11152 8344
rect 8389 8279 8447 8285
rect 8389 8245 8401 8279
rect 8435 8245 8447 8279
rect 8389 8239 8447 8245
rect 9953 8279 10011 8285
rect 9953 8245 9965 8279
rect 9999 8276 10011 8279
rect 10042 8276 10048 8288
rect 9999 8248 10048 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 10980 8276 11008 8316
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 11241 8347 11299 8353
rect 11241 8313 11253 8347
rect 11287 8344 11299 8347
rect 12710 8344 12716 8356
rect 11287 8316 12716 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 11054 8276 11060 8288
rect 10980 8248 11060 8276
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 1104 8186 14812 8208
rect 1104 8134 5579 8186
rect 5631 8134 5643 8186
rect 5695 8134 5707 8186
rect 5759 8134 5771 8186
rect 5823 8134 10176 8186
rect 10228 8134 10240 8186
rect 10292 8134 10304 8186
rect 10356 8134 10368 8186
rect 10420 8134 14812 8186
rect 1104 8112 14812 8134
rect 5442 8072 5448 8084
rect 5403 8044 5448 8072
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6822 8072 6828 8084
rect 6604 8044 6828 8072
rect 6604 8032 6610 8044
rect 6822 8032 6828 8044
rect 6880 8072 6886 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 6880 8044 7297 8072
rect 6880 8032 6886 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10100 8044 11100 8072
rect 10100 8032 10106 8044
rect 2777 8007 2835 8013
rect 2777 7973 2789 8007
rect 2823 8004 2835 8007
rect 2866 8004 2872 8016
rect 2823 7976 2872 8004
rect 2823 7973 2835 7976
rect 2777 7967 2835 7973
rect 2866 7964 2872 7976
rect 2924 7964 2930 8016
rect 3602 7964 3608 8016
rect 3660 7964 3666 8016
rect 3970 7964 3976 8016
rect 4028 8004 4034 8016
rect 5258 8004 5264 8016
rect 4028 7976 5264 8004
rect 4028 7964 4034 7976
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 6914 7964 6920 8016
rect 6972 8004 6978 8016
rect 6972 7976 8616 8004
rect 6972 7964 6978 7976
rect 3620 7936 3648 7964
rect 2884 7908 3648 7936
rect 2130 7828 2136 7880
rect 2188 7868 2194 7880
rect 2406 7868 2412 7880
rect 2188 7840 2412 7868
rect 2188 7828 2194 7840
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2884 7877 2912 7908
rect 3786 7896 3792 7948
rect 3844 7936 3850 7948
rect 4321 7939 4379 7945
rect 4321 7936 4333 7939
rect 3844 7908 4333 7936
rect 3844 7896 3850 7908
rect 4321 7905 4333 7908
rect 4367 7905 4379 7939
rect 4321 7899 4379 7905
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 8481 7939 8539 7945
rect 8481 7936 8493 7939
rect 4948 7908 8493 7936
rect 4948 7896 4954 7908
rect 8481 7905 8493 7908
rect 8527 7905 8539 7939
rect 8588 7936 8616 7976
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 8588 7908 10057 7936
rect 8481 7899 8539 7905
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 11072 7936 11100 8044
rect 11416 8007 11474 8013
rect 11416 7973 11428 8007
rect 11462 8004 11474 8007
rect 11514 8004 11520 8016
rect 11462 7976 11520 8004
rect 11462 7973 11474 7976
rect 11416 7967 11474 7973
rect 11514 7964 11520 7976
rect 11572 7964 11578 8016
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 11072 7908 11161 7936
rect 10045 7899 10103 7905
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 11790 7896 11796 7948
rect 11848 7936 11854 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 11848 7908 13369 7936
rect 11848 7896 11854 7908
rect 13357 7905 13369 7908
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3602 7868 3608 7880
rect 3099 7840 3608 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 7374 7868 7380 7880
rect 7335 7840 7380 7868
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7868 7619 7871
rect 7650 7868 7656 7880
rect 7607 7840 7656 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 10870 7868 10876 7880
rect 10192 7840 10876 7868
rect 10192 7828 10198 7840
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 8665 7803 8723 7809
rect 8665 7769 8677 7803
rect 8711 7800 8723 7803
rect 10962 7800 10968 7812
rect 8711 7772 10968 7800
rect 8711 7769 8723 7772
rect 8665 7763 8723 7769
rect 10962 7760 10968 7772
rect 11020 7760 11026 7812
rect 2409 7735 2467 7741
rect 2409 7701 2421 7735
rect 2455 7732 2467 7735
rect 4338 7732 4344 7744
rect 2455 7704 4344 7732
rect 2455 7701 2467 7704
rect 2409 7695 2467 7701
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 6914 7732 6920 7744
rect 6875 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 10229 7735 10287 7741
rect 10229 7701 10241 7735
rect 10275 7732 10287 7735
rect 10870 7732 10876 7744
rect 10275 7704 10876 7732
rect 10275 7701 10287 7704
rect 10229 7695 10287 7701
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 12529 7735 12587 7741
rect 12529 7701 12541 7735
rect 12575 7732 12587 7735
rect 12986 7732 12992 7744
rect 12575 7704 12992 7732
rect 12575 7701 12587 7704
rect 12529 7695 12587 7701
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 13538 7732 13544 7744
rect 13499 7704 13544 7732
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 1104 7642 14812 7664
rect 1104 7590 3280 7642
rect 3332 7590 3344 7642
rect 3396 7590 3408 7642
rect 3460 7590 3472 7642
rect 3524 7590 7878 7642
rect 7930 7590 7942 7642
rect 7994 7590 8006 7642
rect 8058 7590 8070 7642
rect 8122 7590 12475 7642
rect 12527 7590 12539 7642
rect 12591 7590 12603 7642
rect 12655 7590 12667 7642
rect 12719 7590 14812 7642
rect 1104 7568 14812 7590
rect 3697 7531 3755 7537
rect 3697 7497 3709 7531
rect 3743 7528 3755 7531
rect 3786 7528 3792 7540
rect 3743 7500 3792 7528
rect 3743 7497 3755 7500
rect 3697 7491 3755 7497
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 4525 7531 4583 7537
rect 4525 7497 4537 7531
rect 4571 7528 4583 7531
rect 4614 7528 4620 7540
rect 4571 7500 4620 7528
rect 4571 7497 4583 7500
rect 4525 7491 4583 7497
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 7374 7488 7380 7540
rect 7432 7528 7438 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7432 7500 7665 7528
rect 7432 7488 7438 7500
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 10594 7488 10600 7540
rect 10652 7528 10658 7540
rect 11514 7528 11520 7540
rect 10652 7500 11520 7528
rect 10652 7488 10658 7500
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 12802 7528 12808 7540
rect 12483 7500 12808 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 4706 7420 4712 7472
rect 4764 7460 4770 7472
rect 5258 7460 5264 7472
rect 4764 7432 5264 7460
rect 4764 7420 4770 7432
rect 5258 7420 5264 7432
rect 5316 7420 5322 7472
rect 7466 7420 7472 7472
rect 7524 7460 7530 7472
rect 11054 7460 11060 7472
rect 7524 7432 11060 7460
rect 7524 7420 7530 7432
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 4890 7392 4896 7404
rect 3344 7364 4896 7392
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7324 2375 7327
rect 2406 7324 2412 7336
rect 2363 7296 2412 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 3344 7324 3372 7364
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7392 5043 7395
rect 5074 7392 5080 7404
rect 5031 7364 5080 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5442 7392 5448 7404
rect 5215 7364 5448 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 8202 7392 8208 7404
rect 8163 7364 8208 7392
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 10778 7352 10784 7404
rect 10836 7392 10842 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 10836 7364 10885 7392
rect 10836 7352 10842 7364
rect 10873 7361 10885 7364
rect 10919 7392 10931 7395
rect 13078 7392 13084 7404
rect 10919 7364 13084 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 2924 7296 3372 7324
rect 2924 7284 2930 7296
rect 3970 7284 3976 7336
rect 4028 7324 4034 7336
rect 5350 7324 5356 7336
rect 4028 7296 5356 7324
rect 4028 7284 4034 7296
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 8021 7327 8079 7333
rect 8021 7324 8033 7327
rect 7616 7296 8033 7324
rect 7616 7284 7622 7296
rect 8021 7293 8033 7296
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 9217 7327 9275 7333
rect 9217 7324 9229 7327
rect 8720 7296 9229 7324
rect 8720 7284 8726 7296
rect 9217 7293 9229 7296
rect 9263 7293 9275 7327
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 9217 7287 9275 7293
rect 9508 7296 10701 7324
rect 2584 7259 2642 7265
rect 2584 7225 2596 7259
rect 2630 7256 2642 7259
rect 2682 7256 2688 7268
rect 2630 7228 2688 7256
rect 2630 7225 2642 7228
rect 2584 7219 2642 7225
rect 2682 7216 2688 7228
rect 2740 7216 2746 7268
rect 3418 7216 3424 7268
rect 3476 7256 3482 7268
rect 5442 7256 5448 7268
rect 3476 7228 5448 7256
rect 3476 7216 3482 7228
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 6270 7216 6276 7268
rect 6328 7256 6334 7268
rect 6454 7256 6460 7268
rect 6328 7228 6460 7256
rect 6328 7216 6334 7228
rect 6454 7216 6460 7228
rect 6512 7216 6518 7268
rect 9508 7256 9536 7296
rect 10689 7293 10701 7296
rect 10735 7324 10747 7327
rect 11790 7324 11796 7336
rect 10735 7296 11796 7324
rect 10735 7293 10747 7296
rect 10689 7287 10747 7293
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 8036 7228 9536 7256
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3050 7188 3056 7200
rect 2832 7160 3056 7188
rect 2832 7148 2838 7160
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4430 7188 4436 7200
rect 4304 7160 4436 7188
rect 4304 7148 4310 7160
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 4890 7188 4896 7200
rect 4851 7160 4896 7188
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 8036 7188 8064 7228
rect 9950 7216 9956 7268
rect 10008 7256 10014 7268
rect 10781 7259 10839 7265
rect 10781 7256 10793 7259
rect 10008 7228 10793 7256
rect 10008 7216 10014 7228
rect 10781 7225 10793 7228
rect 10827 7225 10839 7259
rect 12802 7256 12808 7268
rect 12763 7228 12808 7256
rect 10781 7219 10839 7225
rect 12802 7216 12808 7228
rect 12860 7216 12866 7268
rect 5224 7160 8064 7188
rect 8113 7191 8171 7197
rect 5224 7148 5230 7160
rect 8113 7157 8125 7191
rect 8159 7188 8171 7191
rect 8294 7188 8300 7200
rect 8159 7160 8300 7188
rect 8159 7157 8171 7160
rect 8113 7151 8171 7157
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 9122 7148 9128 7200
rect 9180 7188 9186 7200
rect 9401 7191 9459 7197
rect 9401 7188 9413 7191
rect 9180 7160 9413 7188
rect 9180 7148 9186 7160
rect 9401 7157 9413 7160
rect 9447 7157 9459 7191
rect 9401 7151 9459 7157
rect 10321 7191 10379 7197
rect 10321 7157 10333 7191
rect 10367 7188 10379 7191
rect 10502 7188 10508 7200
rect 10367 7160 10508 7188
rect 10367 7157 10379 7160
rect 10321 7151 10379 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 1104 7098 14812 7120
rect 1104 7046 5579 7098
rect 5631 7046 5643 7098
rect 5695 7046 5707 7098
rect 5759 7046 5771 7098
rect 5823 7046 10176 7098
rect 10228 7046 10240 7098
rect 10292 7046 10304 7098
rect 10356 7046 10368 7098
rect 10420 7046 14812 7098
rect 1104 7024 14812 7046
rect 2406 6944 2412 6996
rect 2464 6984 2470 6996
rect 4062 6984 4068 6996
rect 2464 6956 4068 6984
rect 2464 6944 2470 6956
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 4890 6944 4896 6996
rect 4948 6984 4954 6996
rect 8849 6987 8907 6993
rect 8849 6984 8861 6987
rect 4948 6956 8861 6984
rect 4948 6944 4954 6956
rect 8849 6953 8861 6956
rect 8895 6984 8907 6987
rect 11422 6984 11428 6996
rect 8895 6956 11428 6984
rect 8895 6953 8907 6956
rect 8849 6947 8907 6953
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 13136 6956 13553 6984
rect 13136 6944 13142 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13541 6947 13599 6953
rect 2777 6919 2835 6925
rect 2777 6885 2789 6919
rect 2823 6916 2835 6919
rect 4430 6916 4436 6928
rect 2823 6888 4436 6916
rect 2823 6885 2835 6888
rect 2777 6879 2835 6885
rect 4430 6876 4436 6888
rect 4488 6876 4494 6928
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 4065 6851 4123 6857
rect 1443 6820 4016 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2498 6740 2504 6792
rect 2556 6780 2562 6792
rect 2869 6783 2927 6789
rect 2869 6780 2881 6783
rect 2556 6752 2881 6780
rect 2556 6740 2562 6752
rect 2869 6749 2881 6752
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6780 3111 6783
rect 3786 6780 3792 6792
rect 3099 6752 3792 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 3988 6780 4016 6820
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4908 6848 4936 6944
rect 7006 6916 7012 6928
rect 4111 6820 4936 6848
rect 5000 6888 7012 6916
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 5000 6780 5028 6888
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 8205 6919 8263 6925
rect 8205 6916 8217 6919
rect 8168 6888 8217 6916
rect 8168 6876 8174 6888
rect 8205 6885 8217 6888
rect 8251 6885 8263 6919
rect 8205 6879 8263 6885
rect 12428 6919 12486 6925
rect 12428 6885 12440 6919
rect 12474 6916 12486 6919
rect 12986 6916 12992 6928
rect 12474 6888 12992 6916
rect 12474 6885 12486 6888
rect 12428 6879 12486 6885
rect 12986 6876 12992 6888
rect 13044 6876 13050 6928
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 6641 6851 6699 6857
rect 6641 6848 6653 6851
rect 6595 6820 6653 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 6641 6817 6653 6820
rect 6687 6817 6699 6851
rect 6641 6811 6699 6817
rect 3988 6752 5028 6780
rect 5368 6780 5396 6811
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 7558 6848 7564 6860
rect 6880 6820 7564 6848
rect 6880 6808 6886 6820
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 8128 6780 8156 6876
rect 9490 6848 9496 6860
rect 8956 6820 9496 6848
rect 8956 6792 8984 6820
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 10042 6848 10048 6860
rect 9640 6820 10048 6848
rect 9640 6808 9646 6820
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10220 6851 10278 6857
rect 10220 6817 10232 6851
rect 10266 6848 10278 6851
rect 10778 6848 10784 6860
rect 10266 6820 10784 6848
rect 10266 6817 10278 6820
rect 10220 6811 10278 6817
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 8938 6780 8944 6792
rect 5368 6752 8156 6780
rect 8899 6752 8944 6780
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9306 6780 9312 6792
rect 9171 6752 9312 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 6549 6715 6607 6721
rect 6549 6712 6561 6715
rect 4764 6684 6561 6712
rect 4764 6672 4770 6684
rect 6549 6681 6561 6684
rect 6595 6681 6607 6715
rect 6549 6675 6607 6681
rect 8202 6672 8208 6724
rect 8260 6712 8266 6724
rect 9140 6712 9168 6743
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6749 12219 6783
rect 12161 6743 12219 6749
rect 8260 6684 9168 6712
rect 8260 6672 8266 6684
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 3050 6644 3056 6656
rect 2455 6616 3056 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 4249 6647 4307 6653
rect 4249 6613 4261 6647
rect 4295 6644 4307 6647
rect 5074 6644 5080 6656
rect 4295 6616 5080 6644
rect 4295 6613 4307 6616
rect 4249 6607 4307 6613
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5902 6644 5908 6656
rect 5215 6616 5908 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 8478 6644 8484 6656
rect 8439 6616 8484 6644
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 9968 6644 9996 6743
rect 10962 6672 10968 6724
rect 11020 6712 11026 6724
rect 11330 6712 11336 6724
rect 11020 6684 11336 6712
rect 11020 6672 11026 6684
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 12176 6644 12204 6743
rect 9548 6616 12204 6644
rect 9548 6604 9554 6616
rect 1104 6554 14812 6576
rect 1104 6502 3280 6554
rect 3332 6502 3344 6554
rect 3396 6502 3408 6554
rect 3460 6502 3472 6554
rect 3524 6502 7878 6554
rect 7930 6502 7942 6554
rect 7994 6502 8006 6554
rect 8058 6502 8070 6554
rect 8122 6502 12475 6554
rect 12527 6502 12539 6554
rect 12591 6502 12603 6554
rect 12655 6502 12667 6554
rect 12719 6502 14812 6554
rect 1104 6480 14812 6502
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 3789 6443 3847 6449
rect 3789 6440 3801 6443
rect 2740 6412 3801 6440
rect 2740 6400 2746 6412
rect 3436 6384 3464 6412
rect 3789 6409 3801 6412
rect 3835 6409 3847 6443
rect 3789 6403 3847 6409
rect 1302 6332 1308 6384
rect 1360 6372 1366 6384
rect 1946 6372 1952 6384
rect 1360 6344 1952 6372
rect 1360 6332 1366 6344
rect 1946 6332 1952 6344
rect 2004 6332 2010 6384
rect 3418 6332 3424 6384
rect 3476 6332 3482 6384
rect 2406 6304 2412 6316
rect 2367 6276 2412 6304
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 3602 6264 3608 6316
rect 3660 6264 3666 6316
rect 3804 6304 3832 6403
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 6641 6443 6699 6449
rect 6641 6440 6653 6443
rect 6512 6412 6653 6440
rect 6512 6400 6518 6412
rect 6641 6409 6653 6412
rect 6687 6440 6699 6443
rect 9030 6440 9036 6452
rect 6687 6412 9036 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 9364 6412 10885 6440
rect 9364 6400 9370 6412
rect 10873 6409 10885 6412
rect 10919 6409 10931 6443
rect 10873 6403 10931 6409
rect 12621 6443 12679 6449
rect 12621 6409 12633 6443
rect 12667 6440 12679 6443
rect 12894 6440 12900 6452
rect 12667 6412 12900 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 12894 6400 12900 6412
rect 12952 6400 12958 6452
rect 4430 6372 4436 6384
rect 4391 6344 4436 6372
rect 4430 6332 4436 6344
rect 4488 6332 4494 6384
rect 4798 6332 4804 6384
rect 4856 6372 4862 6384
rect 4856 6344 5304 6372
rect 4856 6332 4862 6344
rect 5276 6313 5304 6344
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 8938 6372 8944 6384
rect 8352 6344 8944 6372
rect 8352 6332 8358 6344
rect 8938 6332 8944 6344
rect 8996 6332 9002 6384
rect 4985 6307 5043 6313
rect 4985 6304 4997 6307
rect 3804 6276 4997 6304
rect 4985 6273 4997 6276
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6273 5319 6307
rect 9490 6304 9496 6316
rect 9451 6276 9496 6304
rect 5261 6267 5319 6273
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 13170 6304 13176 6316
rect 13044 6276 13176 6304
rect 13044 6264 13050 6276
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 2676 6171 2734 6177
rect 2676 6137 2688 6171
rect 2722 6168 2734 6171
rect 3620 6168 3648 6264
rect 4338 6196 4344 6248
rect 4396 6236 4402 6248
rect 4893 6239 4951 6245
rect 4893 6236 4905 6239
rect 4396 6208 4905 6236
rect 4396 6196 4402 6208
rect 4893 6205 4905 6208
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6236 7343 6239
rect 9508 6236 9536 6264
rect 7331 6208 9536 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 13081 6239 13139 6245
rect 13081 6236 13093 6239
rect 9640 6208 13093 6236
rect 9640 6196 9646 6208
rect 13081 6205 13093 6208
rect 13127 6205 13139 6239
rect 13081 6199 13139 6205
rect 3970 6168 3976 6180
rect 2722 6140 3976 6168
rect 2722 6137 2734 6140
rect 2676 6131 2734 6137
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 5528 6171 5586 6177
rect 5528 6137 5540 6171
rect 5574 6168 5586 6171
rect 7552 6171 7610 6177
rect 5574 6140 7512 6168
rect 5574 6137 5586 6140
rect 5528 6131 5586 6137
rect 1397 6103 1455 6109
rect 1397 6069 1409 6103
rect 1443 6100 1455 6103
rect 3142 6100 3148 6112
rect 1443 6072 3148 6100
rect 1443 6069 1455 6072
rect 1397 6063 1455 6069
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 4614 6100 4620 6112
rect 4120 6072 4620 6100
rect 4120 6060 4126 6072
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 4798 6100 4804 6112
rect 4759 6072 4804 6100
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5994 6060 6000 6112
rect 6052 6100 6058 6112
rect 6270 6100 6276 6112
rect 6052 6072 6276 6100
rect 6052 6060 6058 6072
rect 6270 6060 6276 6072
rect 6328 6060 6334 6112
rect 7484 6100 7512 6140
rect 7552 6137 7564 6171
rect 7598 6168 7610 6171
rect 8202 6168 8208 6180
rect 7598 6140 8208 6168
rect 7598 6137 7610 6140
rect 7552 6131 7610 6137
rect 8202 6128 8208 6140
rect 8260 6128 8266 6180
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 9760 6171 9818 6177
rect 8352 6140 9628 6168
rect 8352 6128 8358 6140
rect 7650 6100 7656 6112
rect 7484 6072 7656 6100
rect 7650 6060 7656 6072
rect 7708 6100 7714 6112
rect 8665 6103 8723 6109
rect 8665 6100 8677 6103
rect 7708 6072 8677 6100
rect 7708 6060 7714 6072
rect 8665 6069 8677 6072
rect 8711 6069 8723 6103
rect 9600 6100 9628 6140
rect 9760 6137 9772 6171
rect 9806 6168 9818 6171
rect 11054 6168 11060 6180
rect 9806 6140 11060 6168
rect 9806 6137 9818 6140
rect 9760 6131 9818 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 12989 6171 13047 6177
rect 12989 6137 13001 6171
rect 13035 6168 13047 6171
rect 13630 6168 13636 6180
rect 13035 6140 13636 6168
rect 13035 6137 13047 6140
rect 12989 6131 13047 6137
rect 13630 6128 13636 6140
rect 13688 6128 13694 6180
rect 9950 6100 9956 6112
rect 9600 6072 9956 6100
rect 8665 6063 8723 6069
rect 9950 6060 9956 6072
rect 10008 6100 10014 6112
rect 10870 6100 10876 6112
rect 10008 6072 10876 6100
rect 10008 6060 10014 6072
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 12894 6060 12900 6112
rect 12952 6100 12958 6112
rect 13354 6100 13360 6112
rect 12952 6072 13360 6100
rect 12952 6060 12958 6072
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 1104 6010 14812 6032
rect 1104 5958 5579 6010
rect 5631 5958 5643 6010
rect 5695 5958 5707 6010
rect 5759 5958 5771 6010
rect 5823 5958 10176 6010
rect 10228 5958 10240 6010
rect 10292 5958 10304 6010
rect 10356 5958 10368 6010
rect 10420 5958 14812 6010
rect 1104 5936 14812 5958
rect 8294 5896 8300 5908
rect 1780 5868 8300 5896
rect 934 5720 940 5772
rect 992 5760 998 5772
rect 1780 5769 1808 5868
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 9950 5896 9956 5908
rect 8435 5868 9956 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 11054 5896 11060 5908
rect 11015 5868 11060 5896
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 12621 5899 12679 5905
rect 12621 5865 12633 5899
rect 12667 5896 12679 5899
rect 12802 5896 12808 5908
rect 12667 5868 12808 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 4890 5828 4896 5840
rect 2823 5800 4896 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 4890 5788 4896 5800
rect 4948 5788 4954 5840
rect 5620 5831 5678 5837
rect 5620 5797 5632 5831
rect 5666 5828 5678 5831
rect 6454 5828 6460 5840
rect 5666 5800 6460 5828
rect 5666 5797 5678 5800
rect 5620 5791 5678 5797
rect 6454 5788 6460 5800
rect 6512 5828 6518 5840
rect 7006 5828 7012 5840
rect 6512 5800 7012 5828
rect 6512 5788 6518 5800
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 8481 5831 8539 5837
rect 8481 5797 8493 5831
rect 8527 5828 8539 5831
rect 9214 5828 9220 5840
rect 8527 5800 9220 5828
rect 8527 5797 8539 5800
rect 8481 5791 8539 5797
rect 9214 5788 9220 5800
rect 9272 5788 9278 5840
rect 11072 5828 11100 5856
rect 9600 5800 11100 5828
rect 1397 5763 1455 5769
rect 1397 5760 1409 5763
rect 992 5732 1409 5760
rect 992 5720 998 5732
rect 1397 5729 1409 5732
rect 1443 5729 1455 5763
rect 1397 5723 1455 5729
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5729 1823 5763
rect 3418 5760 3424 5772
rect 1765 5723 1823 5729
rect 2976 5732 3424 5760
rect 2866 5692 2872 5704
rect 2827 5664 2872 5692
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 2976 5701 3004 5732
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 6730 5760 6736 5772
rect 4111 5732 6736 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 5258 5692 5264 5704
rect 4212 5664 5264 5692
rect 4212 5652 4218 5664
rect 5258 5652 5264 5664
rect 5316 5692 5322 5704
rect 5353 5695 5411 5701
rect 5353 5692 5365 5695
rect 5316 5664 5365 5692
rect 5316 5652 5322 5664
rect 5353 5661 5365 5664
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8570 5692 8576 5704
rect 8352 5664 8576 5692
rect 8352 5652 8358 5664
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5692 8723 5695
rect 9600 5692 9628 5800
rect 12250 5788 12256 5840
rect 12308 5828 12314 5840
rect 12989 5831 13047 5837
rect 12989 5828 13001 5831
rect 12308 5800 13001 5828
rect 12308 5788 12314 5800
rect 12989 5797 13001 5800
rect 13035 5797 13047 5831
rect 12989 5791 13047 5797
rect 9944 5763 10002 5769
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 10962 5760 10968 5772
rect 9990 5732 10968 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 8711 5664 9628 5692
rect 9677 5695 9735 5701
rect 8711 5661 8723 5664
rect 8665 5655 8723 5661
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 1946 5624 1952 5636
rect 1907 5596 1952 5624
rect 1946 5584 1952 5596
rect 2004 5584 2010 5636
rect 2317 5627 2375 5633
rect 2317 5593 2329 5627
rect 2363 5624 2375 5627
rect 2363 5596 5396 5624
rect 2363 5593 2375 5596
rect 2317 5587 2375 5593
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 1670 5556 1676 5568
rect 1627 5528 1676 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 2406 5556 2412 5568
rect 2367 5528 2412 5556
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 4154 5516 4160 5568
rect 4212 5556 4218 5568
rect 4249 5559 4307 5565
rect 4249 5556 4261 5559
rect 4212 5528 4261 5556
rect 4212 5516 4218 5528
rect 4249 5525 4261 5528
rect 4295 5525 4307 5559
rect 5368 5556 5396 5596
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 9692 5624 9720 5655
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 12308 5664 13093 5692
rect 12308 5652 12314 5664
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13170 5652 13176 5704
rect 13228 5692 13234 5704
rect 13228 5664 13273 5692
rect 13228 5652 13234 5664
rect 9548 5596 9720 5624
rect 9548 5584 9554 5596
rect 6086 5556 6092 5568
rect 5368 5528 6092 5556
rect 4249 5519 4307 5525
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 6730 5556 6736 5568
rect 6691 5528 6736 5556
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 8021 5559 8079 5565
rect 8021 5525 8033 5559
rect 8067 5556 8079 5559
rect 8202 5556 8208 5568
rect 8067 5528 8208 5556
rect 8067 5525 8079 5528
rect 8021 5519 8079 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 8662 5516 8668 5568
rect 8720 5556 8726 5568
rect 11882 5556 11888 5568
rect 8720 5528 11888 5556
rect 8720 5516 8726 5528
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 1104 5466 14812 5488
rect 1104 5414 3280 5466
rect 3332 5414 3344 5466
rect 3396 5414 3408 5466
rect 3460 5414 3472 5466
rect 3524 5414 7878 5466
rect 7930 5414 7942 5466
rect 7994 5414 8006 5466
rect 8058 5414 8070 5466
rect 8122 5414 12475 5466
rect 12527 5414 12539 5466
rect 12591 5414 12603 5466
rect 12655 5414 12667 5466
rect 12719 5414 14812 5466
rect 1104 5392 14812 5414
rect 1394 5352 1400 5364
rect 1355 5324 1400 5352
rect 1394 5312 1400 5324
rect 1452 5312 1458 5364
rect 3329 5355 3387 5361
rect 3329 5321 3341 5355
rect 3375 5352 3387 5355
rect 4798 5352 4804 5364
rect 3375 5324 4804 5352
rect 3375 5321 3387 5324
rect 3329 5315 3387 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 4948 5324 4993 5352
rect 4948 5312 4954 5324
rect 5258 5312 5264 5364
rect 5316 5352 5322 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 5316 5324 6469 5352
rect 5316 5312 5322 5324
rect 6457 5321 6469 5324
rect 6503 5352 6515 5355
rect 6822 5352 6828 5364
rect 6503 5324 6828 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 9232 5324 9444 5352
rect 6730 5284 6736 5296
rect 2884 5256 6736 5284
rect 1946 5216 1952 5228
rect 1907 5188 1952 5216
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 2222 5176 2228 5228
rect 2280 5216 2286 5228
rect 2498 5216 2504 5228
rect 2280 5188 2504 5216
rect 2280 5176 2286 5188
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 2884 5225 2912 5256
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 7101 5287 7159 5293
rect 7101 5253 7113 5287
rect 7147 5284 7159 5287
rect 9232 5284 9260 5324
rect 7147 5256 9260 5284
rect 9416 5284 9444 5324
rect 9490 5312 9496 5364
rect 9548 5352 9554 5364
rect 9585 5355 9643 5361
rect 9585 5352 9597 5355
rect 9548 5324 9597 5352
rect 9548 5312 9554 5324
rect 9585 5321 9597 5324
rect 9631 5321 9643 5355
rect 9950 5352 9956 5364
rect 9911 5324 9956 5352
rect 9585 5315 9643 5321
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 10502 5352 10508 5364
rect 10376 5324 10508 5352
rect 10376 5312 10382 5324
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 11054 5284 11060 5296
rect 9416 5256 11060 5284
rect 7147 5253 7159 5256
rect 7101 5247 7159 5253
rect 11054 5244 11060 5256
rect 11112 5244 11118 5296
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5185 2927 5219
rect 3510 5216 3516 5228
rect 2869 5179 2927 5185
rect 2976 5188 3516 5216
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5148 1823 5151
rect 2976 5148 3004 5188
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 3694 5176 3700 5228
rect 3752 5216 3758 5228
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 3752 5188 3801 5216
rect 3752 5176 3758 5188
rect 3789 5185 3801 5188
rect 3835 5185 3847 5219
rect 3970 5216 3976 5228
rect 3931 5188 3976 5216
rect 3789 5179 3847 5185
rect 3970 5176 3976 5188
rect 4028 5216 4034 5228
rect 4614 5216 4620 5228
rect 4028 5188 4620 5216
rect 4028 5176 4034 5188
rect 4614 5176 4620 5188
rect 4672 5216 4678 5228
rect 5166 5216 5172 5228
rect 4672 5188 5172 5216
rect 4672 5176 4678 5188
rect 5166 5176 5172 5188
rect 5224 5216 5230 5228
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 5224 5188 5457 5216
rect 5224 5176 5230 5188
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 8481 5219 8539 5225
rect 8481 5216 8493 5219
rect 7340 5188 8493 5216
rect 7340 5176 7346 5188
rect 8481 5185 8493 5188
rect 8527 5185 8539 5219
rect 8481 5179 8539 5185
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5216 8723 5219
rect 9214 5216 9220 5228
rect 8711 5188 9220 5216
rect 8711 5185 8723 5188
rect 8665 5179 8723 5185
rect 4430 5148 4436 5160
rect 1811 5120 3004 5148
rect 3068 5120 4436 5148
rect 1811 5117 1823 5120
rect 1765 5111 1823 5117
rect 3068 5080 3096 5120
rect 4430 5108 4436 5120
rect 4488 5108 4494 5160
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5350 5148 5356 5160
rect 5307 5120 5356 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 6641 5151 6699 5157
rect 6641 5148 6653 5151
rect 5960 5120 6653 5148
rect 5960 5108 5966 5120
rect 6641 5117 6653 5120
rect 6687 5117 6699 5151
rect 6641 5111 6699 5117
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5148 6975 5151
rect 6963 5120 7328 5148
rect 6963 5117 6975 5120
rect 6917 5111 6975 5117
rect 7300 5092 7328 5120
rect 2240 5052 3096 5080
rect 1854 4972 1860 5024
rect 1912 5012 1918 5024
rect 2240 5021 2268 5052
rect 3142 5040 3148 5092
rect 3200 5080 3206 5092
rect 3697 5083 3755 5089
rect 3697 5080 3709 5083
rect 3200 5052 3709 5080
rect 3200 5040 3206 5052
rect 3697 5049 3709 5052
rect 3743 5049 3755 5083
rect 3697 5043 3755 5049
rect 4890 5040 4896 5092
rect 4948 5080 4954 5092
rect 7190 5080 7196 5092
rect 4948 5052 7196 5080
rect 4948 5040 4954 5052
rect 7190 5040 7196 5052
rect 7248 5040 7254 5092
rect 7282 5040 7288 5092
rect 7340 5040 7346 5092
rect 7668 5052 8156 5080
rect 2225 5015 2283 5021
rect 1912 4984 1957 5012
rect 1912 4972 1918 4984
rect 2225 4981 2237 5015
rect 2271 4981 2283 5015
rect 2225 4975 2283 4981
rect 2498 4972 2504 5024
rect 2556 5012 2562 5024
rect 2593 5015 2651 5021
rect 2593 5012 2605 5015
rect 2556 4984 2605 5012
rect 2556 4972 2562 4984
rect 2593 4981 2605 4984
rect 2639 4981 2651 5015
rect 2593 4975 2651 4981
rect 2685 5015 2743 5021
rect 2685 4981 2697 5015
rect 2731 5012 2743 5015
rect 4798 5012 4804 5024
rect 2731 4984 4804 5012
rect 2731 4981 2743 4984
rect 2685 4975 2743 4981
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 5408 4984 5453 5012
rect 5408 4972 5414 4984
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 7668 5012 7696 5052
rect 6512 4984 7696 5012
rect 6512 4972 6518 4984
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7800 4984 8033 5012
rect 7800 4972 7806 4984
rect 8021 4981 8033 4984
rect 8067 4981 8079 5015
rect 8128 5012 8156 5052
rect 8294 5040 8300 5092
rect 8352 5080 8358 5092
rect 8389 5083 8447 5089
rect 8389 5080 8401 5083
rect 8352 5052 8401 5080
rect 8352 5040 8358 5052
rect 8389 5049 8401 5052
rect 8435 5049 8447 5083
rect 8496 5080 8524 5179
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 9582 5176 9588 5228
rect 9640 5216 9646 5228
rect 10226 5216 10232 5228
rect 9640 5188 10232 5216
rect 9640 5176 9646 5188
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 10962 5216 10968 5228
rect 10643 5188 10968 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 13170 5216 13176 5228
rect 13131 5188 13176 5216
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 9766 5148 9772 5160
rect 9727 5120 9772 5148
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 10318 5108 10324 5160
rect 10376 5148 10382 5160
rect 10413 5151 10471 5157
rect 10413 5148 10425 5151
rect 10376 5120 10425 5148
rect 10376 5108 10382 5120
rect 10413 5117 10425 5120
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12492 5120 12909 5148
rect 12492 5108 12498 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 9950 5080 9956 5092
rect 8496 5052 9956 5080
rect 8389 5043 8447 5049
rect 9950 5040 9956 5052
rect 10008 5040 10014 5092
rect 10134 5040 10140 5092
rect 10192 5040 10198 5092
rect 11330 5040 11336 5092
rect 11388 5080 11394 5092
rect 12989 5083 13047 5089
rect 12989 5080 13001 5083
rect 11388 5052 13001 5080
rect 11388 5040 11394 5052
rect 12989 5049 13001 5052
rect 13035 5049 13047 5083
rect 12989 5043 13047 5049
rect 10152 5012 10180 5040
rect 8128 4984 10180 5012
rect 10321 5015 10379 5021
rect 8021 4975 8079 4981
rect 10321 4981 10333 5015
rect 10367 5012 10379 5015
rect 10502 5012 10508 5024
rect 10367 4984 10508 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 10502 4972 10508 4984
rect 10560 4972 10566 5024
rect 12526 5012 12532 5024
rect 12487 4984 12532 5012
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 1104 4922 14812 4944
rect 1104 4870 5579 4922
rect 5631 4870 5643 4922
rect 5695 4870 5707 4922
rect 5759 4870 5771 4922
rect 5823 4870 10176 4922
rect 10228 4870 10240 4922
rect 10292 4870 10304 4922
rect 10356 4870 10368 4922
rect 10420 4870 14812 4922
rect 1104 4848 14812 4870
rect 1397 4811 1455 4817
rect 1397 4777 1409 4811
rect 1443 4808 1455 4811
rect 1854 4808 1860 4820
rect 1443 4780 1860 4808
rect 1443 4777 1455 4780
rect 1397 4771 1455 4777
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 2823 4780 5120 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 1118 4700 1124 4752
rect 1176 4740 1182 4752
rect 2590 4740 2596 4752
rect 1176 4712 2596 4740
rect 1176 4700 1182 4712
rect 2590 4700 2596 4712
rect 2648 4700 2654 4752
rect 4062 4740 4068 4752
rect 3068 4712 4068 4740
rect 1394 4632 1400 4684
rect 1452 4672 1458 4684
rect 1765 4675 1823 4681
rect 1765 4672 1777 4675
rect 1452 4644 1777 4672
rect 1452 4632 1458 4644
rect 1765 4641 1777 4644
rect 1811 4641 1823 4675
rect 1765 4635 1823 4641
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 2682 4672 2688 4684
rect 1903 4644 2688 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4604 2099 4607
rect 2498 4604 2504 4616
rect 2087 4576 2504 4604
rect 2087 4573 2099 4576
rect 2041 4567 2099 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 2590 4564 2596 4616
rect 2648 4604 2654 4616
rect 3068 4613 3096 4712
rect 4062 4700 4068 4712
rect 4120 4740 4126 4752
rect 4310 4743 4368 4749
rect 4310 4740 4322 4743
rect 4120 4712 4322 4740
rect 4120 4700 4126 4712
rect 4310 4709 4322 4712
rect 4356 4709 4368 4743
rect 5092 4740 5120 4780
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5445 4811 5503 4817
rect 5445 4808 5457 4811
rect 5224 4780 5457 4808
rect 5224 4768 5230 4780
rect 5445 4777 5457 4780
rect 5491 4777 5503 4811
rect 7466 4808 7472 4820
rect 5445 4771 5503 4777
rect 5920 4780 7472 4808
rect 5920 4752 5948 4780
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7742 4808 7748 4820
rect 7703 4780 7748 4808
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 7837 4811 7895 4817
rect 7837 4777 7849 4811
rect 7883 4808 7895 4811
rect 8478 4808 8484 4820
rect 7883 4780 8484 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 8938 4768 8944 4820
rect 8996 4808 9002 4820
rect 9306 4808 9312 4820
rect 8996 4780 9312 4808
rect 8996 4768 9002 4780
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 10321 4811 10379 4817
rect 10321 4777 10333 4811
rect 10367 4808 10379 4811
rect 10502 4808 10508 4820
rect 10367 4780 10508 4808
rect 10367 4777 10379 4780
rect 10321 4771 10379 4777
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 10686 4808 10692 4820
rect 10647 4780 10692 4808
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 11146 4768 11152 4820
rect 11204 4808 11210 4820
rect 12069 4811 12127 4817
rect 12069 4808 12081 4811
rect 11204 4780 12081 4808
rect 11204 4768 11210 4780
rect 12069 4777 12081 4780
rect 12115 4777 12127 4811
rect 12526 4808 12532 4820
rect 12487 4780 12532 4808
rect 12069 4771 12127 4777
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 5902 4740 5908 4752
rect 5092 4712 5908 4740
rect 4310 4703 4368 4709
rect 5902 4700 5908 4712
rect 5960 4700 5966 4752
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 6052 4712 10732 4740
rect 6052 4700 6058 4712
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 3878 4672 3884 4684
rect 3283 4644 3884 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 6270 4672 6276 4684
rect 5316 4644 6276 4672
rect 5316 4632 5322 4644
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 10410 4672 10416 4684
rect 6380 4644 10416 4672
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2648 4576 2881 4604
rect 2648 4564 2654 4576
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 842 4496 848 4548
rect 900 4536 906 4548
rect 3436 4536 3464 4567
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 4028 4576 4077 4604
rect 4028 4564 4034 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 5810 4564 5816 4616
rect 5868 4604 5874 4616
rect 6380 4604 6408 4644
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 5868 4576 6408 4604
rect 5868 4564 5874 4576
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7708 4576 7941 4604
rect 7708 4564 7714 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 900 4508 3464 4536
rect 6457 4539 6515 4545
rect 900 4496 906 4508
rect 6457 4505 6469 4539
rect 6503 4536 6515 4539
rect 9582 4536 9588 4548
rect 6503 4508 9588 4536
rect 6503 4505 6515 4508
rect 6457 4499 6515 4505
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 2409 4471 2467 4477
rect 2409 4437 2421 4471
rect 2455 4468 2467 4471
rect 4246 4468 4252 4480
rect 2455 4440 4252 4468
rect 2455 4437 2467 4440
rect 2409 4431 2467 4437
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 7377 4471 7435 4477
rect 7377 4468 7389 4471
rect 7340 4440 7389 4468
rect 7340 4428 7346 4440
rect 7377 4437 7389 4440
rect 7423 4437 7435 4471
rect 10704 4468 10732 4712
rect 10778 4700 10784 4752
rect 10836 4740 10842 4752
rect 10836 4712 10916 4740
rect 10836 4700 10842 4712
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10888 4604 10916 4712
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 11204 4644 12449 4672
rect 11204 4632 11210 4644
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 12437 4635 12495 4641
rect 12986 4632 12992 4684
rect 13044 4672 13050 4684
rect 13722 4672 13728 4684
rect 13044 4644 13728 4672
rect 13044 4632 13050 4644
rect 13722 4632 13728 4644
rect 13780 4632 13786 4684
rect 10965 4607 11023 4613
rect 10965 4604 10977 4607
rect 10888 4576 10977 4604
rect 10781 4567 10839 4573
rect 10965 4573 10977 4576
rect 11011 4604 11023 4607
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 11011 4576 12633 4604
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 12621 4573 12633 4576
rect 12667 4573 12679 4607
rect 12621 4567 12679 4573
rect 10796 4536 10824 4567
rect 11606 4536 11612 4548
rect 10796 4508 11612 4536
rect 11606 4496 11612 4508
rect 11664 4496 11670 4548
rect 11146 4468 11152 4480
rect 10704 4440 11152 4468
rect 7377 4431 7435 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 1104 4378 14812 4400
rect 1104 4326 3280 4378
rect 3332 4326 3344 4378
rect 3396 4326 3408 4378
rect 3460 4326 3472 4378
rect 3524 4326 7878 4378
rect 7930 4326 7942 4378
rect 7994 4326 8006 4378
rect 8058 4326 8070 4378
rect 8122 4326 12475 4378
rect 12527 4326 12539 4378
rect 12591 4326 12603 4378
rect 12655 4326 12667 4378
rect 12719 4326 14812 4378
rect 1104 4304 14812 4326
rect 1946 4224 1952 4276
rect 2004 4264 2010 4276
rect 2004 4236 2636 4264
rect 2004 4224 2010 4236
rect 1486 4156 1492 4208
rect 1544 4196 1550 4208
rect 2225 4199 2283 4205
rect 2225 4196 2237 4199
rect 1544 4168 2237 4196
rect 1544 4156 1550 4168
rect 2225 4165 2237 4168
rect 2271 4165 2283 4199
rect 2608 4196 2636 4236
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 2740 4236 4364 4264
rect 2740 4224 2746 4236
rect 2608 4168 2820 4196
rect 2225 4159 2283 4165
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 1949 4131 2007 4137
rect 1949 4128 1961 4131
rect 1820 4100 1961 4128
rect 1820 4088 1826 4100
rect 1949 4097 1961 4100
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2792 4137 2820 4168
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2188 4100 2697 4128
rect 2188 4088 2194 4100
rect 2685 4097 2697 4100
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 4120 4100 4261 4128
rect 4120 4088 4126 4100
rect 4249 4097 4261 4100
rect 4295 4097 4307 4131
rect 4336 4128 4364 4236
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 9490 4264 9496 4276
rect 7064 4236 7788 4264
rect 7064 4224 7070 4236
rect 5074 4156 5080 4208
rect 5132 4196 5138 4208
rect 5132 4168 6960 4196
rect 5132 4156 5138 4168
rect 6178 4128 6184 4140
rect 4336 4100 6184 4128
rect 4249 4091 4307 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 6932 4128 6960 4168
rect 6932 4100 7236 4128
rect 2222 4060 2228 4072
rect 1780 4032 2228 4060
rect 1780 4001 1808 4032
rect 2222 4020 2228 4032
rect 2280 4020 2286 4072
rect 3050 4060 3056 4072
rect 3011 4032 3056 4060
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4060 4215 4063
rect 4338 4060 4344 4072
rect 4203 4032 4344 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 4338 4020 4344 4032
rect 4396 4020 4402 4072
rect 4525 4063 4583 4069
rect 4525 4029 4537 4063
rect 4571 4060 4583 4063
rect 5074 4060 5080 4072
rect 4571 4032 5080 4060
rect 4571 4029 4583 4032
rect 4525 4023 4583 4029
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5445 4063 5503 4069
rect 5445 4060 5457 4063
rect 5316 4032 5457 4060
rect 5316 4020 5322 4032
rect 5445 4029 5457 4032
rect 5491 4029 5503 4063
rect 5445 4023 5503 4029
rect 6914 4020 6920 4072
rect 6972 4020 6978 4072
rect 7208 4060 7236 4100
rect 7282 4088 7288 4140
rect 7340 4128 7346 4140
rect 7469 4131 7527 4137
rect 7340 4100 7385 4128
rect 7340 4088 7346 4100
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 7760 4128 7788 4236
rect 8404 4236 9496 4264
rect 8404 4137 8432 4236
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 11330 4264 11336 4276
rect 10468 4236 11336 4264
rect 10468 4224 10474 4236
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 13538 4264 13544 4276
rect 13499 4236 13544 4264
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 12434 4196 12440 4208
rect 9824 4168 12440 4196
rect 9824 4156 9830 4168
rect 12434 4156 12440 4168
rect 12492 4156 12498 4208
rect 7515 4100 7788 4128
rect 8389 4131 8447 4137
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 8389 4097 8401 4131
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10778 4128 10784 4140
rect 10100 4100 10784 4128
rect 10100 4088 10106 4100
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11072 4100 11376 4128
rect 8478 4060 8484 4072
rect 7208 4032 8484 4060
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 8662 4069 8668 4072
rect 8656 4060 8668 4069
rect 8623 4032 8668 4060
rect 8656 4023 8668 4032
rect 8662 4020 8668 4023
rect 8720 4020 8726 4072
rect 9030 4020 9036 4072
rect 9088 4060 9094 4072
rect 11072 4060 11100 4100
rect 9088 4032 11100 4060
rect 9088 4020 9094 4032
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 11241 4063 11299 4069
rect 11241 4060 11253 4063
rect 11204 4032 11253 4060
rect 11204 4020 11210 4032
rect 11241 4029 11253 4032
rect 11287 4029 11299 4063
rect 11348 4060 11376 4100
rect 13357 4063 13415 4069
rect 13357 4060 13369 4063
rect 11348 4032 13369 4060
rect 11241 4023 11299 4029
rect 13357 4029 13369 4032
rect 13403 4029 13415 4063
rect 13357 4023 13415 4029
rect 1765 3995 1823 4001
rect 1765 3961 1777 3995
rect 1811 3961 1823 3995
rect 1765 3955 1823 3961
rect 1946 3952 1952 4004
rect 2004 3992 2010 4004
rect 3329 3995 3387 4001
rect 3329 3992 3341 3995
rect 2004 3964 3341 3992
rect 2004 3952 2010 3964
rect 3329 3961 3341 3964
rect 3375 3961 3387 3995
rect 5721 3995 5779 4001
rect 5721 3992 5733 3995
rect 3329 3955 3387 3961
rect 4356 3964 5733 3992
rect 4356 3936 4384 3964
rect 5721 3961 5733 3964
rect 5767 3961 5779 3995
rect 6932 3992 6960 4020
rect 7193 3995 7251 4001
rect 7193 3992 7205 3995
rect 6932 3964 7205 3992
rect 5721 3955 5779 3961
rect 7193 3961 7205 3964
rect 7239 3961 7251 3995
rect 7193 3955 7251 3961
rect 8938 3952 8944 4004
rect 8996 3992 9002 4004
rect 11790 3992 11796 4004
rect 8996 3964 11796 3992
rect 8996 3952 9002 3964
rect 11790 3952 11796 3964
rect 11848 3952 11854 4004
rect 1394 3924 1400 3936
rect 1355 3896 1400 3924
rect 1394 3884 1400 3896
rect 1452 3884 1458 3936
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3924 1915 3927
rect 2130 3924 2136 3936
rect 1903 3896 2136 3924
rect 1903 3893 1915 3896
rect 1857 3887 1915 3893
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 2590 3924 2596 3936
rect 2551 3896 2596 3924
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 2682 3884 2688 3936
rect 2740 3924 2746 3936
rect 3050 3924 3056 3936
rect 2740 3896 3056 3924
rect 2740 3884 2746 3896
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 3694 3924 3700 3936
rect 3655 3896 3700 3924
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 3844 3896 4077 3924
rect 3844 3884 3850 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 4338 3884 4344 3936
rect 4396 3884 4402 3936
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 4580 3896 4721 3924
rect 4580 3884 4586 3896
rect 4709 3893 4721 3896
rect 4755 3893 4767 3927
rect 4709 3887 4767 3893
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 6825 3927 6883 3933
rect 6825 3924 6837 3927
rect 4856 3896 6837 3924
rect 4856 3884 4862 3896
rect 6825 3893 6837 3896
rect 6871 3893 6883 3927
rect 6825 3887 6883 3893
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 9769 3927 9827 3933
rect 9769 3924 9781 3927
rect 6972 3896 9781 3924
rect 6972 3884 6978 3896
rect 9769 3893 9781 3896
rect 9815 3893 9827 3927
rect 11422 3924 11428 3936
rect 11383 3896 11428 3924
rect 9769 3887 9827 3893
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 1104 3834 14812 3856
rect 1104 3782 5579 3834
rect 5631 3782 5643 3834
rect 5695 3782 5707 3834
rect 5759 3782 5771 3834
rect 5823 3782 10176 3834
rect 10228 3782 10240 3834
rect 10292 3782 10304 3834
rect 10356 3782 10368 3834
rect 10420 3782 14812 3834
rect 1104 3760 14812 3782
rect 290 3680 296 3732
rect 348 3720 354 3732
rect 1946 3720 1952 3732
rect 348 3692 1952 3720
rect 348 3680 354 3692
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2869 3723 2927 3729
rect 2869 3720 2881 3723
rect 2648 3692 2881 3720
rect 2648 3680 2654 3692
rect 2869 3689 2881 3692
rect 2915 3689 2927 3723
rect 2869 3683 2927 3689
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 3237 3723 3295 3729
rect 3237 3720 3249 3723
rect 3108 3692 3249 3720
rect 3108 3680 3114 3692
rect 3237 3689 3249 3692
rect 3283 3689 3295 3723
rect 4062 3720 4068 3732
rect 3237 3683 3295 3689
rect 3620 3692 4068 3720
rect 1664 3655 1722 3661
rect 1664 3621 1676 3655
rect 1710 3652 1722 3655
rect 2682 3652 2688 3664
rect 1710 3624 2688 3652
rect 1710 3621 1722 3624
rect 1664 3615 1722 3621
rect 2682 3612 2688 3624
rect 2740 3612 2746 3664
rect 1946 3544 1952 3596
rect 2004 3584 2010 3596
rect 3329 3587 3387 3593
rect 3329 3584 3341 3587
rect 2004 3556 3341 3584
rect 2004 3544 2010 3556
rect 3329 3553 3341 3556
rect 3375 3553 3387 3587
rect 3620 3584 3648 3692
rect 4062 3680 4068 3692
rect 4120 3720 4126 3732
rect 4798 3720 4804 3732
rect 4120 3692 4804 3720
rect 4120 3680 4126 3692
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 5442 3720 5448 3732
rect 5403 3692 5448 3720
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 9858 3720 9864 3732
rect 5650 3692 9864 3720
rect 3694 3612 3700 3664
rect 3752 3652 3758 3664
rect 4433 3655 4491 3661
rect 4433 3652 4445 3655
rect 3752 3624 4445 3652
rect 3752 3612 3758 3624
rect 4433 3621 4445 3624
rect 4479 3621 4491 3655
rect 4433 3615 4491 3621
rect 4522 3612 4528 3664
rect 4580 3652 4586 3664
rect 5534 3652 5540 3664
rect 4580 3624 4625 3652
rect 5184 3624 5540 3652
rect 4580 3612 4586 3624
rect 3329 3547 3387 3553
rect 3436 3556 3648 3584
rect 3436 3516 3464 3556
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4893 3587 4951 3593
rect 4028 3556 4752 3584
rect 4028 3544 4034 3556
rect 2792 3488 3464 3516
rect 3513 3519 3571 3525
rect 2792 3457 2820 3488
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 3878 3516 3884 3528
rect 3559 3488 3884 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 4614 3516 4620 3528
rect 4575 3488 4620 3516
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 4724 3516 4752 3556
rect 4893 3553 4905 3587
rect 4939 3584 4951 3587
rect 5184 3584 5212 3624
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 4939 3556 5212 3584
rect 5261 3587 5319 3593
rect 4939 3553 4951 3556
rect 4893 3547 4951 3553
rect 5261 3553 5273 3587
rect 5307 3584 5319 3587
rect 5442 3584 5448 3596
rect 5307 3556 5448 3584
rect 5307 3553 5319 3556
rect 5261 3547 5319 3553
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 5650 3593 5678 3692
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 10042 3720 10048 3732
rect 9968 3692 10048 3720
rect 7000 3655 7058 3661
rect 7000 3621 7012 3655
rect 7046 3652 7058 3655
rect 8294 3652 8300 3664
rect 7046 3624 8300 3652
rect 7046 3621 7058 3624
rect 7000 3615 7058 3621
rect 8294 3612 8300 3624
rect 8352 3612 8358 3664
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 9766 3652 9772 3664
rect 8444 3624 9772 3652
rect 8444 3612 8450 3624
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 9968 3661 9996 3692
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 12342 3680 12348 3732
rect 12400 3720 12406 3732
rect 12437 3723 12495 3729
rect 12437 3720 12449 3723
rect 12400 3692 12449 3720
rect 12400 3680 12406 3692
rect 12437 3689 12449 3692
rect 12483 3689 12495 3723
rect 12437 3683 12495 3689
rect 13541 3723 13599 3729
rect 13541 3689 13553 3723
rect 13587 3720 13599 3723
rect 13630 3720 13636 3732
rect 13587 3692 13636 3720
rect 13587 3689 13599 3692
rect 13541 3683 13599 3689
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 9953 3655 10011 3661
rect 9953 3621 9965 3655
rect 9999 3621 10011 3655
rect 9953 3615 10011 3621
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3553 5687 3587
rect 5629 3547 5687 3553
rect 6733 3587 6791 3593
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 6822 3584 6828 3596
rect 6779 3556 6828 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 7558 3544 7564 3596
rect 7616 3584 7622 3596
rect 7616 3556 7788 3584
rect 7616 3544 7622 3556
rect 6362 3516 6368 3528
rect 4724 3488 6368 3516
rect 6362 3476 6368 3488
rect 6420 3476 6426 3528
rect 7760 3516 7788 3556
rect 8202 3544 8208 3596
rect 8260 3584 8266 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 8260 3556 9689 3584
rect 8260 3544 8266 3556
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 9775 3556 9996 3584
rect 9775 3516 9803 3556
rect 7760 3488 9803 3516
rect 9968 3516 9996 3556
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 10100 3556 11161 3584
rect 10100 3544 10106 3556
rect 11149 3553 11161 3556
rect 11195 3553 11207 3587
rect 11149 3547 11207 3553
rect 12253 3587 12311 3593
rect 12253 3553 12265 3587
rect 12299 3553 12311 3587
rect 12253 3547 12311 3553
rect 12268 3516 12296 3547
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 13357 3587 13415 3593
rect 13357 3584 13369 3587
rect 12492 3556 13369 3584
rect 12492 3544 12498 3556
rect 13357 3553 13369 3556
rect 13403 3553 13415 3587
rect 13357 3547 13415 3553
rect 9968 3488 12296 3516
rect 2777 3451 2835 3457
rect 2777 3417 2789 3451
rect 2823 3417 2835 3451
rect 2777 3411 2835 3417
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 4065 3451 4123 3457
rect 4065 3448 4077 3451
rect 2924 3420 4077 3448
rect 2924 3408 2930 3420
rect 4065 3417 4077 3420
rect 4111 3417 4123 3451
rect 6270 3448 6276 3460
rect 4065 3411 4123 3417
rect 4172 3420 6276 3448
rect 3602 3340 3608 3392
rect 3660 3380 3666 3392
rect 4172 3380 4200 3420
rect 6270 3408 6276 3420
rect 6328 3408 6334 3460
rect 9674 3448 9680 3460
rect 8036 3420 9680 3448
rect 3660 3352 4200 3380
rect 3660 3340 3666 3352
rect 4246 3340 4252 3392
rect 4304 3380 4310 3392
rect 4522 3380 4528 3392
rect 4304 3352 4528 3380
rect 4304 3340 4310 3352
rect 4522 3340 4528 3352
rect 4580 3340 4586 3392
rect 4614 3340 4620 3392
rect 4672 3380 4678 3392
rect 4890 3380 4896 3392
rect 4672 3352 4896 3380
rect 4672 3340 4678 3352
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5074 3380 5080 3392
rect 5035 3352 5080 3380
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 5813 3383 5871 3389
rect 5813 3349 5825 3383
rect 5859 3380 5871 3383
rect 8036 3380 8064 3420
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 5859 3352 8064 3380
rect 8113 3383 8171 3389
rect 5859 3349 5871 3352
rect 5813 3343 5871 3349
rect 8113 3349 8125 3383
rect 8159 3380 8171 3383
rect 8202 3380 8208 3392
rect 8159 3352 8208 3380
rect 8159 3349 8171 3352
rect 8113 3343 8171 3349
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 9858 3340 9864 3392
rect 9916 3380 9922 3392
rect 10594 3380 10600 3392
rect 9916 3352 10600 3380
rect 9916 3340 9922 3352
rect 10594 3340 10600 3352
rect 10652 3340 10658 3392
rect 11333 3383 11391 3389
rect 11333 3349 11345 3383
rect 11379 3380 11391 3383
rect 11514 3380 11520 3392
rect 11379 3352 11520 3380
rect 11379 3349 11391 3352
rect 11333 3343 11391 3349
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 1104 3290 14812 3312
rect 1104 3238 3280 3290
rect 3332 3238 3344 3290
rect 3396 3238 3408 3290
rect 3460 3238 3472 3290
rect 3524 3238 7878 3290
rect 7930 3238 7942 3290
rect 7994 3238 8006 3290
rect 8058 3238 8070 3290
rect 8122 3238 12475 3290
rect 12527 3238 12539 3290
rect 12591 3238 12603 3290
rect 12655 3238 12667 3290
rect 12719 3238 14812 3290
rect 1104 3216 14812 3238
rect 2498 3136 2504 3188
rect 2556 3176 2562 3188
rect 10134 3176 10140 3188
rect 2556 3148 10140 3176
rect 2556 3136 2562 3148
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 13541 3179 13599 3185
rect 13541 3145 13553 3179
rect 13587 3176 13599 3179
rect 13722 3176 13728 3188
rect 13587 3148 13728 3176
rect 13587 3145 13599 3148
rect 13541 3139 13599 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 5350 3108 5356 3120
rect 4387 3080 5356 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 5350 3068 5356 3080
rect 5408 3068 5414 3120
rect 9217 3111 9275 3117
rect 9217 3077 9229 3111
rect 9263 3108 9275 3111
rect 15746 3108 15752 3120
rect 9263 3080 15752 3108
rect 9263 3077 9275 3080
rect 9217 3071 9275 3077
rect 15746 3068 15752 3080
rect 15804 3068 15810 3120
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 4488 3012 4844 3040
rect 4488 3000 4494 3012
rect 1664 2975 1722 2981
rect 1664 2941 1676 2975
rect 1710 2972 1722 2975
rect 2406 2972 2412 2984
rect 1710 2944 2412 2972
rect 1710 2941 1722 2944
rect 1664 2935 1722 2941
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 2866 2972 2872 2984
rect 2827 2944 2872 2972
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 4338 2972 4344 2984
rect 3068 2944 4344 2972
rect 1394 2864 1400 2916
rect 1452 2904 1458 2916
rect 3068 2904 3096 2944
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 4522 2932 4528 2984
rect 4580 2972 4586 2984
rect 4816 2972 4844 3012
rect 4890 3000 4896 3052
rect 4948 3040 4954 3052
rect 4948 3012 4993 3040
rect 4948 3000 4954 3012
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 10778 3040 10784 3052
rect 5592 3012 10784 3040
rect 5592 3000 5598 3012
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 5169 2975 5227 2981
rect 5169 2972 5181 2975
rect 4580 2944 4660 2972
rect 4816 2944 5181 2972
rect 4580 2932 4586 2944
rect 1452 2876 2452 2904
rect 1452 2864 1458 2876
rect 2424 2836 2452 2876
rect 2608 2876 3096 2904
rect 3136 2907 3194 2913
rect 2608 2836 2636 2876
rect 3136 2873 3148 2907
rect 3182 2904 3194 2907
rect 3326 2904 3332 2916
rect 3182 2876 3332 2904
rect 3182 2873 3194 2876
rect 3136 2867 3194 2873
rect 3326 2864 3332 2876
rect 3384 2864 3390 2916
rect 4632 2904 4660 2944
rect 5169 2941 5181 2944
rect 5215 2941 5227 2975
rect 5169 2935 5227 2941
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 5902 2972 5908 2984
rect 5767 2944 5908 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2972 6883 2975
rect 6914 2972 6920 2984
rect 6871 2944 6920 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 6914 2932 6920 2944
rect 6972 2972 6978 2984
rect 7282 2972 7288 2984
rect 6972 2944 7288 2972
rect 6972 2932 6978 2944
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7929 2975 7987 2981
rect 7929 2941 7941 2975
rect 7975 2972 7987 2975
rect 8202 2972 8208 2984
rect 7975 2944 8208 2972
rect 7975 2941 7987 2944
rect 7929 2935 7987 2941
rect 4801 2907 4859 2913
rect 4801 2904 4813 2907
rect 4632 2876 4813 2904
rect 4801 2873 4813 2876
rect 4847 2873 4859 2907
rect 5442 2904 5448 2916
rect 5403 2876 5448 2904
rect 4801 2867 4859 2873
rect 5442 2864 5448 2876
rect 5500 2864 5506 2916
rect 5994 2864 6000 2916
rect 6052 2904 6058 2916
rect 7944 2904 7972 2935
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 9033 2975 9091 2981
rect 9033 2941 9045 2975
rect 9079 2972 9091 2975
rect 9398 2972 9404 2984
rect 9079 2944 9404 2972
rect 9079 2941 9091 2944
rect 9033 2935 9091 2941
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 9490 2932 9496 2984
rect 9548 2972 9554 2984
rect 10137 2975 10195 2981
rect 10137 2972 10149 2975
rect 9548 2944 10149 2972
rect 9548 2932 9554 2944
rect 10137 2941 10149 2944
rect 10183 2941 10195 2975
rect 10137 2935 10195 2941
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11330 2972 11336 2984
rect 11287 2944 11336 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 13262 2932 13268 2984
rect 13320 2972 13326 2984
rect 13357 2975 13415 2981
rect 13357 2972 13369 2975
rect 13320 2944 13369 2972
rect 13320 2932 13326 2944
rect 13357 2941 13369 2944
rect 13403 2941 13415 2975
rect 13357 2935 13415 2941
rect 6052 2876 7972 2904
rect 6052 2864 6058 2876
rect 8478 2864 8484 2916
rect 8536 2904 8542 2916
rect 11790 2904 11796 2916
rect 8536 2876 11796 2904
rect 8536 2864 8542 2876
rect 11790 2864 11796 2876
rect 11848 2864 11854 2916
rect 2424 2808 2636 2836
rect 2777 2839 2835 2845
rect 2777 2805 2789 2839
rect 2823 2836 2835 2839
rect 4154 2836 4160 2848
rect 2823 2808 4160 2836
rect 2823 2805 2835 2808
rect 2777 2799 2835 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 4249 2839 4307 2845
rect 4249 2805 4261 2839
rect 4295 2836 4307 2839
rect 4614 2836 4620 2848
rect 4295 2808 4620 2836
rect 4295 2805 4307 2808
rect 4249 2799 4307 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 4890 2836 4896 2848
rect 4755 2808 4896 2836
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 4890 2796 4896 2808
rect 4948 2796 4954 2848
rect 5902 2836 5908 2848
rect 5863 2808 5908 2836
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 7009 2839 7067 2845
rect 7009 2836 7021 2839
rect 6420 2808 7021 2836
rect 6420 2796 6426 2808
rect 7009 2805 7021 2808
rect 7055 2805 7067 2839
rect 7009 2799 7067 2805
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 8113 2839 8171 2845
rect 8113 2836 8125 2839
rect 7524 2808 8125 2836
rect 7524 2796 7530 2808
rect 8113 2805 8125 2808
rect 8159 2805 8171 2839
rect 8113 2799 8171 2805
rect 8202 2796 8208 2848
rect 8260 2836 8266 2848
rect 9674 2836 9680 2848
rect 8260 2808 9680 2836
rect 8260 2796 8266 2808
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 11054 2836 11060 2848
rect 10367 2808 11060 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 1104 2746 14812 2768
rect 1104 2694 5579 2746
rect 5631 2694 5643 2746
rect 5695 2694 5707 2746
rect 5759 2694 5771 2746
rect 5823 2694 10176 2746
rect 10228 2694 10240 2746
rect 10292 2694 10304 2746
rect 10356 2694 10368 2746
rect 10420 2694 14812 2746
rect 1104 2672 14812 2694
rect 5994 2632 6000 2644
rect 1872 2604 6000 2632
rect 1664 2567 1722 2573
rect 1664 2533 1676 2567
rect 1710 2564 1722 2567
rect 1872 2564 1900 2604
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 13538 2632 13544 2644
rect 13499 2604 13544 2632
rect 13538 2592 13544 2604
rect 13596 2592 13602 2644
rect 1710 2536 1900 2564
rect 1710 2533 1722 2536
rect 1664 2527 1722 2533
rect 1946 2524 1952 2576
rect 2004 2564 2010 2576
rect 4341 2567 4399 2573
rect 4341 2564 4353 2567
rect 2004 2536 4353 2564
rect 2004 2524 2010 2536
rect 4341 2533 4353 2536
rect 4387 2533 4399 2567
rect 5626 2564 5632 2576
rect 4341 2527 4399 2533
rect 4448 2536 5632 2564
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 2866 2496 2872 2508
rect 1443 2468 2872 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 4062 2496 4068 2508
rect 3283 2468 3924 2496
rect 4023 2468 4068 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 3694 2428 3700 2440
rect 3559 2400 3700 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 2406 2320 2412 2372
rect 2464 2360 2470 2372
rect 2777 2363 2835 2369
rect 2777 2360 2789 2363
rect 2464 2332 2789 2360
rect 2464 2320 2470 2332
rect 2777 2329 2789 2332
rect 2823 2360 2835 2363
rect 3050 2360 3056 2372
rect 2823 2332 3056 2360
rect 2823 2329 2835 2332
rect 2777 2323 2835 2329
rect 3050 2320 3056 2332
rect 3108 2320 3114 2372
rect 3344 2360 3372 2391
rect 3694 2388 3700 2400
rect 3752 2388 3758 2440
rect 3896 2428 3924 2468
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4448 2428 4476 2536
rect 5626 2524 5632 2536
rect 5684 2524 5690 2576
rect 7184 2567 7242 2573
rect 6012 2536 6500 2564
rect 4522 2456 4528 2508
rect 4580 2496 4586 2508
rect 4873 2499 4931 2505
rect 4873 2496 4885 2499
rect 4580 2468 4885 2496
rect 4580 2456 4586 2468
rect 4873 2465 4885 2468
rect 4919 2496 4931 2499
rect 6012 2496 6040 2536
rect 4919 2468 6040 2496
rect 6089 2499 6147 2505
rect 4919 2465 4931 2468
rect 4873 2459 4931 2465
rect 6089 2465 6101 2499
rect 6135 2496 6147 2499
rect 6178 2496 6184 2508
rect 6135 2468 6184 2496
rect 6135 2465 6147 2468
rect 6089 2459 6147 2465
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 6472 2505 6500 2536
rect 7184 2533 7196 2567
rect 7230 2564 7242 2567
rect 7282 2564 7288 2576
rect 7230 2536 7288 2564
rect 7230 2533 7242 2536
rect 7184 2527 7242 2533
rect 7282 2524 7288 2536
rect 7340 2524 7346 2576
rect 6457 2499 6515 2505
rect 6457 2465 6469 2499
rect 6503 2465 6515 2499
rect 6457 2459 6515 2465
rect 6822 2456 6828 2508
rect 6880 2496 6886 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6880 2468 6929 2496
rect 6880 2456 6886 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 8312 2496 8340 2592
rect 9950 2524 9956 2576
rect 10008 2564 10014 2576
rect 15194 2564 15200 2576
rect 10008 2536 15200 2564
rect 10008 2524 10014 2536
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 8312 2468 9781 2496
rect 6917 2459 6975 2465
rect 9769 2465 9781 2468
rect 9815 2465 9827 2499
rect 9769 2459 9827 2465
rect 10226 2456 10232 2508
rect 10284 2496 10290 2508
rect 10870 2496 10876 2508
rect 10284 2468 10876 2496
rect 10284 2456 10290 2468
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 12250 2496 12256 2508
rect 11471 2468 12256 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 12250 2456 12256 2468
rect 12308 2456 12314 2508
rect 13354 2496 13360 2508
rect 13315 2468 13360 2496
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 4614 2428 4620 2440
rect 3896 2400 4476 2428
rect 4575 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 6638 2428 6644 2440
rect 5684 2400 6644 2428
rect 5684 2388 5690 2400
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 3602 2360 3608 2372
rect 3344 2332 3608 2360
rect 3602 2320 3608 2332
rect 3660 2320 3666 2372
rect 5997 2363 6055 2369
rect 5997 2329 6009 2363
rect 6043 2360 6055 2363
rect 6546 2360 6552 2372
rect 6043 2332 6552 2360
rect 6043 2329 6055 2332
rect 5997 2323 6055 2329
rect 2866 2252 2872 2304
rect 2924 2292 2930 2304
rect 2924 2264 2969 2292
rect 2924 2252 2930 2264
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 6012 2292 6040 2323
rect 6546 2320 6552 2332
rect 6604 2320 6610 2372
rect 6270 2292 6276 2304
rect 4212 2264 6040 2292
rect 6231 2264 6276 2292
rect 4212 2252 4218 2264
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 6641 2295 6699 2301
rect 6641 2261 6653 2295
rect 6687 2292 6699 2295
rect 8570 2292 8576 2304
rect 6687 2264 8576 2292
rect 6687 2261 6699 2264
rect 6641 2255 6699 2261
rect 8570 2252 8576 2264
rect 8628 2252 8634 2304
rect 9950 2292 9956 2304
rect 9911 2264 9956 2292
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 1104 2202 14812 2224
rect 1104 2150 3280 2202
rect 3332 2150 3344 2202
rect 3396 2150 3408 2202
rect 3460 2150 3472 2202
rect 3524 2150 7878 2202
rect 7930 2150 7942 2202
rect 7994 2150 8006 2202
rect 8058 2150 8070 2202
rect 8122 2150 12475 2202
rect 12527 2150 12539 2202
rect 12591 2150 12603 2202
rect 12655 2150 12667 2202
rect 12719 2150 14812 2202
rect 1104 2128 14812 2150
rect 3602 2048 3608 2100
rect 3660 2088 3666 2100
rect 7098 2088 7104 2100
rect 3660 2060 7104 2088
rect 3660 2048 3666 2060
rect 7098 2048 7104 2060
rect 7156 2048 7162 2100
rect 6270 1980 6276 2032
rect 6328 2020 6334 2032
rect 10962 2020 10968 2032
rect 6328 1992 10968 2020
rect 6328 1980 6334 1992
rect 10962 1980 10968 1992
rect 11020 1980 11026 2032
rect 4062 1912 4068 1964
rect 4120 1952 4126 1964
rect 11698 1952 11704 1964
rect 4120 1924 11704 1952
rect 4120 1912 4126 1924
rect 11698 1912 11704 1924
rect 11756 1912 11762 1964
rect 3050 1844 3056 1896
rect 3108 1884 3114 1896
rect 7374 1884 7380 1896
rect 3108 1856 7380 1884
rect 3108 1844 3114 1856
rect 7374 1844 7380 1856
rect 7432 1844 7438 1896
rect 2866 1776 2872 1828
rect 2924 1816 2930 1828
rect 8846 1816 8852 1828
rect 2924 1788 8852 1816
rect 2924 1776 2930 1788
rect 8846 1776 8852 1788
rect 8904 1776 8910 1828
rect 12986 1640 12992 1692
rect 13044 1680 13050 1692
rect 13446 1680 13452 1692
rect 13044 1652 13452 1680
rect 13044 1640 13050 1652
rect 13446 1640 13452 1652
rect 13504 1640 13510 1692
rect 3050 1436 3056 1488
rect 3108 1476 3114 1488
rect 5442 1476 5448 1488
rect 3108 1448 5448 1476
rect 3108 1436 3114 1448
rect 5442 1436 5448 1448
rect 5500 1436 5506 1488
rect 6914 1368 6920 1420
rect 6972 1408 6978 1420
rect 9950 1408 9956 1420
rect 6972 1380 9956 1408
rect 6972 1368 6978 1380
rect 9950 1368 9956 1380
rect 10008 1368 10014 1420
rect 9582 1300 9588 1352
rect 9640 1340 9646 1352
rect 12618 1340 12624 1352
rect 9640 1312 12624 1340
rect 9640 1300 9646 1312
rect 12618 1300 12624 1312
rect 12676 1300 12682 1352
rect 2682 960 2688 1012
rect 2740 1000 2746 1012
rect 3602 1000 3608 1012
rect 2740 972 3608 1000
rect 2740 960 2746 972
rect 3602 960 3608 972
rect 3660 960 3666 1012
rect 2774 756 2780 808
rect 2832 796 2838 808
rect 5166 796 5172 808
rect 2832 768 5172 796
rect 2832 756 2838 768
rect 5166 756 5172 768
rect 5224 756 5230 808
rect 2866 688 2872 740
rect 2924 728 2930 740
rect 5902 728 5908 740
rect 2924 700 5908 728
rect 2924 688 2930 700
rect 5902 688 5908 700
rect 5960 688 5966 740
<< via1 >>
rect 3332 15036 3384 15088
rect 6828 15036 6880 15088
rect 2780 14220 2832 14272
rect 7288 14220 7340 14272
rect 4068 14152 4120 14204
rect 6920 14152 6972 14204
rect 4344 14016 4396 14068
rect 8484 14016 8536 14068
rect 5080 13948 5132 14000
rect 11244 13948 11296 14000
rect 5264 13880 5316 13932
rect 11060 13880 11112 13932
rect 4068 13812 4120 13864
rect 5448 13812 5500 13864
rect 4804 13744 4856 13796
rect 7748 13812 7800 13864
rect 11152 13812 11204 13864
rect 1952 13676 2004 13728
rect 6184 13676 6236 13728
rect 5579 13574 5631 13626
rect 5643 13574 5695 13626
rect 5707 13574 5759 13626
rect 5771 13574 5823 13626
rect 10176 13574 10228 13626
rect 10240 13574 10292 13626
rect 10304 13574 10356 13626
rect 10368 13574 10420 13626
rect 1124 13472 1176 13524
rect 11520 13515 11572 13524
rect 11520 13481 11529 13515
rect 11529 13481 11563 13515
rect 11563 13481 11572 13515
rect 11520 13472 11572 13481
rect 3056 13404 3108 13456
rect 8208 13404 8260 13456
rect 4804 13336 4856 13388
rect 4896 13336 4948 13388
rect 5264 13336 5316 13388
rect 7104 13336 7156 13388
rect 10600 13404 10652 13456
rect 9128 13336 9180 13388
rect 10508 13336 10560 13388
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 9220 13268 9272 13320
rect 1676 13132 1728 13184
rect 4160 13132 4212 13184
rect 5356 13175 5408 13184
rect 5356 13141 5365 13175
rect 5365 13141 5399 13175
rect 5399 13141 5408 13175
rect 5356 13132 5408 13141
rect 8852 13200 8904 13252
rect 10048 13200 10100 13252
rect 7380 13132 7432 13184
rect 9312 13132 9364 13184
rect 9772 13175 9824 13184
rect 9772 13141 9781 13175
rect 9781 13141 9815 13175
rect 9815 13141 9824 13175
rect 9772 13132 9824 13141
rect 3280 13030 3332 13082
rect 3344 13030 3396 13082
rect 3408 13030 3460 13082
rect 3472 13030 3524 13082
rect 7878 13030 7930 13082
rect 7942 13030 7994 13082
rect 8006 13030 8058 13082
rect 8070 13030 8122 13082
rect 12475 13030 12527 13082
rect 12539 13030 12591 13082
rect 12603 13030 12655 13082
rect 12667 13030 12719 13082
rect 2044 12928 2096 12980
rect 5172 12928 5224 12980
rect 13544 12928 13596 12980
rect 2504 12860 2556 12912
rect 2136 12767 2188 12776
rect 2136 12733 2145 12767
rect 2145 12733 2179 12767
rect 2179 12733 2188 12767
rect 2136 12724 2188 12733
rect 3240 12767 3292 12776
rect 3240 12733 3249 12767
rect 3249 12733 3283 12767
rect 3283 12733 3292 12767
rect 3240 12724 3292 12733
rect 3700 12724 3752 12776
rect 7288 12860 7340 12912
rect 6092 12792 6144 12844
rect 11060 12792 11112 12844
rect 2872 12588 2924 12640
rect 3516 12588 3568 12640
rect 4436 12588 4488 12640
rect 5080 12588 5132 12640
rect 7012 12724 7064 12776
rect 7656 12724 7708 12776
rect 9680 12724 9732 12776
rect 9864 12656 9916 12708
rect 6000 12588 6052 12640
rect 9772 12588 9824 12640
rect 11336 12724 11388 12776
rect 13084 12724 13136 12776
rect 11152 12656 11204 12708
rect 10968 12588 11020 12640
rect 5579 12486 5631 12538
rect 5643 12486 5695 12538
rect 5707 12486 5759 12538
rect 5771 12486 5823 12538
rect 10176 12486 10228 12538
rect 10240 12486 10292 12538
rect 10304 12486 10356 12538
rect 10368 12486 10420 12538
rect 3240 12384 3292 12436
rect 6644 12384 6696 12436
rect 7104 12384 7156 12436
rect 8484 12384 8536 12436
rect 9772 12384 9824 12436
rect 4988 12316 5040 12368
rect 7012 12316 7064 12368
rect 7196 12316 7248 12368
rect 8392 12316 8444 12368
rect 2688 12248 2740 12300
rect 4252 12248 4304 12300
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 9036 12248 9088 12300
rect 10692 12316 10744 12368
rect 11428 12316 11480 12368
rect 11796 12316 11848 12368
rect 11980 12316 12032 12368
rect 14740 12384 14792 12436
rect 14096 12316 14148 12368
rect 388 12180 440 12232
rect 7104 12180 7156 12232
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 11336 12248 11388 12300
rect 2044 12044 2096 12096
rect 2412 12044 2464 12096
rect 4804 12044 4856 12096
rect 6736 12044 6788 12096
rect 11980 12180 12032 12232
rect 8944 12112 8996 12164
rect 9680 12112 9732 12164
rect 13912 12112 13964 12164
rect 9036 12044 9088 12096
rect 10508 12044 10560 12096
rect 13452 12044 13504 12096
rect 3280 11942 3332 11994
rect 3344 11942 3396 11994
rect 3408 11942 3460 11994
rect 3472 11942 3524 11994
rect 7878 11942 7930 11994
rect 7942 11942 7994 11994
rect 8006 11942 8058 11994
rect 8070 11942 8122 11994
rect 12475 11942 12527 11994
rect 12539 11942 12591 11994
rect 12603 11942 12655 11994
rect 12667 11942 12719 11994
rect 3608 11840 3660 11892
rect 4528 11840 4580 11892
rect 5908 11883 5960 11892
rect 5908 11849 5917 11883
rect 5917 11849 5951 11883
rect 5951 11849 5960 11883
rect 5908 11840 5960 11849
rect 7196 11840 7248 11892
rect 7472 11840 7524 11892
rect 9220 11840 9272 11892
rect 9864 11840 9916 11892
rect 12256 11840 12308 11892
rect 1952 11772 2004 11824
rect 2780 11636 2832 11688
rect 3516 11772 3568 11824
rect 4252 11772 4304 11824
rect 6184 11772 6236 11824
rect 9680 11772 9732 11824
rect 9772 11772 9824 11824
rect 10048 11772 10100 11824
rect 12808 11772 12860 11824
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 5080 11704 5132 11756
rect 6552 11704 6604 11756
rect 6644 11704 6696 11756
rect 4068 11568 4120 11620
rect 5908 11636 5960 11688
rect 7012 11636 7064 11688
rect 7564 11704 7616 11756
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 9312 11704 9364 11756
rect 11060 11704 11112 11756
rect 11520 11704 11572 11756
rect 8852 11679 8904 11688
rect 8392 11568 8444 11620
rect 8852 11645 8861 11679
rect 8861 11645 8895 11679
rect 8895 11645 8904 11679
rect 8852 11636 8904 11645
rect 9220 11636 9272 11688
rect 11152 11679 11204 11688
rect 10876 11568 10928 11620
rect 1584 11500 1636 11552
rect 3056 11543 3108 11552
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3056 11500 3108 11509
rect 3792 11500 3844 11552
rect 4344 11500 4396 11552
rect 6644 11500 6696 11552
rect 7472 11500 7524 11552
rect 8944 11500 8996 11552
rect 9404 11500 9456 11552
rect 10784 11500 10836 11552
rect 11152 11645 11161 11679
rect 11161 11645 11195 11679
rect 11195 11645 11204 11679
rect 11152 11636 11204 11645
rect 12900 11679 12952 11688
rect 12900 11645 12909 11679
rect 12909 11645 12943 11679
rect 12943 11645 12952 11679
rect 12900 11636 12952 11645
rect 13544 11568 13596 11620
rect 15568 11568 15620 11620
rect 11612 11500 11664 11552
rect 12900 11500 12952 11552
rect 5579 11398 5631 11450
rect 5643 11398 5695 11450
rect 5707 11398 5759 11450
rect 5771 11398 5823 11450
rect 10176 11398 10228 11450
rect 10240 11398 10292 11450
rect 10304 11398 10356 11450
rect 10368 11398 10420 11450
rect 6460 11296 6512 11348
rect 3056 11228 3108 11280
rect 2136 11160 2188 11212
rect 10140 11228 10192 11280
rect 6828 11160 6880 11212
rect 9220 11160 9272 11212
rect 9772 11160 9824 11212
rect 11060 11160 11112 11212
rect 2228 11092 2280 11144
rect 3148 11092 3200 11144
rect 3608 11092 3660 11144
rect 1400 11024 1452 11076
rect 2412 11024 2464 11076
rect 3884 11024 3936 11076
rect 4252 11024 4304 11076
rect 7656 11092 7708 11144
rect 8484 11135 8536 11144
rect 6368 11024 6420 11076
rect 6736 11024 6788 11076
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 8944 11024 8996 11076
rect 3976 10956 4028 11008
rect 9312 10956 9364 11008
rect 10692 11092 10744 11144
rect 12072 11024 12124 11076
rect 12348 11024 12400 11076
rect 10968 10956 11020 11008
rect 3280 10854 3332 10906
rect 3344 10854 3396 10906
rect 3408 10854 3460 10906
rect 3472 10854 3524 10906
rect 7878 10854 7930 10906
rect 7942 10854 7994 10906
rect 8006 10854 8058 10906
rect 8070 10854 8122 10906
rect 12475 10854 12527 10906
rect 12539 10854 12591 10906
rect 12603 10854 12655 10906
rect 12667 10854 12719 10906
rect 9128 10752 9180 10804
rect 2504 10548 2556 10600
rect 3148 10591 3200 10600
rect 3148 10557 3182 10591
rect 3182 10557 3200 10591
rect 3148 10548 3200 10557
rect 2964 10480 3016 10532
rect 5816 10684 5868 10736
rect 6000 10684 6052 10736
rect 9496 10684 9548 10736
rect 6184 10616 6236 10668
rect 7564 10616 7616 10668
rect 8024 10616 8076 10668
rect 8576 10616 8628 10668
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 6092 10480 6144 10532
rect 8392 10548 8444 10600
rect 11060 10616 11112 10668
rect 13544 10684 13596 10736
rect 11704 10616 11756 10668
rect 12072 10616 12124 10668
rect 9312 10548 9364 10600
rect 11152 10548 11204 10600
rect 2320 10412 2372 10464
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 4252 10412 4304 10421
rect 5264 10455 5316 10464
rect 5264 10421 5273 10455
rect 5273 10421 5307 10455
rect 5307 10421 5316 10455
rect 5264 10412 5316 10421
rect 7104 10412 7156 10464
rect 7564 10412 7616 10464
rect 8760 10412 8812 10464
rect 9680 10412 9732 10464
rect 11704 10480 11756 10532
rect 11612 10412 11664 10464
rect 13176 10455 13228 10464
rect 13176 10421 13185 10455
rect 13185 10421 13219 10455
rect 13219 10421 13228 10455
rect 13176 10412 13228 10421
rect 5579 10310 5631 10362
rect 5643 10310 5695 10362
rect 5707 10310 5759 10362
rect 5771 10310 5823 10362
rect 10176 10310 10228 10362
rect 10240 10310 10292 10362
rect 10304 10310 10356 10362
rect 10368 10310 10420 10362
rect 2504 10208 2556 10260
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 2504 10072 2556 10124
rect 2688 10140 2740 10192
rect 4252 10140 4304 10192
rect 4620 10004 4672 10056
rect 3976 9936 4028 9988
rect 4252 9936 4304 9988
rect 5816 9936 5868 9988
rect 2412 9868 2464 9920
rect 6000 9868 6052 9920
rect 7196 10208 7248 10260
rect 7472 10208 7524 10260
rect 8576 10251 8628 10260
rect 8576 10217 8585 10251
rect 8585 10217 8619 10251
rect 8619 10217 8628 10251
rect 8576 10208 8628 10217
rect 9036 10208 9088 10260
rect 9128 10208 9180 10260
rect 12256 10208 12308 10260
rect 7012 10140 7064 10192
rect 7472 10115 7524 10124
rect 7472 10081 7506 10115
rect 7506 10081 7524 10115
rect 7472 10072 7524 10081
rect 8024 10072 8076 10124
rect 8208 10072 8260 10124
rect 9312 10072 9364 10124
rect 10048 10140 10100 10192
rect 7196 10047 7248 10056
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 10968 10072 11020 10124
rect 11612 10072 11664 10124
rect 11704 10072 11756 10124
rect 12164 9936 12216 9988
rect 10600 9868 10652 9920
rect 12992 9868 13044 9920
rect 3280 9766 3332 9818
rect 3344 9766 3396 9818
rect 3408 9766 3460 9818
rect 3472 9766 3524 9818
rect 7878 9766 7930 9818
rect 7942 9766 7994 9818
rect 8006 9766 8058 9818
rect 8070 9766 8122 9818
rect 12475 9766 12527 9818
rect 12539 9766 12591 9818
rect 12603 9766 12655 9818
rect 12667 9766 12719 9818
rect 1492 9664 1544 9716
rect 2872 9664 2924 9716
rect 4252 9664 4304 9716
rect 2228 9639 2280 9648
rect 2228 9605 2237 9639
rect 2237 9605 2271 9639
rect 2271 9605 2280 9639
rect 2228 9596 2280 9605
rect 5816 9664 5868 9716
rect 6184 9664 6236 9716
rect 6276 9596 6328 9648
rect 2504 9528 2556 9580
rect 5080 9528 5132 9580
rect 7380 9596 7432 9648
rect 7196 9528 7248 9580
rect 9772 9596 9824 9648
rect 10048 9528 10100 9580
rect 11152 9664 11204 9716
rect 13084 9664 13136 9716
rect 13360 9664 13412 9716
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 1032 9460 1084 9512
rect 1676 9460 1728 9512
rect 2596 9503 2648 9512
rect 2596 9469 2605 9503
rect 2605 9469 2639 9503
rect 2639 9469 2648 9503
rect 2596 9460 2648 9469
rect 3608 9460 3660 9512
rect 3976 9460 4028 9512
rect 4620 9460 4672 9512
rect 5172 9460 5224 9512
rect 5448 9460 5500 9512
rect 7012 9460 7064 9512
rect 7564 9460 7616 9512
rect 8576 9460 8628 9512
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 3332 9392 3384 9444
rect 4160 9435 4212 9444
rect 4160 9401 4172 9435
rect 4172 9401 4212 9435
rect 4160 9392 4212 9401
rect 1676 9324 1728 9376
rect 4620 9324 4672 9376
rect 7288 9324 7340 9376
rect 12072 9392 12124 9444
rect 11612 9324 11664 9376
rect 12716 9324 12768 9376
rect 5579 9222 5631 9274
rect 5643 9222 5695 9274
rect 5707 9222 5759 9274
rect 5771 9222 5823 9274
rect 10176 9222 10228 9274
rect 10240 9222 10292 9274
rect 10304 9222 10356 9274
rect 10368 9222 10420 9274
rect 2688 9120 2740 9172
rect 4068 9163 4120 9172
rect 4068 9129 4077 9163
rect 4077 9129 4111 9163
rect 4111 9129 4120 9163
rect 4068 9120 4120 9129
rect 7012 9120 7064 9172
rect 7748 9120 7800 9172
rect 8576 9120 8628 9172
rect 11060 9120 11112 9172
rect 12716 9163 12768 9172
rect 12716 9129 12725 9163
rect 12725 9129 12759 9163
rect 12759 9129 12768 9163
rect 12716 9120 12768 9129
rect 13268 9120 13320 9172
rect 13820 9120 13872 9172
rect 4160 9052 4212 9104
rect 5448 9052 5500 9104
rect 5816 9052 5868 9104
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 4436 9027 4488 9036
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 6276 8984 6328 9036
rect 2504 8916 2556 8968
rect 3332 8916 3384 8968
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 5816 8916 5868 8968
rect 7012 8984 7064 9036
rect 8208 8984 8260 9036
rect 10048 8984 10100 9036
rect 12992 9052 13044 9104
rect 13268 8984 13320 9036
rect 848 8848 900 8900
rect 5908 8848 5960 8900
rect 7656 8916 7708 8968
rect 12808 8959 12860 8968
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 8300 8848 8352 8900
rect 9220 8848 9272 8900
rect 11520 8891 11572 8900
rect 4068 8780 4120 8832
rect 8484 8780 8536 8832
rect 9772 8780 9824 8832
rect 11520 8857 11529 8891
rect 11529 8857 11563 8891
rect 11563 8857 11572 8891
rect 11520 8848 11572 8857
rect 10784 8780 10836 8832
rect 11704 8780 11756 8832
rect 3280 8678 3332 8730
rect 3344 8678 3396 8730
rect 3408 8678 3460 8730
rect 3472 8678 3524 8730
rect 7878 8678 7930 8730
rect 7942 8678 7994 8730
rect 8006 8678 8058 8730
rect 8070 8678 8122 8730
rect 12475 8678 12527 8730
rect 12539 8678 12591 8730
rect 12603 8678 12655 8730
rect 12667 8678 12719 8730
rect 2136 8619 2188 8628
rect 2136 8585 2145 8619
rect 2145 8585 2179 8619
rect 2179 8585 2188 8619
rect 2136 8576 2188 8585
rect 3792 8619 3844 8628
rect 1400 8508 1452 8560
rect 2596 8508 2648 8560
rect 3792 8585 3801 8619
rect 3801 8585 3835 8619
rect 3835 8585 3844 8619
rect 3792 8576 3844 8585
rect 10416 8576 10468 8628
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 10784 8576 10836 8585
rect 12808 8576 12860 8628
rect 3976 8508 4028 8560
rect 4620 8440 4672 8492
rect 2504 8415 2556 8424
rect 2504 8381 2513 8415
rect 2513 8381 2547 8415
rect 2547 8381 2556 8415
rect 2504 8372 2556 8381
rect 4896 8372 4948 8424
rect 5908 8440 5960 8492
rect 9036 8508 9088 8560
rect 6828 8372 6880 8424
rect 6920 8372 6972 8424
rect 7656 8440 7708 8492
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 9128 8440 9180 8492
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 2228 8304 2280 8356
rect 4068 8236 4120 8288
rect 4620 8236 4672 8288
rect 7380 8236 7432 8288
rect 8484 8304 8536 8356
rect 9036 8304 9088 8356
rect 9772 8372 9824 8424
rect 10416 8372 10468 8424
rect 11152 8347 11204 8356
rect 10048 8236 10100 8288
rect 11152 8313 11161 8347
rect 11161 8313 11195 8347
rect 11195 8313 11204 8347
rect 11152 8304 11204 8313
rect 12716 8304 12768 8356
rect 11060 8236 11112 8288
rect 5579 8134 5631 8186
rect 5643 8134 5695 8186
rect 5707 8134 5759 8186
rect 5771 8134 5823 8186
rect 10176 8134 10228 8186
rect 10240 8134 10292 8186
rect 10304 8134 10356 8186
rect 10368 8134 10420 8186
rect 5448 8075 5500 8084
rect 5448 8041 5457 8075
rect 5457 8041 5491 8075
rect 5491 8041 5500 8075
rect 5448 8032 5500 8041
rect 6552 8032 6604 8084
rect 6828 8032 6880 8084
rect 10048 8032 10100 8084
rect 2872 7964 2924 8016
rect 3608 7964 3660 8016
rect 3976 7964 4028 8016
rect 5264 7964 5316 8016
rect 6920 7964 6972 8016
rect 2136 7828 2188 7880
rect 2412 7828 2464 7880
rect 3792 7896 3844 7948
rect 4896 7896 4948 7948
rect 11520 7964 11572 8016
rect 11796 7896 11848 7948
rect 3608 7828 3660 7880
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 7656 7828 7708 7880
rect 10140 7828 10192 7880
rect 10876 7828 10928 7880
rect 10968 7760 11020 7812
rect 4344 7692 4396 7744
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 10876 7692 10928 7744
rect 12992 7692 13044 7744
rect 13544 7735 13596 7744
rect 13544 7701 13553 7735
rect 13553 7701 13587 7735
rect 13587 7701 13596 7735
rect 13544 7692 13596 7701
rect 3280 7590 3332 7642
rect 3344 7590 3396 7642
rect 3408 7590 3460 7642
rect 3472 7590 3524 7642
rect 7878 7590 7930 7642
rect 7942 7590 7994 7642
rect 8006 7590 8058 7642
rect 8070 7590 8122 7642
rect 12475 7590 12527 7642
rect 12539 7590 12591 7642
rect 12603 7590 12655 7642
rect 12667 7590 12719 7642
rect 3792 7488 3844 7540
rect 4620 7488 4672 7540
rect 7380 7488 7432 7540
rect 10600 7488 10652 7540
rect 11520 7488 11572 7540
rect 12808 7488 12860 7540
rect 4712 7420 4764 7472
rect 5264 7420 5316 7472
rect 7472 7420 7524 7472
rect 11060 7420 11112 7472
rect 2412 7284 2464 7336
rect 2872 7284 2924 7336
rect 4896 7352 4948 7404
rect 5080 7352 5132 7404
rect 5448 7352 5500 7404
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 10784 7352 10836 7404
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 3976 7284 4028 7336
rect 5356 7284 5408 7336
rect 7564 7284 7616 7336
rect 8668 7284 8720 7336
rect 2688 7216 2740 7268
rect 3424 7216 3476 7268
rect 5448 7216 5500 7268
rect 6276 7216 6328 7268
rect 6460 7216 6512 7268
rect 11796 7284 11848 7336
rect 2780 7148 2832 7200
rect 3056 7148 3108 7200
rect 4252 7148 4304 7200
rect 4436 7148 4488 7200
rect 4896 7191 4948 7200
rect 4896 7157 4905 7191
rect 4905 7157 4939 7191
rect 4939 7157 4948 7191
rect 4896 7148 4948 7157
rect 5172 7148 5224 7200
rect 9956 7216 10008 7268
rect 12808 7259 12860 7268
rect 12808 7225 12817 7259
rect 12817 7225 12851 7259
rect 12851 7225 12860 7259
rect 12808 7216 12860 7225
rect 8300 7148 8352 7200
rect 9128 7148 9180 7200
rect 10508 7148 10560 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 5579 7046 5631 7098
rect 5643 7046 5695 7098
rect 5707 7046 5759 7098
rect 5771 7046 5823 7098
rect 10176 7046 10228 7098
rect 10240 7046 10292 7098
rect 10304 7046 10356 7098
rect 10368 7046 10420 7098
rect 2412 6944 2464 6996
rect 4068 6944 4120 6996
rect 4896 6944 4948 6996
rect 11428 6944 11480 6996
rect 13084 6944 13136 6996
rect 4436 6876 4488 6928
rect 2504 6740 2556 6792
rect 3792 6740 3844 6792
rect 7012 6876 7064 6928
rect 8116 6876 8168 6928
rect 12992 6876 13044 6928
rect 6828 6808 6880 6860
rect 7564 6808 7616 6860
rect 9496 6808 9548 6860
rect 9588 6808 9640 6860
rect 10048 6808 10100 6860
rect 10784 6808 10836 6860
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 4712 6672 4764 6724
rect 8208 6672 8260 6724
rect 9312 6740 9364 6792
rect 3056 6604 3108 6656
rect 5080 6604 5132 6656
rect 5908 6604 5960 6656
rect 8484 6647 8536 6656
rect 8484 6613 8493 6647
rect 8493 6613 8527 6647
rect 8527 6613 8536 6647
rect 8484 6604 8536 6613
rect 9496 6604 9548 6656
rect 10968 6672 11020 6724
rect 11336 6715 11388 6724
rect 11336 6681 11345 6715
rect 11345 6681 11379 6715
rect 11379 6681 11388 6715
rect 11336 6672 11388 6681
rect 3280 6502 3332 6554
rect 3344 6502 3396 6554
rect 3408 6502 3460 6554
rect 3472 6502 3524 6554
rect 7878 6502 7930 6554
rect 7942 6502 7994 6554
rect 8006 6502 8058 6554
rect 8070 6502 8122 6554
rect 12475 6502 12527 6554
rect 12539 6502 12591 6554
rect 12603 6502 12655 6554
rect 12667 6502 12719 6554
rect 2688 6400 2740 6452
rect 1308 6332 1360 6384
rect 1952 6332 2004 6384
rect 3424 6332 3476 6384
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 3608 6264 3660 6316
rect 6460 6400 6512 6452
rect 9036 6400 9088 6452
rect 9312 6400 9364 6452
rect 12900 6400 12952 6452
rect 4436 6375 4488 6384
rect 4436 6341 4445 6375
rect 4445 6341 4479 6375
rect 4479 6341 4488 6375
rect 4436 6332 4488 6341
rect 4804 6332 4856 6384
rect 8300 6332 8352 6384
rect 8944 6332 8996 6384
rect 9496 6307 9548 6316
rect 9496 6273 9505 6307
rect 9505 6273 9539 6307
rect 9539 6273 9548 6307
rect 9496 6264 9548 6273
rect 12992 6264 13044 6316
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 4344 6196 4396 6248
rect 9588 6196 9640 6248
rect 3976 6128 4028 6180
rect 3148 6060 3200 6112
rect 4068 6060 4120 6112
rect 4620 6060 4672 6112
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 6000 6060 6052 6112
rect 6276 6060 6328 6112
rect 8208 6128 8260 6180
rect 8300 6128 8352 6180
rect 7656 6060 7708 6112
rect 11060 6128 11112 6180
rect 13636 6128 13688 6180
rect 9956 6060 10008 6112
rect 10876 6060 10928 6112
rect 12900 6060 12952 6112
rect 13360 6060 13412 6112
rect 5579 5958 5631 6010
rect 5643 5958 5695 6010
rect 5707 5958 5759 6010
rect 5771 5958 5823 6010
rect 10176 5958 10228 6010
rect 10240 5958 10292 6010
rect 10304 5958 10356 6010
rect 10368 5958 10420 6010
rect 940 5720 992 5772
rect 8300 5856 8352 5908
rect 9956 5856 10008 5908
rect 11060 5899 11112 5908
rect 11060 5865 11069 5899
rect 11069 5865 11103 5899
rect 11103 5865 11112 5899
rect 11060 5856 11112 5865
rect 12808 5856 12860 5908
rect 4896 5788 4948 5840
rect 6460 5788 6512 5840
rect 7012 5788 7064 5840
rect 9220 5788 9272 5840
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 3424 5720 3476 5772
rect 6736 5720 6788 5772
rect 4160 5652 4212 5704
rect 5264 5652 5316 5704
rect 8300 5652 8352 5704
rect 8576 5652 8628 5704
rect 12256 5788 12308 5840
rect 10968 5720 11020 5772
rect 1952 5627 2004 5636
rect 1952 5593 1961 5627
rect 1961 5593 1995 5627
rect 1995 5593 2004 5627
rect 1952 5584 2004 5593
rect 1676 5516 1728 5568
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 4160 5516 4212 5568
rect 9496 5584 9548 5636
rect 12256 5652 12308 5704
rect 13176 5695 13228 5704
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 6092 5516 6144 5568
rect 6736 5559 6788 5568
rect 6736 5525 6745 5559
rect 6745 5525 6779 5559
rect 6779 5525 6788 5559
rect 6736 5516 6788 5525
rect 8208 5516 8260 5568
rect 8668 5516 8720 5568
rect 11888 5516 11940 5568
rect 3280 5414 3332 5466
rect 3344 5414 3396 5466
rect 3408 5414 3460 5466
rect 3472 5414 3524 5466
rect 7878 5414 7930 5466
rect 7942 5414 7994 5466
rect 8006 5414 8058 5466
rect 8070 5414 8122 5466
rect 12475 5414 12527 5466
rect 12539 5414 12591 5466
rect 12603 5414 12655 5466
rect 12667 5414 12719 5466
rect 1400 5355 1452 5364
rect 1400 5321 1409 5355
rect 1409 5321 1443 5355
rect 1443 5321 1452 5355
rect 1400 5312 1452 5321
rect 4804 5312 4856 5364
rect 4896 5355 4948 5364
rect 4896 5321 4905 5355
rect 4905 5321 4939 5355
rect 4939 5321 4948 5355
rect 4896 5312 4948 5321
rect 5264 5312 5316 5364
rect 6828 5312 6880 5364
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 2228 5176 2280 5228
rect 2504 5176 2556 5228
rect 6736 5244 6788 5296
rect 9496 5312 9548 5364
rect 9956 5355 10008 5364
rect 9956 5321 9965 5355
rect 9965 5321 9999 5355
rect 9999 5321 10008 5355
rect 9956 5312 10008 5321
rect 10324 5312 10376 5364
rect 10508 5312 10560 5364
rect 11060 5244 11112 5296
rect 3516 5176 3568 5228
rect 3700 5176 3752 5228
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 4620 5176 4672 5228
rect 5172 5176 5224 5228
rect 7288 5176 7340 5228
rect 4436 5108 4488 5160
rect 5356 5108 5408 5160
rect 5908 5108 5960 5160
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 3148 5040 3200 5092
rect 4896 5040 4948 5092
rect 7196 5040 7248 5092
rect 7288 5040 7340 5092
rect 1860 4972 1912 4981
rect 2504 4972 2556 5024
rect 4804 4972 4856 5024
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 6460 4972 6512 5024
rect 7748 4972 7800 5024
rect 8300 5040 8352 5092
rect 9220 5176 9272 5228
rect 9588 5176 9640 5228
rect 10232 5176 10284 5228
rect 10968 5176 11020 5228
rect 13176 5219 13228 5228
rect 13176 5185 13185 5219
rect 13185 5185 13219 5219
rect 13219 5185 13228 5219
rect 13176 5176 13228 5185
rect 9772 5151 9824 5160
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 9772 5108 9824 5117
rect 10324 5108 10376 5160
rect 12440 5108 12492 5160
rect 9956 5040 10008 5092
rect 10140 5040 10192 5092
rect 11336 5040 11388 5092
rect 10508 4972 10560 5024
rect 12532 5015 12584 5024
rect 12532 4981 12541 5015
rect 12541 4981 12575 5015
rect 12575 4981 12584 5015
rect 12532 4972 12584 4981
rect 5579 4870 5631 4922
rect 5643 4870 5695 4922
rect 5707 4870 5759 4922
rect 5771 4870 5823 4922
rect 10176 4870 10228 4922
rect 10240 4870 10292 4922
rect 10304 4870 10356 4922
rect 10368 4870 10420 4922
rect 1860 4768 1912 4820
rect 1124 4700 1176 4752
rect 2596 4700 2648 4752
rect 1400 4632 1452 4684
rect 2688 4632 2740 4684
rect 2504 4564 2556 4616
rect 2596 4564 2648 4616
rect 4068 4700 4120 4752
rect 5172 4768 5224 4820
rect 7472 4768 7524 4820
rect 7748 4811 7800 4820
rect 7748 4777 7757 4811
rect 7757 4777 7791 4811
rect 7791 4777 7800 4811
rect 7748 4768 7800 4777
rect 8484 4768 8536 4820
rect 8944 4768 8996 4820
rect 9312 4768 9364 4820
rect 10508 4768 10560 4820
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 11152 4768 11204 4820
rect 12532 4811 12584 4820
rect 12532 4777 12541 4811
rect 12541 4777 12575 4811
rect 12575 4777 12584 4811
rect 12532 4768 12584 4777
rect 5908 4700 5960 4752
rect 6000 4700 6052 4752
rect 3884 4632 3936 4684
rect 5264 4632 5316 4684
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 848 4496 900 4548
rect 3976 4564 4028 4616
rect 5816 4564 5868 4616
rect 10416 4632 10468 4684
rect 7656 4564 7708 4616
rect 9588 4496 9640 4548
rect 4252 4428 4304 4480
rect 7288 4428 7340 4480
rect 10784 4700 10836 4752
rect 11152 4632 11204 4684
rect 12992 4632 13044 4684
rect 13728 4632 13780 4684
rect 11612 4496 11664 4548
rect 11152 4428 11204 4480
rect 3280 4326 3332 4378
rect 3344 4326 3396 4378
rect 3408 4326 3460 4378
rect 3472 4326 3524 4378
rect 7878 4326 7930 4378
rect 7942 4326 7994 4378
rect 8006 4326 8058 4378
rect 8070 4326 8122 4378
rect 12475 4326 12527 4378
rect 12539 4326 12591 4378
rect 12603 4326 12655 4378
rect 12667 4326 12719 4378
rect 1952 4224 2004 4276
rect 1492 4156 1544 4208
rect 2688 4224 2740 4276
rect 1768 4088 1820 4140
rect 2136 4088 2188 4140
rect 4068 4088 4120 4140
rect 7012 4224 7064 4276
rect 5080 4156 5132 4208
rect 6184 4088 6236 4140
rect 2228 4020 2280 4072
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 4344 4020 4396 4072
rect 5080 4020 5132 4072
rect 5264 4020 5316 4072
rect 6920 4020 6972 4072
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 9496 4224 9548 4276
rect 10416 4224 10468 4276
rect 11336 4224 11388 4276
rect 13544 4267 13596 4276
rect 13544 4233 13553 4267
rect 13553 4233 13587 4267
rect 13587 4233 13596 4267
rect 13544 4224 13596 4233
rect 9772 4156 9824 4208
rect 12440 4156 12492 4208
rect 10048 4088 10100 4140
rect 10784 4088 10836 4140
rect 8484 4020 8536 4072
rect 8668 4063 8720 4072
rect 8668 4029 8702 4063
rect 8702 4029 8720 4063
rect 8668 4020 8720 4029
rect 9036 4020 9088 4072
rect 11152 4020 11204 4072
rect 1952 3952 2004 4004
rect 8944 3952 8996 4004
rect 11796 3952 11848 4004
rect 1400 3927 1452 3936
rect 1400 3893 1409 3927
rect 1409 3893 1443 3927
rect 1443 3893 1452 3927
rect 1400 3884 1452 3893
rect 2136 3884 2188 3936
rect 2596 3927 2648 3936
rect 2596 3893 2605 3927
rect 2605 3893 2639 3927
rect 2639 3893 2648 3927
rect 2596 3884 2648 3893
rect 2688 3884 2740 3936
rect 3056 3884 3108 3936
rect 3700 3927 3752 3936
rect 3700 3893 3709 3927
rect 3709 3893 3743 3927
rect 3743 3893 3752 3927
rect 3700 3884 3752 3893
rect 3792 3884 3844 3936
rect 4344 3884 4396 3936
rect 4528 3884 4580 3936
rect 4804 3884 4856 3936
rect 6920 3884 6972 3936
rect 11428 3927 11480 3936
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 5579 3782 5631 3834
rect 5643 3782 5695 3834
rect 5707 3782 5759 3834
rect 5771 3782 5823 3834
rect 10176 3782 10228 3834
rect 10240 3782 10292 3834
rect 10304 3782 10356 3834
rect 10368 3782 10420 3834
rect 296 3680 348 3732
rect 1952 3680 2004 3732
rect 2596 3680 2648 3732
rect 3056 3680 3108 3732
rect 2688 3612 2740 3664
rect 1952 3544 2004 3596
rect 4068 3680 4120 3732
rect 4804 3680 4856 3732
rect 5448 3723 5500 3732
rect 5448 3689 5457 3723
rect 5457 3689 5491 3723
rect 5491 3689 5500 3723
rect 5448 3680 5500 3689
rect 3700 3612 3752 3664
rect 4528 3655 4580 3664
rect 4528 3621 4537 3655
rect 4537 3621 4571 3655
rect 4571 3621 4580 3655
rect 4528 3612 4580 3621
rect 3976 3544 4028 3596
rect 3884 3476 3936 3528
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 5540 3612 5592 3664
rect 5448 3544 5500 3596
rect 9864 3680 9916 3732
rect 8300 3612 8352 3664
rect 8392 3612 8444 3664
rect 9772 3612 9824 3664
rect 10048 3680 10100 3732
rect 12348 3680 12400 3732
rect 13636 3680 13688 3732
rect 6828 3544 6880 3596
rect 7564 3544 7616 3596
rect 6368 3476 6420 3528
rect 8208 3544 8260 3596
rect 10048 3544 10100 3596
rect 12440 3544 12492 3596
rect 2872 3408 2924 3460
rect 3608 3340 3660 3392
rect 6276 3408 6328 3460
rect 4252 3340 4304 3392
rect 4528 3340 4580 3392
rect 4620 3340 4672 3392
rect 4896 3340 4948 3392
rect 5080 3383 5132 3392
rect 5080 3349 5089 3383
rect 5089 3349 5123 3383
rect 5123 3349 5132 3383
rect 5080 3340 5132 3349
rect 9680 3408 9732 3460
rect 8208 3340 8260 3392
rect 9864 3340 9916 3392
rect 10600 3340 10652 3392
rect 11520 3340 11572 3392
rect 3280 3238 3332 3290
rect 3344 3238 3396 3290
rect 3408 3238 3460 3290
rect 3472 3238 3524 3290
rect 7878 3238 7930 3290
rect 7942 3238 7994 3290
rect 8006 3238 8058 3290
rect 8070 3238 8122 3290
rect 12475 3238 12527 3290
rect 12539 3238 12591 3290
rect 12603 3238 12655 3290
rect 12667 3238 12719 3290
rect 2504 3136 2556 3188
rect 10140 3136 10192 3188
rect 13728 3136 13780 3188
rect 5356 3068 5408 3120
rect 15752 3068 15804 3120
rect 4436 3000 4488 3052
rect 2412 2932 2464 2984
rect 2872 2975 2924 2984
rect 2872 2941 2881 2975
rect 2881 2941 2915 2975
rect 2915 2941 2924 2975
rect 2872 2932 2924 2941
rect 1400 2864 1452 2916
rect 4344 2932 4396 2984
rect 4528 2932 4580 2984
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 5540 3000 5592 3052
rect 10784 3000 10836 3052
rect 3332 2864 3384 2916
rect 5908 2932 5960 2984
rect 6920 2932 6972 2984
rect 7288 2932 7340 2984
rect 5448 2907 5500 2916
rect 5448 2873 5457 2907
rect 5457 2873 5491 2907
rect 5491 2873 5500 2907
rect 5448 2864 5500 2873
rect 6000 2864 6052 2916
rect 8208 2932 8260 2984
rect 9404 2932 9456 2984
rect 9496 2932 9548 2984
rect 11336 2932 11388 2984
rect 13268 2932 13320 2984
rect 8484 2864 8536 2916
rect 11796 2864 11848 2916
rect 4160 2796 4212 2848
rect 4620 2796 4672 2848
rect 4896 2796 4948 2848
rect 5908 2839 5960 2848
rect 5908 2805 5917 2839
rect 5917 2805 5951 2839
rect 5951 2805 5960 2839
rect 5908 2796 5960 2805
rect 6368 2796 6420 2848
rect 7472 2796 7524 2848
rect 8208 2796 8260 2848
rect 9680 2796 9732 2848
rect 11060 2796 11112 2848
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 5579 2694 5631 2746
rect 5643 2694 5695 2746
rect 5707 2694 5759 2746
rect 5771 2694 5823 2746
rect 10176 2694 10228 2746
rect 10240 2694 10292 2746
rect 10304 2694 10356 2746
rect 10368 2694 10420 2746
rect 6000 2592 6052 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 13544 2635 13596 2644
rect 13544 2601 13553 2635
rect 13553 2601 13587 2635
rect 13587 2601 13596 2635
rect 13544 2592 13596 2601
rect 1952 2524 2004 2576
rect 2872 2456 2924 2508
rect 4068 2499 4120 2508
rect 2412 2320 2464 2372
rect 3056 2320 3108 2372
rect 3700 2388 3752 2440
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 5632 2524 5684 2576
rect 4528 2456 4580 2508
rect 6184 2456 6236 2508
rect 7288 2524 7340 2576
rect 6828 2456 6880 2508
rect 9956 2524 10008 2576
rect 15200 2524 15252 2576
rect 10232 2456 10284 2508
rect 10876 2456 10928 2508
rect 12256 2456 12308 2508
rect 13360 2499 13412 2508
rect 13360 2465 13369 2499
rect 13369 2465 13403 2499
rect 13403 2465 13412 2499
rect 13360 2456 13412 2465
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5632 2388 5684 2440
rect 6644 2388 6696 2440
rect 3608 2320 3660 2372
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 4160 2252 4212 2304
rect 6552 2320 6604 2372
rect 6276 2295 6328 2304
rect 6276 2261 6285 2295
rect 6285 2261 6319 2295
rect 6319 2261 6328 2295
rect 6276 2252 6328 2261
rect 8576 2252 8628 2304
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 3280 2150 3332 2202
rect 3344 2150 3396 2202
rect 3408 2150 3460 2202
rect 3472 2150 3524 2202
rect 7878 2150 7930 2202
rect 7942 2150 7994 2202
rect 8006 2150 8058 2202
rect 8070 2150 8122 2202
rect 12475 2150 12527 2202
rect 12539 2150 12591 2202
rect 12603 2150 12655 2202
rect 12667 2150 12719 2202
rect 3608 2048 3660 2100
rect 7104 2048 7156 2100
rect 6276 1980 6328 2032
rect 10968 1980 11020 2032
rect 4068 1912 4120 1964
rect 11704 1912 11756 1964
rect 3056 1844 3108 1896
rect 7380 1844 7432 1896
rect 2872 1776 2924 1828
rect 8852 1776 8904 1828
rect 12992 1640 13044 1692
rect 13452 1640 13504 1692
rect 3056 1436 3108 1488
rect 5448 1436 5500 1488
rect 6920 1368 6972 1420
rect 9956 1368 10008 1420
rect 9588 1300 9640 1352
rect 12624 1300 12676 1352
rect 2688 960 2740 1012
rect 3608 960 3660 1012
rect 2780 756 2832 808
rect 5172 756 5224 808
rect 2872 688 2924 740
rect 5908 688 5960 740
<< metal2 >>
rect 386 15520 442 16000
rect 1122 15520 1178 16000
rect 1950 15520 2006 16000
rect 2778 15520 2834 16000
rect 3330 15872 3386 15881
rect 3330 15807 3386 15816
rect 400 12238 428 15520
rect 1136 13530 1164 15520
rect 1490 14648 1546 14657
rect 1490 14583 1546 14592
rect 1124 13524 1176 13530
rect 1124 13466 1176 13472
rect 388 12232 440 12238
rect 388 12174 440 12180
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1032 9512 1084 9518
rect 1032 9454 1084 9460
rect 848 8900 900 8906
rect 848 8842 900 8848
rect 860 6633 888 8842
rect 938 7984 994 7993
rect 938 7919 994 7928
rect 846 6624 902 6633
rect 846 6559 902 6568
rect 952 5778 980 7919
rect 940 5772 992 5778
rect 940 5714 992 5720
rect 848 4548 900 4554
rect 848 4490 900 4496
rect 296 3732 348 3738
rect 296 3674 348 3680
rect 308 480 336 3674
rect 860 480 888 4490
rect 1044 3777 1072 9454
rect 1412 8650 1440 11018
rect 1504 9722 1532 14583
rect 1964 13734 1992 15520
rect 2594 15056 2650 15065
rect 2594 14991 2650 15000
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1492 9716 1544 9722
rect 1492 9658 1544 9664
rect 1228 8622 1440 8650
rect 1122 8256 1178 8265
rect 1122 8191 1178 8200
rect 1136 4758 1164 8191
rect 1124 4752 1176 4758
rect 1124 4694 1176 4700
rect 1228 4593 1256 8622
rect 1400 8560 1452 8566
rect 1400 8502 1452 8508
rect 1308 6384 1360 6390
rect 1308 6326 1360 6332
rect 1320 5250 1348 6326
rect 1412 5370 1440 8502
rect 1490 7304 1546 7313
rect 1490 7239 1546 7248
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1320 5222 1440 5250
rect 1412 4690 1440 5222
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1214 4584 1270 4593
rect 1214 4519 1270 4528
rect 1504 4214 1532 7239
rect 1492 4208 1544 4214
rect 1492 4150 1544 4156
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1030 3768 1086 3777
rect 1030 3703 1086 3712
rect 1412 3097 1440 3878
rect 1398 3088 1454 3097
rect 1398 3023 1454 3032
rect 1400 2916 1452 2922
rect 1400 2858 1452 2864
rect 1412 480 1440 2858
rect 1596 1329 1624 11494
rect 1688 9518 1716 13126
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 2056 12322 2084 12922
rect 2504 12912 2556 12918
rect 2504 12854 2556 12860
rect 2136 12776 2188 12782
rect 2134 12744 2136 12753
rect 2188 12744 2190 12753
rect 2134 12679 2190 12688
rect 1872 12294 2084 12322
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1766 9344 1822 9353
rect 1688 5681 1716 9318
rect 1766 9279 1822 9288
rect 1780 5953 1808 9279
rect 1766 5944 1822 5953
rect 1766 5879 1822 5888
rect 1674 5672 1730 5681
rect 1674 5607 1730 5616
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1688 3641 1716 5510
rect 1780 4536 1808 5879
rect 1872 5409 1900 12294
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 1952 11824 2004 11830
rect 1952 11766 2004 11772
rect 1964 6390 1992 11766
rect 1952 6384 2004 6390
rect 1952 6326 2004 6332
rect 1950 6080 2006 6089
rect 1950 6015 2006 6024
rect 1964 5642 1992 6015
rect 1952 5636 2004 5642
rect 1952 5578 2004 5584
rect 1950 5536 2006 5545
rect 1950 5471 2006 5480
rect 1858 5400 1914 5409
rect 1858 5335 1914 5344
rect 1964 5234 1992 5471
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1872 4826 1900 4966
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1780 4508 1900 4536
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1674 3632 1730 3641
rect 1674 3567 1730 3576
rect 1780 2689 1808 4082
rect 1872 3584 1900 4508
rect 1964 4282 1992 5170
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 1964 3738 1992 3946
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1952 3596 2004 3602
rect 1872 3556 1952 3584
rect 1952 3538 2004 3544
rect 1766 2680 1822 2689
rect 1766 2615 1822 2624
rect 1952 2576 2004 2582
rect 1952 2518 2004 2524
rect 1582 1320 1638 1329
rect 1582 1255 1638 1264
rect 1964 480 1992 2518
rect 2056 1737 2084 12038
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2148 8634 2176 11154
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2240 9654 2268 11086
rect 2424 11082 2452 12038
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2516 10690 2544 12854
rect 2424 10662 2544 10690
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2148 4146 2176 7822
rect 2240 5234 2268 8298
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2226 5128 2282 5137
rect 2226 5063 2282 5072
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2240 4078 2268 5063
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2148 3505 2176 3878
rect 2134 3496 2190 3505
rect 2134 3431 2190 3440
rect 2042 1728 2098 1737
rect 2042 1663 2098 1672
rect 2332 921 2360 10406
rect 2424 10033 2452 10662
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2516 10266 2544 10542
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2608 10180 2636 14991
rect 2792 14278 2820 15520
rect 3344 15094 3372 15807
rect 3514 15520 3570 16000
rect 4342 15520 4398 16000
rect 5170 15520 5226 16000
rect 5906 15520 5962 16000
rect 6734 15520 6790 16000
rect 7562 15520 7618 16000
rect 8390 15520 8446 16000
rect 9126 15520 9182 16000
rect 9954 15520 10010 16000
rect 10782 15520 10838 16000
rect 11518 15520 11574 16000
rect 11610 15872 11666 15881
rect 11610 15807 11666 15816
rect 3332 15088 3384 15094
rect 3332 15030 3384 15036
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 3528 13682 3556 15520
rect 4066 14240 4122 14249
rect 4066 14175 4068 14184
rect 4120 14175 4122 14184
rect 4068 14146 4120 14152
rect 4356 14074 4384 15520
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 5080 14000 5132 14006
rect 5080 13942 5132 13948
rect 4068 13864 4120 13870
rect 4066 13832 4068 13841
rect 4120 13832 4122 13841
rect 4066 13767 4122 13776
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 3528 13654 3648 13682
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 3068 13025 3096 13398
rect 3254 13084 3550 13104
rect 3310 13082 3334 13084
rect 3390 13082 3414 13084
rect 3470 13082 3494 13084
rect 3332 13030 3334 13082
rect 3396 13030 3408 13082
rect 3470 13030 3472 13082
rect 3310 13028 3334 13030
rect 3390 13028 3414 13030
rect 3470 13028 3494 13030
rect 3054 13016 3110 13025
rect 3254 13008 3550 13028
rect 3054 12951 3110 12960
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2700 11121 2728 12242
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2686 11112 2742 11121
rect 2686 11047 2742 11056
rect 2688 10192 2740 10198
rect 2608 10152 2688 10180
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2410 10024 2466 10033
rect 2410 9959 2466 9968
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2424 7886 2452 9862
rect 2516 9586 2544 10066
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2516 9058 2544 9522
rect 2608 9518 2636 10152
rect 2688 10134 2740 10140
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2686 9344 2742 9353
rect 2686 9279 2742 9288
rect 2700 9178 2728 9279
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2792 9081 2820 11630
rect 2884 10112 2912 12582
rect 3252 12481 3280 12718
rect 3516 12640 3568 12646
rect 3514 12608 3516 12617
rect 3568 12608 3570 12617
rect 3514 12543 3570 12552
rect 3238 12472 3294 12481
rect 3238 12407 3240 12416
rect 3292 12407 3294 12416
rect 3240 12378 3292 12384
rect 3252 12347 3280 12378
rect 3254 11996 3550 12016
rect 3310 11994 3334 11996
rect 3390 11994 3414 11996
rect 3470 11994 3494 11996
rect 3332 11942 3334 11994
rect 3396 11942 3408 11994
rect 3470 11942 3472 11994
rect 3310 11940 3334 11942
rect 3390 11940 3414 11942
rect 3470 11940 3494 11942
rect 3254 11920 3550 11940
rect 3620 11898 3648 13654
rect 3882 13424 3938 13433
rect 4816 13394 4844 13738
rect 3882 13359 3938 13368
rect 4804 13388 4856 13394
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3068 11286 3096 11494
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3054 10976 3110 10985
rect 3054 10911 3110 10920
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2976 10305 3004 10474
rect 2962 10296 3018 10305
rect 2962 10231 3018 10240
rect 2884 10084 3004 10112
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2778 9072 2834 9081
rect 2516 9030 2636 9058
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2516 8430 2544 8910
rect 2608 8566 2636 9030
rect 2778 9007 2780 9016
rect 2832 9007 2834 9016
rect 2780 8978 2832 8984
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2792 7392 2820 8978
rect 2884 8022 2912 9658
rect 2872 8016 2924 8022
rect 2872 7958 2924 7964
rect 2608 7364 2820 7392
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2424 7002 2452 7278
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2424 6322 2452 6938
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2516 5658 2544 6734
rect 2424 5630 2544 5658
rect 2424 5574 2452 5630
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2608 5352 2636 7364
rect 2884 7342 2912 7958
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2700 6458 2728 7210
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2792 6338 2820 7142
rect 2424 5324 2636 5352
rect 2700 6310 2820 6338
rect 2424 4026 2452 5324
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2516 5030 2544 5170
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2594 4856 2650 4865
rect 2594 4791 2650 4800
rect 2608 4758 2636 4791
rect 2596 4752 2648 4758
rect 2502 4720 2558 4729
rect 2596 4694 2648 4700
rect 2502 4655 2558 4664
rect 2516 4622 2544 4655
rect 2608 4622 2636 4694
rect 2700 4690 2728 6310
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2700 4282 2728 4626
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2424 3998 2728 4026
rect 2700 3942 2728 3998
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2608 3738 2636 3878
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2424 2378 2452 2926
rect 2412 2372 2464 2378
rect 2412 2314 2464 2320
rect 2318 912 2374 921
rect 2318 847 2374 856
rect 2516 480 2544 3130
rect 2700 1018 2728 3606
rect 2884 3466 2912 5646
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2884 2514 2912 2926
rect 2976 2553 3004 10084
rect 3068 7206 3096 10911
rect 3160 10606 3188 11086
rect 3528 10996 3556 11766
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3620 11150 3648 11698
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3528 10968 3648 10996
rect 3254 10908 3550 10928
rect 3310 10906 3334 10908
rect 3390 10906 3414 10908
rect 3470 10906 3494 10908
rect 3332 10854 3334 10906
rect 3396 10854 3408 10906
rect 3470 10854 3472 10906
rect 3310 10852 3334 10854
rect 3390 10852 3414 10854
rect 3470 10852 3494 10854
rect 3254 10832 3550 10852
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3160 10266 3188 10542
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3146 10024 3202 10033
rect 3146 9959 3202 9968
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 4078 3096 6598
rect 3160 6202 3188 9959
rect 3254 9820 3550 9840
rect 3310 9818 3334 9820
rect 3390 9818 3414 9820
rect 3470 9818 3494 9820
rect 3332 9766 3334 9818
rect 3396 9766 3408 9818
rect 3470 9766 3472 9818
rect 3310 9764 3334 9766
rect 3390 9764 3414 9766
rect 3470 9764 3494 9766
rect 3254 9744 3550 9764
rect 3620 9518 3648 10968
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3344 8974 3372 9386
rect 3606 9344 3662 9353
rect 3606 9279 3662 9288
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3254 8732 3550 8752
rect 3310 8730 3334 8732
rect 3390 8730 3414 8732
rect 3470 8730 3494 8732
rect 3332 8678 3334 8730
rect 3396 8678 3408 8730
rect 3470 8678 3472 8730
rect 3310 8676 3334 8678
rect 3390 8676 3414 8678
rect 3470 8676 3494 8678
rect 3254 8656 3550 8676
rect 3620 8022 3648 9279
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3254 7644 3550 7664
rect 3310 7642 3334 7644
rect 3390 7642 3414 7644
rect 3470 7642 3494 7644
rect 3332 7590 3334 7642
rect 3396 7590 3408 7642
rect 3470 7590 3472 7642
rect 3310 7588 3334 7590
rect 3390 7588 3414 7590
rect 3470 7588 3494 7590
rect 3254 7568 3550 7588
rect 3422 7440 3478 7449
rect 3422 7375 3478 7384
rect 3436 7274 3464 7375
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3254 6556 3550 6576
rect 3310 6554 3334 6556
rect 3390 6554 3414 6556
rect 3470 6554 3494 6556
rect 3332 6502 3334 6554
rect 3396 6502 3408 6554
rect 3470 6502 3472 6554
rect 3310 6500 3334 6502
rect 3390 6500 3414 6502
rect 3470 6500 3494 6502
rect 3254 6480 3550 6500
rect 3424 6384 3476 6390
rect 3424 6326 3476 6332
rect 3160 6174 3280 6202
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5098 3188 6054
rect 3252 5556 3280 6174
rect 3436 5778 3464 6326
rect 3620 6322 3648 7822
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3252 5528 3648 5556
rect 3254 5468 3550 5488
rect 3310 5466 3334 5468
rect 3390 5466 3414 5468
rect 3470 5466 3494 5468
rect 3332 5414 3334 5466
rect 3396 5414 3408 5466
rect 3470 5414 3472 5466
rect 3310 5412 3334 5414
rect 3390 5412 3414 5414
rect 3470 5412 3494 5414
rect 3254 5392 3550 5412
rect 3514 5264 3570 5273
rect 3514 5199 3516 5208
rect 3568 5199 3570 5208
rect 3516 5170 3568 5176
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3146 4584 3202 4593
rect 3146 4519 3202 4528
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3068 3738 3096 3878
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 2962 2544 3018 2553
rect 2872 2508 2924 2514
rect 3160 2496 3188 4519
rect 3254 4380 3550 4400
rect 3310 4378 3334 4380
rect 3390 4378 3414 4380
rect 3470 4378 3494 4380
rect 3332 4326 3334 4378
rect 3396 4326 3408 4378
rect 3470 4326 3472 4378
rect 3310 4324 3334 4326
rect 3390 4324 3414 4326
rect 3470 4324 3494 4326
rect 3254 4304 3550 4324
rect 3620 4185 3648 5528
rect 3712 5234 3740 12718
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3804 8634 3832 11494
rect 3896 11257 3924 13359
rect 4804 13330 4856 13336
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3882 11248 3938 11257
rect 3882 11183 3938 11192
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3804 7546 3832 7890
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3804 6798 3832 7482
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3896 4690 3924 11018
rect 3976 11008 4028 11014
rect 3974 10976 3976 10985
rect 4028 10976 4030 10985
rect 3974 10911 4030 10920
rect 3974 10160 4030 10169
rect 3974 10095 4030 10104
rect 3988 9994 4016 10095
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 8566 4016 9454
rect 4080 9178 4108 11562
rect 4172 9568 4200 13126
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4250 12336 4306 12345
rect 4250 12271 4252 12280
rect 4304 12271 4306 12280
rect 4252 12242 4304 12248
rect 4264 11830 4292 12242
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4264 10470 4292 11018
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4264 10198 4292 10406
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4264 9722 4292 9930
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4172 9540 4292 9568
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4172 9110 4200 9386
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3988 8106 4016 8502
rect 4080 8294 4108 8774
rect 4264 8344 4292 9540
rect 4172 8316 4292 8344
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3988 8078 4108 8106
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3988 7857 4016 7958
rect 4080 7886 4108 8078
rect 4068 7880 4120 7886
rect 3974 7848 4030 7857
rect 4068 7822 4120 7828
rect 3974 7783 4030 7792
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3988 7177 4016 7278
rect 3974 7168 4030 7177
rect 3974 7103 4030 7112
rect 4080 7002 4108 7822
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4080 6497 4108 6938
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 4066 6216 4122 6225
rect 3976 6180 4028 6186
rect 4172 6202 4200 8316
rect 4356 7834 4384 11494
rect 4448 9042 4476 12582
rect 4710 12200 4766 12209
rect 4710 12135 4766 12144
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4356 7806 4476 7834
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4122 6174 4200 6202
rect 4066 6151 4122 6160
rect 3976 6122 4028 6128
rect 3988 5234 4016 6122
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5817 4108 6054
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4160 5704 4212 5710
rect 4080 5664 4160 5692
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4080 5114 4108 5664
rect 4160 5646 4212 5652
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 3988 5086 4108 5114
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3988 4622 4016 5086
rect 4066 4992 4122 5001
rect 4172 4978 4200 5510
rect 4122 4950 4200 4978
rect 4066 4927 4122 4936
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3882 4448 3938 4457
rect 3882 4383 3938 4392
rect 3606 4176 3662 4185
rect 3606 4111 3662 4120
rect 3700 3936 3752 3942
rect 3792 3936 3844 3942
rect 3700 3878 3752 3884
rect 3790 3904 3792 3913
rect 3844 3904 3846 3913
rect 3712 3670 3740 3878
rect 3790 3839 3846 3848
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3896 3534 3924 4383
rect 3988 3913 4016 4558
rect 4080 4146 4108 4694
rect 4264 4570 4292 7142
rect 4356 6254 4384 7686
rect 4448 7206 4476 7806
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 4448 6390 4476 6870
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4172 4542 4292 4570
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3974 3904 4030 3913
rect 3974 3839 4030 3848
rect 3974 3768 4030 3777
rect 4080 3738 4108 4082
rect 3974 3703 4030 3712
rect 4068 3732 4120 3738
rect 3988 3602 4016 3703
rect 4068 3674 4120 3680
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3254 3292 3550 3312
rect 3310 3290 3334 3292
rect 3390 3290 3414 3292
rect 3470 3290 3494 3292
rect 3332 3238 3334 3290
rect 3396 3238 3408 3290
rect 3470 3238 3472 3290
rect 3310 3236 3334 3238
rect 3390 3236 3414 3238
rect 3470 3236 3494 3238
rect 3254 3216 3550 3236
rect 3620 3176 3648 3334
rect 3344 3148 3648 3176
rect 3344 2922 3372 3148
rect 4066 2952 4122 2961
rect 3332 2916 3384 2922
rect 4172 2938 4200 4542
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4264 3398 4292 4422
rect 4342 4312 4398 4321
rect 4342 4247 4398 4256
rect 4356 4078 4384 4247
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4356 2990 4384 3878
rect 4448 3058 4476 5102
rect 4540 3942 4568 11834
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4632 9518 4660 9998
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 8974 4660 9318
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4632 8498 4660 8910
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4632 7546 4660 8230
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4724 7478 4752 12135
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4816 6882 4844 12038
rect 4908 8430 4936 13330
rect 5092 12646 5120 13942
rect 5184 12986 5212 15520
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5276 13394 5304 13874
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4908 7410 4936 7890
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 7002 4936 7142
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4632 6854 4844 6882
rect 4632 6118 4660 6854
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4540 3398 4568 3606
rect 4632 3534 4660 5170
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4526 3224 4582 3233
rect 4526 3159 4582 3168
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4540 2990 4568 3159
rect 4122 2910 4200 2938
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4066 2887 4122 2896
rect 3332 2858 3384 2864
rect 4632 2854 4660 3334
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4172 2666 4200 2790
rect 4172 2638 4476 2666
rect 2962 2479 3018 2488
rect 2872 2450 2924 2456
rect 3068 2468 3188 2496
rect 3698 2544 3754 2553
rect 4448 2530 4476 2638
rect 4632 2553 4660 2790
rect 4618 2544 4674 2553
rect 4448 2514 4568 2530
rect 3698 2479 3754 2488
rect 4068 2508 4120 2514
rect 2884 2417 2912 2450
rect 2870 2408 2926 2417
rect 3068 2378 3096 2468
rect 3712 2446 3740 2479
rect 4448 2508 4580 2514
rect 4448 2502 4528 2508
rect 4068 2450 4120 2456
rect 4618 2479 4674 2488
rect 4528 2450 4580 2456
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 2870 2343 2926 2352
rect 3056 2372 3108 2378
rect 3056 2314 3108 2320
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2884 1834 2912 2246
rect 3254 2204 3550 2224
rect 3310 2202 3334 2204
rect 3390 2202 3414 2204
rect 3470 2202 3494 2204
rect 3332 2150 3334 2202
rect 3396 2150 3408 2202
rect 3470 2150 3472 2202
rect 3310 2148 3334 2150
rect 3390 2148 3414 2150
rect 3470 2148 3494 2150
rect 3054 2136 3110 2145
rect 3254 2128 3550 2148
rect 3620 2106 3648 2314
rect 3054 2071 3110 2080
rect 3608 2100 3660 2106
rect 3068 1902 3096 2071
rect 3608 2042 3660 2048
rect 4080 1970 4108 2450
rect 4620 2440 4672 2446
rect 4618 2408 4620 2417
rect 4672 2408 4674 2417
rect 4618 2343 4674 2352
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 3056 1896 3108 1902
rect 3056 1838 3108 1844
rect 2872 1828 2924 1834
rect 2872 1770 2924 1776
rect 3056 1488 3108 1494
rect 3056 1430 3108 1436
rect 2688 1012 2740 1018
rect 2688 954 2740 960
rect 2780 808 2832 814
rect 2780 750 2832 756
rect 2792 513 2820 750
rect 2872 740 2924 746
rect 2872 682 2924 688
rect 2778 504 2834 513
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 2778 439 2834 448
rect 2884 241 2912 682
rect 3068 480 3096 1430
rect 3608 1012 3660 1018
rect 3608 954 3660 960
rect 3620 480 3648 954
rect 4172 480 4200 2246
rect 4724 480 4752 6666
rect 4802 6488 4858 6497
rect 4802 6423 4858 6432
rect 4816 6390 4844 6423
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4816 5370 4844 6054
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4908 5370 4936 5782
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4816 3942 4844 4966
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4816 3040 4844 3674
rect 4908 3398 4936 5034
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4896 3052 4948 3058
rect 4816 3012 4896 3040
rect 4896 2994 4948 3000
rect 4896 2848 4948 2854
rect 4894 2816 4896 2825
rect 4948 2816 4950 2825
rect 4894 2751 4950 2760
rect 5000 626 5028 12310
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5184 12209 5212 12242
rect 5170 12200 5226 12209
rect 5170 12135 5226 12144
rect 5078 11792 5134 11801
rect 5078 11727 5080 11736
rect 5132 11727 5134 11736
rect 5080 11698 5132 11704
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5092 8945 5120 9522
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5078 8936 5134 8945
rect 5078 8871 5134 8880
rect 5078 8528 5134 8537
rect 5078 8463 5134 8472
rect 5092 7410 5120 8463
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5092 6769 5120 7346
rect 5184 7206 5212 9454
rect 5276 8022 5304 10406
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5078 6760 5134 6769
rect 5078 6695 5134 6704
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 4706 5120 6598
rect 5276 5794 5304 7414
rect 5368 7342 5396 13126
rect 5460 9518 5488 13806
rect 5553 13628 5849 13648
rect 5609 13626 5633 13628
rect 5689 13626 5713 13628
rect 5769 13626 5793 13628
rect 5631 13574 5633 13626
rect 5695 13574 5707 13626
rect 5769 13574 5771 13626
rect 5609 13572 5633 13574
rect 5689 13572 5713 13574
rect 5769 13572 5793 13574
rect 5553 13552 5849 13572
rect 5553 12540 5849 12560
rect 5609 12538 5633 12540
rect 5689 12538 5713 12540
rect 5769 12538 5793 12540
rect 5631 12486 5633 12538
rect 5695 12486 5707 12538
rect 5769 12486 5771 12538
rect 5609 12484 5633 12486
rect 5689 12484 5713 12486
rect 5769 12484 5793 12486
rect 5553 12464 5849 12484
rect 5920 11898 5948 15520
rect 6458 15464 6514 15473
rect 6458 15399 6514 15408
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5553 11452 5849 11472
rect 5609 11450 5633 11452
rect 5689 11450 5713 11452
rect 5769 11450 5793 11452
rect 5631 11398 5633 11450
rect 5695 11398 5707 11450
rect 5769 11398 5771 11450
rect 5609 11396 5633 11398
rect 5689 11396 5713 11398
rect 5769 11396 5793 11398
rect 5553 11376 5849 11396
rect 5920 11234 5948 11630
rect 5828 11206 5948 11234
rect 5828 10742 5856 11206
rect 6012 10826 6040 12582
rect 6104 12345 6132 12786
rect 6090 12336 6146 12345
rect 6090 12271 6146 12280
rect 6196 11830 6224 13670
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6472 11354 6500 15399
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6656 11762 6684 12378
rect 6748 12102 6776 15520
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6458 11248 6514 11257
rect 6458 11183 6514 11192
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 5920 10798 6040 10826
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5553 10364 5849 10384
rect 5609 10362 5633 10364
rect 5689 10362 5713 10364
rect 5769 10362 5793 10364
rect 5631 10310 5633 10362
rect 5695 10310 5707 10362
rect 5769 10310 5771 10362
rect 5609 10308 5633 10310
rect 5689 10308 5713 10310
rect 5769 10308 5793 10310
rect 5553 10288 5849 10308
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5828 9722 5856 9930
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5553 9276 5849 9296
rect 5609 9274 5633 9276
rect 5689 9274 5713 9276
rect 5769 9274 5793 9276
rect 5631 9222 5633 9274
rect 5695 9222 5707 9274
rect 5769 9222 5771 9274
rect 5609 9220 5633 9222
rect 5689 9220 5713 9222
rect 5769 9220 5793 9222
rect 5553 9200 5849 9220
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5460 8090 5488 9046
rect 5828 8974 5856 9046
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5920 8906 5948 10798
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 6012 9926 6040 10678
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5553 8188 5849 8208
rect 5609 8186 5633 8188
rect 5689 8186 5713 8188
rect 5769 8186 5793 8188
rect 5631 8134 5633 8186
rect 5695 8134 5707 8186
rect 5769 8134 5771 8186
rect 5609 8132 5633 8134
rect 5689 8132 5713 8134
rect 5769 8132 5793 8134
rect 5553 8112 5849 8132
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5460 7410 5488 8026
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5354 5808 5410 5817
rect 5276 5766 5354 5794
rect 5354 5743 5410 5752
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5276 5370 5304 5646
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5184 4826 5212 5170
rect 5368 5166 5396 5743
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5262 4856 5318 4865
rect 5172 4820 5224 4826
rect 5262 4791 5318 4800
rect 5172 4762 5224 4768
rect 5092 4678 5212 4706
rect 5276 4690 5304 4791
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5092 4078 5120 4150
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 3097 5120 3334
rect 5078 3088 5134 3097
rect 5078 3023 5134 3032
rect 5184 814 5212 4678
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5264 4072 5316 4078
rect 5262 4040 5264 4049
rect 5316 4040 5318 4049
rect 5262 3975 5318 3984
rect 5368 3126 5396 4966
rect 5460 3738 5488 7210
rect 5553 7100 5849 7120
rect 5609 7098 5633 7100
rect 5689 7098 5713 7100
rect 5769 7098 5793 7100
rect 5631 7046 5633 7098
rect 5695 7046 5707 7098
rect 5769 7046 5771 7098
rect 5609 7044 5633 7046
rect 5689 7044 5713 7046
rect 5769 7044 5793 7046
rect 5553 7024 5849 7044
rect 5920 6662 5948 8434
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5553 6012 5849 6032
rect 5609 6010 5633 6012
rect 5689 6010 5713 6012
rect 5769 6010 5793 6012
rect 5631 5958 5633 6010
rect 5695 5958 5707 6010
rect 5769 5958 5771 6010
rect 5609 5956 5633 5958
rect 5689 5956 5713 5958
rect 5769 5956 5793 5958
rect 5553 5936 5849 5956
rect 5920 5166 5948 6598
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5553 4924 5849 4944
rect 5609 4922 5633 4924
rect 5689 4922 5713 4924
rect 5769 4922 5793 4924
rect 5631 4870 5633 4922
rect 5695 4870 5707 4922
rect 5769 4870 5771 4922
rect 5609 4868 5633 4870
rect 5689 4868 5713 4870
rect 5769 4868 5793 4870
rect 5553 4848 5849 4868
rect 6012 4758 6040 6054
rect 6104 5953 6132 10474
rect 6196 9722 6224 10610
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6090 5944 6146 5953
rect 6090 5879 6146 5888
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5816 4616 5868 4622
rect 5814 4584 5816 4593
rect 5868 4584 5870 4593
rect 5814 4519 5870 4528
rect 5553 3836 5849 3856
rect 5609 3834 5633 3836
rect 5689 3834 5713 3836
rect 5769 3834 5793 3836
rect 5631 3782 5633 3834
rect 5695 3782 5707 3834
rect 5769 3782 5771 3834
rect 5609 3780 5633 3782
rect 5689 3780 5713 3782
rect 5769 3780 5793 3782
rect 5553 3760 5849 3780
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 3505 5488 3538
rect 5446 3496 5502 3505
rect 5446 3431 5502 3440
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5552 3058 5580 3606
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5920 2990 5948 4694
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 5460 1494 5488 2858
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5553 2748 5849 2768
rect 5609 2746 5633 2748
rect 5689 2746 5713 2748
rect 5769 2746 5793 2748
rect 5631 2694 5633 2746
rect 5695 2694 5707 2746
rect 5769 2694 5771 2746
rect 5609 2692 5633 2694
rect 5689 2692 5713 2694
rect 5769 2692 5793 2694
rect 5553 2672 5849 2692
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 5644 2446 5672 2518
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5448 1488 5500 1494
rect 5448 1430 5500 1436
rect 5172 808 5224 814
rect 5172 750 5224 756
rect 5920 746 5948 2790
rect 6012 2650 6040 2858
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5908 740 5960 746
rect 5908 682 5960 688
rect 6104 626 6132 5510
rect 6196 4570 6224 9658
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6288 9042 6316 9590
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6288 6118 6316 7210
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6274 5944 6330 5953
rect 6274 5879 6330 5888
rect 6288 4690 6316 5879
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6196 4542 6316 4570
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6196 2514 6224 4082
rect 6288 3466 6316 4542
rect 6380 3534 6408 11018
rect 6472 7274 6500 11183
rect 6564 8090 6592 11698
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6472 5846 6500 6394
rect 6550 6352 6606 6361
rect 6550 6287 6606 6296
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6458 5400 6514 5409
rect 6458 5335 6514 5344
rect 6472 5030 6500 5335
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6288 2038 6316 2246
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 5000 598 5304 626
rect 5276 480 5304 598
rect 5828 598 6132 626
rect 5828 480 5856 598
rect 6380 480 6408 2790
rect 6564 2378 6592 6287
rect 6656 2446 6684 11494
rect 6840 11218 6868 15030
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 6920 14204 6972 14210
rect 6920 14146 6972 14152
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6748 5778 6776 11018
rect 6840 8430 6868 11154
rect 6932 8430 6960 14146
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 7024 12374 7052 12718
rect 7116 12442 7144 13330
rect 7300 12918 7328 14214
rect 7576 13410 7604 15520
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7576 13382 7696 13410
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7288 12912 7340 12918
rect 7288 12854 7340 12860
rect 7194 12744 7250 12753
rect 7194 12679 7250 12688
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7208 12374 7236 12679
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7024 10305 7052 11630
rect 7116 10577 7144 12174
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7102 10568 7158 10577
rect 7102 10503 7158 10512
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7010 10296 7066 10305
rect 7010 10231 7066 10240
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 7024 9518 7052 10134
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7024 9178 7052 9454
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6840 6866 6868 8026
rect 6932 8022 6960 8366
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6748 5302 6776 5510
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6748 4729 6776 5238
rect 6734 4720 6790 4729
rect 6734 4655 6790 4664
rect 6840 3602 6868 5306
rect 6932 4078 6960 7686
rect 7024 6934 7052 8978
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 7024 4282 7052 5782
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6840 2514 6868 3538
rect 6932 2990 6960 3878
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 7116 2106 7144 10406
rect 7208 10266 7236 11834
rect 7392 11132 7420 13126
rect 7576 12322 7604 13262
rect 7668 12782 7696 13382
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7484 12294 7604 12322
rect 7484 11898 7512 12294
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7576 11762 7604 12174
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7300 11104 7420 11132
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 9586 7236 9998
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7194 9480 7250 9489
rect 7300 9466 7328 11104
rect 7484 10588 7512 11494
rect 7576 10674 7604 11698
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7392 10560 7512 10588
rect 7392 9654 7420 10560
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7484 10130 7512 10202
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7484 9489 7512 10066
rect 7576 9625 7604 10406
rect 7562 9616 7618 9625
rect 7562 9551 7618 9560
rect 7564 9512 7616 9518
rect 7470 9480 7526 9489
rect 7300 9438 7420 9466
rect 7194 9415 7250 9424
rect 7208 5098 7236 9415
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 6066 7328 9318
rect 7392 8294 7420 9438
rect 7564 9454 7616 9460
rect 7470 9415 7526 9424
rect 7470 9344 7526 9353
rect 7470 9279 7526 9288
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7546 7420 7822
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7484 7478 7512 9279
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7300 6038 7420 6066
rect 7286 5672 7342 5681
rect 7286 5607 7342 5616
rect 7300 5234 7328 5607
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7286 5128 7342 5137
rect 7196 5092 7248 5098
rect 7286 5063 7288 5072
rect 7196 5034 7248 5040
rect 7340 5063 7342 5072
rect 7288 5034 7340 5040
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 4146 7328 4422
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7300 2582 7328 2926
rect 7288 2576 7340 2582
rect 7288 2518 7340 2524
rect 7104 2100 7156 2106
rect 7104 2042 7156 2048
rect 7392 1902 7420 6038
rect 7484 4826 7512 7414
rect 7576 7342 7604 9454
rect 7668 9058 7696 11086
rect 7760 9178 7788 13806
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 7852 13084 8148 13104
rect 7908 13082 7932 13084
rect 7988 13082 8012 13084
rect 8068 13082 8092 13084
rect 7930 13030 7932 13082
rect 7994 13030 8006 13082
rect 8068 13030 8070 13082
rect 7908 13028 7932 13030
rect 7988 13028 8012 13030
rect 8068 13028 8092 13030
rect 7852 13008 8148 13028
rect 8220 12424 8248 13398
rect 8220 12396 8340 12424
rect 7852 11996 8148 12016
rect 7908 11994 7932 11996
rect 7988 11994 8012 11996
rect 8068 11994 8092 11996
rect 7930 11942 7932 11994
rect 7994 11942 8006 11994
rect 8068 11942 8070 11994
rect 7908 11940 7932 11942
rect 7988 11940 8012 11942
rect 8068 11940 8092 11942
rect 7852 11920 8148 11940
rect 7852 10908 8148 10928
rect 7908 10906 7932 10908
rect 7988 10906 8012 10908
rect 8068 10906 8092 10908
rect 7930 10854 7932 10906
rect 7994 10854 8006 10906
rect 8068 10854 8070 10906
rect 7908 10852 7932 10854
rect 7988 10852 8012 10854
rect 8068 10852 8092 10854
rect 7852 10832 8148 10852
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8036 10130 8064 10610
rect 8206 10568 8262 10577
rect 8206 10503 8262 10512
rect 8220 10130 8248 10503
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8312 10010 8340 12396
rect 8404 12374 8432 15520
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8496 12442 8524 14010
rect 9140 13512 9168 15520
rect 8772 13484 9168 13512
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8482 12336 8538 12345
rect 8482 12271 8538 12280
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8404 10606 8432 11562
rect 8496 11150 8524 12271
rect 8772 11540 8800 13484
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8864 11778 8892 13194
rect 8942 12744 8998 12753
rect 8942 12679 8998 12688
rect 8956 12170 8984 12679
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 8944 12164 8996 12170
rect 8944 12106 8996 12112
rect 9048 12102 9076 12242
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8864 11750 8984 11778
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8680 11512 8800 11540
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8588 10674 8616 11086
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8220 9982 8340 10010
rect 7852 9820 8148 9840
rect 7908 9818 7932 9820
rect 7988 9818 8012 9820
rect 8068 9818 8092 9820
rect 7930 9766 7932 9818
rect 7994 9766 8006 9818
rect 8068 9766 8070 9818
rect 7908 9764 7932 9766
rect 7988 9764 8012 9766
rect 8068 9764 8092 9766
rect 7852 9744 8148 9764
rect 7748 9172 7800 9178
rect 8220 9160 8248 9982
rect 8588 9518 8616 10202
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8576 9172 8628 9178
rect 8220 9132 8432 9160
rect 7748 9114 7800 9120
rect 7668 9030 7788 9058
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7668 8498 7696 8910
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7668 7886 7696 8434
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7576 3602 7604 6802
rect 7668 6118 7696 7822
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7668 4622 7696 6054
rect 7760 5137 7788 9030
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 7852 8732 8148 8752
rect 7908 8730 7932 8732
rect 7988 8730 8012 8732
rect 8068 8730 8092 8732
rect 7930 8678 7932 8730
rect 7994 8678 8006 8730
rect 8068 8678 8070 8730
rect 7908 8676 7932 8678
rect 7988 8676 8012 8678
rect 8068 8676 8092 8678
rect 7852 8656 8148 8676
rect 7852 7644 8148 7664
rect 7908 7642 7932 7644
rect 7988 7642 8012 7644
rect 8068 7642 8092 7644
rect 7930 7590 7932 7642
rect 7994 7590 8006 7642
rect 8068 7590 8070 7642
rect 7908 7588 7932 7590
rect 7988 7588 8012 7590
rect 8068 7588 8092 7590
rect 7852 7568 8148 7588
rect 8220 7528 8248 8978
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8128 7500 8248 7528
rect 8128 6934 8156 7500
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8220 6730 8248 7346
rect 8312 7206 8340 8842
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 7852 6556 8148 6576
rect 7908 6554 7932 6556
rect 7988 6554 8012 6556
rect 8068 6554 8092 6556
rect 7930 6502 7932 6554
rect 7994 6502 8006 6554
rect 8068 6502 8070 6554
rect 7908 6500 7932 6502
rect 7988 6500 8012 6502
rect 8068 6500 8092 6502
rect 7852 6480 8148 6500
rect 8220 6186 8248 6666
rect 8312 6390 8340 7142
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8312 5914 8340 6122
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 7852 5468 8148 5488
rect 7908 5466 7932 5468
rect 7988 5466 8012 5468
rect 8068 5466 8092 5468
rect 7930 5414 7932 5466
rect 7994 5414 8006 5466
rect 8068 5414 8070 5466
rect 7908 5412 7932 5414
rect 7988 5412 8012 5414
rect 8068 5412 8092 5414
rect 7852 5392 8148 5412
rect 7746 5128 7802 5137
rect 7746 5063 7802 5072
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4826 7788 4966
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7852 4380 8148 4400
rect 7908 4378 7932 4380
rect 7988 4378 8012 4380
rect 8068 4378 8092 4380
rect 7930 4326 7932 4378
rect 7994 4326 8006 4378
rect 8068 4326 8070 4378
rect 7908 4324 7932 4326
rect 7988 4324 8012 4326
rect 8068 4324 8092 4326
rect 7852 4304 8148 4324
rect 8220 3602 8248 5510
rect 8312 5098 8340 5646
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8404 3670 8432 9132
rect 8576 9114 8628 9120
rect 8588 9081 8616 9114
rect 8574 9072 8630 9081
rect 8574 9007 8630 9016
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8496 8362 8524 8774
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 4826 8524 6598
rect 8588 5710 8616 9007
rect 8680 7993 8708 11512
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8666 7984 8722 7993
rect 8666 7919 8722 7928
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8680 6361 8708 7278
rect 8666 6352 8722 6361
rect 8666 6287 8722 6296
rect 8666 6080 8722 6089
rect 8666 6015 8722 6024
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8680 5574 8708 6015
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8666 4720 8722 4729
rect 8666 4655 8722 4664
rect 8680 4078 8708 4655
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8300 3664 8352 3670
rect 8300 3606 8352 3612
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 7852 3292 8148 3312
rect 7908 3290 7932 3292
rect 7988 3290 8012 3292
rect 8068 3290 8092 3292
rect 7930 3238 7932 3290
rect 7994 3238 8006 3290
rect 8068 3238 8070 3290
rect 7908 3236 7932 3238
rect 7988 3236 8012 3238
rect 8068 3236 8092 3238
rect 7852 3216 8148 3236
rect 8220 2990 8248 3334
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 7380 1896 7432 1902
rect 7380 1838 7432 1844
rect 6920 1420 6972 1426
rect 6920 1362 6972 1368
rect 6932 480 6960 1362
rect 7484 480 7512 2790
rect 7852 2204 8148 2224
rect 7908 2202 7932 2204
rect 7988 2202 8012 2204
rect 8068 2202 8092 2204
rect 7930 2150 7932 2202
rect 7994 2150 8006 2202
rect 8068 2150 8070 2202
rect 7908 2148 7932 2150
rect 7988 2148 8012 2150
rect 8068 2148 8092 2150
rect 7852 2128 8148 2148
rect 8220 1986 8248 2790
rect 8312 2650 8340 3606
rect 8496 2922 8524 4014
rect 8772 2961 8800 10406
rect 8758 2952 8814 2961
rect 8484 2916 8536 2922
rect 8758 2887 8814 2896
rect 8484 2858 8536 2864
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8036 1958 8248 1986
rect 8036 480 8064 1958
rect 8588 480 8616 2246
rect 8864 1834 8892 11630
rect 8956 11558 8984 11750
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8956 10674 8984 11018
rect 9048 10674 9076 11698
rect 9140 10810 9168 13330
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9232 11898 9260 13262
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9324 11762 9352 13126
rect 9784 12889 9812 13126
rect 9770 12880 9826 12889
rect 9770 12815 9826 12824
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9862 12744 9918 12753
rect 9692 12322 9720 12718
rect 9862 12679 9864 12688
rect 9916 12679 9918 12688
rect 9864 12650 9916 12656
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 12442 9812 12582
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9600 12294 9720 12322
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9220 11688 9272 11694
rect 9600 11676 9628 12294
rect 9680 12164 9732 12170
rect 9732 12124 9904 12152
rect 9680 12106 9732 12112
rect 9678 12064 9734 12073
rect 9678 11999 9734 12008
rect 9692 11830 9720 11999
rect 9876 11898 9904 12124
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9600 11648 9720 11676
rect 9220 11630 9272 11636
rect 9232 11218 9260 11630
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9048 10266 9076 10610
rect 9324 10606 9352 10950
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9126 10296 9182 10305
rect 9036 10260 9088 10266
rect 9126 10231 9128 10240
rect 9036 10202 9088 10208
rect 9180 10231 9182 10240
rect 9128 10202 9180 10208
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9324 10033 9352 10066
rect 9310 10024 9366 10033
rect 9310 9959 9366 9968
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 6882 8984 8434
rect 9048 8362 9076 8502
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9140 7313 9168 8434
rect 9126 7304 9182 7313
rect 9126 7239 9182 7248
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 8956 6854 9076 6882
rect 8944 6792 8996 6798
rect 8942 6760 8944 6769
rect 8996 6760 8998 6769
rect 8942 6695 8998 6704
rect 9048 6458 9076 6854
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 8956 4826 8984 6326
rect 9034 5264 9090 5273
rect 9034 5199 9090 5208
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9048 4078 9076 5199
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8956 3505 8984 3946
rect 8942 3496 8998 3505
rect 8942 3431 8998 3440
rect 8852 1828 8904 1834
rect 8852 1770 8904 1776
rect 9140 480 9168 7142
rect 9232 5846 9260 8842
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9324 6458 9352 6734
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9220 5228 9272 5234
rect 9324 5216 9352 6394
rect 9272 5188 9352 5216
rect 9220 5170 9272 5176
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9324 2836 9352 4762
rect 9416 2990 9444 11494
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9508 6866 9536 10678
rect 9692 10554 9720 11648
rect 9784 11218 9812 11766
rect 9772 11212 9824 11218
rect 9968 11200 9996 15520
rect 10690 13832 10746 13841
rect 10690 13767 10746 13776
rect 10150 13628 10446 13648
rect 10206 13626 10230 13628
rect 10286 13626 10310 13628
rect 10366 13626 10390 13628
rect 10228 13574 10230 13626
rect 10292 13574 10304 13626
rect 10366 13574 10368 13626
rect 10206 13572 10230 13574
rect 10286 13572 10310 13574
rect 10366 13572 10390 13574
rect 10150 13552 10446 13572
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 10060 11830 10088 13194
rect 10150 12540 10446 12560
rect 10206 12538 10230 12540
rect 10286 12538 10310 12540
rect 10366 12538 10390 12540
rect 10228 12486 10230 12538
rect 10292 12486 10304 12538
rect 10366 12486 10368 12538
rect 10206 12484 10230 12486
rect 10286 12484 10310 12486
rect 10366 12484 10390 12486
rect 10150 12464 10446 12484
rect 10520 12102 10548 13330
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10150 11452 10446 11472
rect 10206 11450 10230 11452
rect 10286 11450 10310 11452
rect 10366 11450 10390 11452
rect 10228 11398 10230 11450
rect 10292 11398 10304 11450
rect 10366 11398 10368 11450
rect 10206 11396 10230 11398
rect 10286 11396 10310 11398
rect 10366 11396 10390 11398
rect 10150 11376 10446 11396
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 9772 11154 9824 11160
rect 9876 11172 9996 11200
rect 9600 10526 9720 10554
rect 9600 6866 9628 10526
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6322 9536 6598
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9508 5642 9536 6258
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9600 5953 9628 6190
rect 9586 5944 9642 5953
rect 9586 5879 9642 5888
rect 9586 5808 9642 5817
rect 9586 5743 9642 5752
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9508 5370 9536 5578
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9508 4282 9536 5306
rect 9600 5234 9628 5743
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9508 2836 9536 2926
rect 9324 2808 9536 2836
rect 9600 1358 9628 4490
rect 9692 3777 9720 10406
rect 9784 9654 9812 11154
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8430 9812 8774
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9784 5166 9812 8366
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9678 3768 9734 3777
rect 9678 3703 9734 3712
rect 9784 3670 9812 4150
rect 9876 3738 9904 11172
rect 10152 11098 10180 11222
rect 9968 11070 10180 11098
rect 9968 7274 9996 11070
rect 10150 10364 10446 10384
rect 10206 10362 10230 10364
rect 10286 10362 10310 10364
rect 10366 10362 10390 10364
rect 10228 10310 10230 10362
rect 10292 10310 10304 10362
rect 10366 10310 10368 10362
rect 10206 10308 10230 10310
rect 10286 10308 10310 10310
rect 10366 10308 10390 10310
rect 10150 10288 10446 10308
rect 10048 10192 10100 10198
rect 10046 10160 10048 10169
rect 10100 10160 10102 10169
rect 10046 10095 10102 10104
rect 10046 9752 10102 9761
rect 10046 9687 10102 9696
rect 10060 9586 10088 9687
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10060 9042 10088 9522
rect 10150 9276 10446 9296
rect 10206 9274 10230 9276
rect 10286 9274 10310 9276
rect 10366 9274 10390 9276
rect 10228 9222 10230 9274
rect 10292 9222 10304 9274
rect 10366 9222 10368 9274
rect 10206 9220 10230 9222
rect 10286 9220 10310 9222
rect 10366 9220 10390 9222
rect 10150 9200 10446 9220
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10060 8294 10088 8978
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10428 8430 10456 8570
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 8090 10088 8230
rect 10150 8188 10446 8208
rect 10206 8186 10230 8188
rect 10286 8186 10310 8188
rect 10366 8186 10390 8188
rect 10228 8134 10230 8186
rect 10292 8134 10304 8186
rect 10366 8134 10368 8186
rect 10206 8132 10230 8134
rect 10286 8132 10310 8134
rect 10366 8132 10390 8134
rect 10150 8112 10446 8132
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10140 7880 10192 7886
rect 10060 7840 10140 7868
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 10060 7018 10088 7840
rect 10140 7822 10192 7828
rect 10520 7290 10548 12038
rect 10612 11268 10640 13398
rect 10704 12374 10732 13767
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 10704 12209 10732 12310
rect 10690 12200 10746 12209
rect 10690 12135 10746 12144
rect 10796 11558 10824 15520
rect 11058 15056 11114 15065
rect 11058 14991 11114 15000
rect 11072 13938 11100 14991
rect 11242 14648 11298 14657
rect 11242 14583 11298 14592
rect 11150 14240 11206 14249
rect 11150 14175 11206 14184
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 11164 13870 11192 14175
rect 11256 14006 11284 14583
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11532 13530 11560 15520
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11242 12880 11298 12889
rect 11060 12844 11112 12850
rect 11242 12815 11298 12824
rect 11060 12786 11112 12792
rect 10968 12640 11020 12646
rect 11072 12617 11100 12786
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 10968 12582 11020 12588
rect 11058 12608 11114 12617
rect 10980 12073 11008 12582
rect 11058 12543 11114 12552
rect 11058 12200 11114 12209
rect 11058 12135 11114 12144
rect 10966 12064 11022 12073
rect 10966 11999 11022 12008
rect 11072 11914 11100 12135
rect 10888 11886 11100 11914
rect 10888 11626 10916 11886
rect 11058 11792 11114 11801
rect 11058 11727 11060 11736
rect 11112 11727 11114 11736
rect 11060 11698 11112 11704
rect 11164 11694 11192 12650
rect 11256 12345 11284 12815
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11242 12336 11298 12345
rect 11348 12306 11376 12718
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11242 12271 11298 12280
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 11058 11384 11114 11393
rect 11058 11319 11114 11328
rect 10612 11240 10916 11268
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10612 7546 10640 9862
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10520 7262 10640 7290
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10150 7100 10446 7120
rect 10206 7098 10230 7100
rect 10286 7098 10310 7100
rect 10366 7098 10390 7100
rect 10228 7046 10230 7098
rect 10292 7046 10304 7098
rect 10366 7046 10368 7098
rect 10206 7044 10230 7046
rect 10286 7044 10310 7046
rect 10366 7044 10390 7046
rect 10150 7024 10446 7044
rect 9968 6990 10088 7018
rect 9968 6118 9996 6990
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9968 5370 9996 5850
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9968 3584 9996 5034
rect 10060 4146 10088 6802
rect 10150 6012 10446 6032
rect 10206 6010 10230 6012
rect 10286 6010 10310 6012
rect 10366 6010 10390 6012
rect 10228 5958 10230 6010
rect 10292 5958 10304 6010
rect 10366 5958 10368 6010
rect 10206 5956 10230 5958
rect 10286 5956 10310 5958
rect 10366 5956 10390 5958
rect 10150 5936 10446 5956
rect 10520 5370 10548 7142
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10138 5264 10194 5273
rect 10138 5199 10194 5208
rect 10232 5228 10284 5234
rect 10152 5098 10180 5199
rect 10232 5170 10284 5176
rect 10244 5137 10272 5170
rect 10336 5166 10364 5306
rect 10324 5160 10376 5166
rect 10230 5128 10286 5137
rect 10140 5092 10192 5098
rect 10324 5102 10376 5108
rect 10230 5063 10286 5072
rect 10140 5034 10192 5040
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10150 4924 10446 4944
rect 10206 4922 10230 4924
rect 10286 4922 10310 4924
rect 10366 4922 10390 4924
rect 10228 4870 10230 4922
rect 10292 4870 10304 4922
rect 10366 4870 10368 4922
rect 10206 4868 10230 4870
rect 10286 4868 10310 4870
rect 10366 4868 10390 4870
rect 10150 4848 10446 4868
rect 10520 4826 10548 4966
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10428 4282 10456 4626
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10150 3836 10446 3856
rect 10206 3834 10230 3836
rect 10286 3834 10310 3836
rect 10366 3834 10390 3836
rect 10228 3782 10230 3834
rect 10292 3782 10304 3834
rect 10366 3782 10368 3834
rect 10206 3780 10230 3782
rect 10286 3780 10310 3782
rect 10366 3780 10390 3782
rect 10150 3760 10446 3780
rect 10048 3732 10100 3738
rect 10100 3692 10180 3720
rect 10048 3674 10100 3680
rect 10048 3596 10100 3602
rect 9968 3556 10048 3584
rect 10048 3538 10100 3544
rect 9680 3460 9732 3466
rect 9784 3454 9996 3482
rect 9784 3448 9812 3454
rect 9732 3420 9812 3448
rect 9680 3402 9732 3408
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9678 2952 9734 2961
rect 9678 2887 9734 2896
rect 9692 2854 9720 2887
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9876 2666 9904 3334
rect 9692 2638 9904 2666
rect 9588 1352 9640 1358
rect 9588 1294 9640 1300
rect 9692 480 9720 2638
rect 9968 2582 9996 3454
rect 10152 3194 10180 3692
rect 10612 3398 10640 7262
rect 10704 4826 10732 11086
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8634 10824 8774
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10888 7886 10916 11240
rect 11072 11218 11100 11319
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10980 10130 11008 10950
rect 11058 10704 11114 10713
rect 11058 10639 11060 10648
rect 11112 10639 11114 10648
rect 11060 10610 11112 10616
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 9761 11008 10066
rect 10966 9752 11022 9761
rect 11164 9722 11192 10542
rect 10966 9687 11022 9696
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11058 9344 11114 9353
rect 11058 9279 11114 9288
rect 11072 9178 11100 9279
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11348 8673 11376 12242
rect 11440 9194 11468 12310
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11532 10112 11560 11698
rect 11624 11558 11652 15807
rect 11900 15558 12112 15586
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 10470 11652 11494
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11716 10538 11744 10610
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11612 10124 11664 10130
rect 11532 10084 11612 10112
rect 11612 10066 11664 10072
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11624 9382 11652 10066
rect 11716 10033 11744 10066
rect 11702 10024 11758 10033
rect 11702 9959 11758 9968
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11440 9166 11652 9194
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11334 8664 11390 8673
rect 11334 8599 11390 8608
rect 11426 8528 11482 8537
rect 11336 8492 11388 8498
rect 11426 8463 11482 8472
rect 11336 8434 11388 8440
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10876 7880 10928 7886
rect 11072 7857 11100 8230
rect 10876 7822 10928 7828
rect 11058 7848 11114 7857
rect 10968 7812 11020 7818
rect 11058 7783 11114 7792
rect 10968 7754 11020 7760
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10796 6866 10824 7346
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10796 4758 10824 6802
rect 10888 6225 10916 7686
rect 10980 6882 11008 7754
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11072 7313 11100 7414
rect 11058 7304 11114 7313
rect 11058 7239 11114 7248
rect 11058 6896 11114 6905
rect 10980 6854 11058 6882
rect 11058 6831 11114 6840
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10874 6216 10930 6225
rect 10874 6151 10930 6160
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10796 3058 10824 4082
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10150 2748 10446 2768
rect 10206 2746 10230 2748
rect 10286 2746 10310 2748
rect 10366 2746 10390 2748
rect 10228 2694 10230 2746
rect 10292 2694 10304 2746
rect 10366 2694 10368 2746
rect 10206 2692 10230 2694
rect 10286 2692 10310 2694
rect 10366 2692 10390 2694
rect 10150 2672 10446 2692
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9968 1426 9996 2246
rect 9956 1420 10008 1426
rect 9956 1362 10008 1368
rect 10244 480 10272 2450
rect 10796 480 10824 2994
rect 10888 2514 10916 6054
rect 10980 5778 11008 6666
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11072 5914 11100 6122
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10980 5234 11008 5714
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 11072 3890 11100 5238
rect 11164 4826 11192 8298
rect 11348 6730 11376 8434
rect 11440 7002 11468 8463
rect 11532 8022 11560 8842
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11532 7041 11560 7482
rect 11518 7032 11574 7041
rect 11428 6996 11480 7002
rect 11518 6967 11574 6976
rect 11428 6938 11480 6944
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11164 4486 11192 4626
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4078 11192 4422
rect 11348 4282 11376 5034
rect 11624 4554 11652 9166
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11072 3862 11192 3890
rect 10966 2952 11022 2961
rect 10966 2887 11022 2896
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10980 2038 11008 2887
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11072 2417 11100 2790
rect 11058 2408 11114 2417
rect 11058 2343 11114 2352
rect 10968 2032 11020 2038
rect 10968 1974 11020 1980
rect 11164 513 11192 3862
rect 11348 2990 11376 4218
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3505 11468 3878
rect 11426 3496 11482 3505
rect 11426 3431 11482 3440
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11428 2848 11480 2854
rect 11334 2816 11390 2825
rect 11428 2790 11480 2796
rect 11334 2751 11390 2760
rect 11150 504 11206 513
rect 2870 232 2926 241
rect 2870 167 2926 176
rect 3054 0 3110 480
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4710 0 4766 480
rect 5262 0 5318 480
rect 5814 0 5870 480
rect 6366 0 6422 480
rect 6918 0 6974 480
rect 7470 0 7526 480
rect 8022 0 8078 480
rect 8574 0 8630 480
rect 9126 0 9182 480
rect 9678 0 9734 480
rect 10230 0 10286 480
rect 10782 0 10838 480
rect 11348 480 11376 2751
rect 11440 1737 11468 2790
rect 11426 1728 11482 1737
rect 11426 1663 11482 1672
rect 11532 1329 11560 3334
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11518 1320 11574 1329
rect 11518 1255 11574 1264
rect 11624 921 11652 2246
rect 11716 1970 11744 8774
rect 11808 8129 11836 12310
rect 11794 8120 11850 8129
rect 11794 8055 11850 8064
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11808 7342 11836 7890
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11794 7168 11850 7177
rect 11794 7103 11850 7112
rect 11808 4010 11836 7103
rect 11900 5574 11928 15558
rect 11978 15464 12034 15473
rect 12084 15450 12112 15558
rect 12346 15520 12402 16000
rect 13174 15520 13230 16000
rect 13910 15520 13966 16000
rect 14738 15520 14794 16000
rect 15566 15520 15622 16000
rect 12360 15450 12388 15520
rect 12084 15422 12388 15450
rect 11978 15399 12034 15408
rect 11992 12374 12020 15399
rect 12898 13424 12954 13433
rect 12898 13359 12954 13368
rect 12449 13084 12745 13104
rect 12505 13082 12529 13084
rect 12585 13082 12609 13084
rect 12665 13082 12689 13084
rect 12527 13030 12529 13082
rect 12591 13030 12603 13082
rect 12665 13030 12667 13082
rect 12505 13028 12529 13030
rect 12585 13028 12609 13030
rect 12665 13028 12689 13030
rect 12449 13008 12745 13028
rect 12912 12753 12940 13359
rect 13188 13138 13216 15520
rect 13188 13110 13768 13138
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13084 12776 13136 12782
rect 12898 12744 12954 12753
rect 13084 12718 13136 12724
rect 12898 12679 12954 12688
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 11808 2802 11836 2858
rect 11992 2802 12020 12174
rect 12449 11996 12745 12016
rect 12505 11994 12529 11996
rect 12585 11994 12609 11996
rect 12665 11994 12689 11996
rect 12527 11942 12529 11994
rect 12591 11942 12603 11994
rect 12665 11942 12667 11994
rect 12505 11940 12529 11942
rect 12585 11940 12609 11942
rect 12665 11940 12689 11942
rect 12449 11920 12745 11940
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12084 10674 12112 11018
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12084 9450 12112 10610
rect 12268 10577 12296 11834
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12254 10568 12310 10577
rect 12254 10503 12310 10512
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12084 4593 12112 9386
rect 12070 4584 12126 4593
rect 12070 4519 12126 4528
rect 11808 2774 12020 2802
rect 11808 2292 11836 2774
rect 12176 2553 12204 9930
rect 12268 8945 12296 10202
rect 12254 8936 12310 8945
rect 12254 8871 12310 8880
rect 12268 5846 12296 8871
rect 12360 7449 12388 11018
rect 12449 10908 12745 10928
rect 12505 10906 12529 10908
rect 12585 10906 12609 10908
rect 12665 10906 12689 10908
rect 12527 10854 12529 10906
rect 12591 10854 12603 10906
rect 12665 10854 12667 10906
rect 12505 10852 12529 10854
rect 12585 10852 12609 10854
rect 12665 10852 12689 10854
rect 12449 10832 12745 10852
rect 12449 9820 12745 9840
rect 12505 9818 12529 9820
rect 12585 9818 12609 9820
rect 12665 9818 12689 9820
rect 12527 9766 12529 9818
rect 12591 9766 12603 9818
rect 12665 9766 12667 9818
rect 12505 9764 12529 9766
rect 12585 9764 12609 9766
rect 12665 9764 12689 9766
rect 12449 9744 12745 9764
rect 12820 9518 12848 11766
rect 12912 11694 12940 12679
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 9586 12940 11494
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9586 13032 9862
rect 13096 9722 13124 12718
rect 13556 12186 13584 12922
rect 13280 12158 13584 12186
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 9178 12756 9318
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 13004 9110 13032 9522
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12449 8732 12745 8752
rect 12505 8730 12529 8732
rect 12585 8730 12609 8732
rect 12665 8730 12689 8732
rect 12527 8678 12529 8730
rect 12591 8678 12603 8730
rect 12665 8678 12667 8730
rect 12505 8676 12529 8678
rect 12585 8676 12609 8678
rect 12665 8676 12689 8678
rect 12449 8656 12745 8676
rect 12820 8634 12848 8910
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 13004 8498 13032 9046
rect 13188 8537 13216 10406
rect 13280 9178 13308 12158
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13174 8528 13230 8537
rect 12992 8492 13044 8498
rect 13174 8463 13230 8472
rect 12992 8434 13044 8440
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12728 8242 12756 8298
rect 12728 8214 12848 8242
rect 12449 7644 12745 7664
rect 12505 7642 12529 7644
rect 12585 7642 12609 7644
rect 12665 7642 12689 7644
rect 12527 7590 12529 7642
rect 12591 7590 12603 7642
rect 12665 7590 12667 7642
rect 12505 7588 12529 7590
rect 12585 7588 12609 7590
rect 12665 7588 12689 7590
rect 12449 7568 12745 7588
rect 12820 7546 12848 8214
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12346 7440 12402 7449
rect 12346 7375 12402 7384
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12449 6556 12745 6576
rect 12505 6554 12529 6556
rect 12585 6554 12609 6556
rect 12665 6554 12689 6556
rect 12527 6502 12529 6554
rect 12591 6502 12603 6554
rect 12665 6502 12667 6554
rect 12505 6500 12529 6502
rect 12585 6500 12609 6502
rect 12665 6500 12689 6502
rect 12449 6480 12745 6500
rect 12820 5914 12848 7210
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6458 12940 7142
rect 13004 6934 13032 7686
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13096 7002 13124 7346
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 13004 6322 13032 6870
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12268 4185 12296 5646
rect 12449 5468 12745 5488
rect 12505 5466 12529 5468
rect 12585 5466 12609 5468
rect 12665 5466 12689 5468
rect 12527 5414 12529 5466
rect 12591 5414 12603 5466
rect 12665 5414 12667 5466
rect 12505 5412 12529 5414
rect 12585 5412 12609 5414
rect 12665 5412 12689 5414
rect 12449 5392 12745 5412
rect 12438 5264 12494 5273
rect 12438 5199 12494 5208
rect 12452 5166 12480 5199
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12544 4826 12572 4966
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12449 4380 12745 4400
rect 12505 4378 12529 4380
rect 12585 4378 12609 4380
rect 12665 4378 12689 4380
rect 12527 4326 12529 4378
rect 12591 4326 12603 4378
rect 12665 4326 12667 4378
rect 12505 4324 12529 4326
rect 12585 4324 12609 4326
rect 12665 4324 12689 4326
rect 12449 4304 12745 4324
rect 12440 4208 12492 4214
rect 12254 4176 12310 4185
rect 12440 4150 12492 4156
rect 12254 4111 12310 4120
rect 12162 2544 12218 2553
rect 12268 2514 12296 4111
rect 12346 3768 12402 3777
rect 12346 3703 12348 3712
rect 12400 3703 12402 3712
rect 12348 3674 12400 3680
rect 12452 3602 12480 4150
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12449 3292 12745 3312
rect 12505 3290 12529 3292
rect 12585 3290 12609 3292
rect 12665 3290 12689 3292
rect 12527 3238 12529 3290
rect 12591 3238 12603 3290
rect 12665 3238 12667 3290
rect 12505 3236 12529 3238
rect 12585 3236 12609 3238
rect 12665 3236 12689 3238
rect 12449 3216 12745 3236
rect 12912 2802 12940 6054
rect 13188 5710 13216 6258
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13188 5234 13216 5646
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 13004 3097 13032 4626
rect 12990 3088 13046 3097
rect 12990 3023 13046 3032
rect 13280 2990 13308 8978
rect 13372 6118 13400 9658
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13358 5128 13414 5137
rect 13358 5063 13414 5072
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 12820 2774 12940 2802
rect 12162 2479 12218 2488
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 11808 2264 11928 2292
rect 11704 1964 11756 1970
rect 11704 1906 11756 1912
rect 11610 912 11666 921
rect 11610 847 11666 856
rect 11900 480 11928 2264
rect 12449 2204 12745 2224
rect 12505 2202 12529 2204
rect 12585 2202 12609 2204
rect 12665 2202 12689 2204
rect 12527 2150 12529 2202
rect 12591 2150 12603 2202
rect 12665 2150 12667 2202
rect 12505 2148 12529 2150
rect 12585 2148 12609 2150
rect 12665 2148 12689 2150
rect 12449 2128 12745 2148
rect 12820 1442 12848 2774
rect 13372 2514 13400 5063
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13464 1698 13492 12038
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13556 10742 13584 11562
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13634 8256 13690 8265
rect 13634 8191 13690 8200
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 5817 13584 7686
rect 13648 7313 13676 8191
rect 13634 7304 13690 7313
rect 13634 7239 13690 7248
rect 13648 6186 13676 7239
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13542 5808 13598 5817
rect 13542 5743 13598 5752
rect 13542 5400 13598 5409
rect 13542 5335 13598 5344
rect 13556 4282 13584 5335
rect 13634 4992 13690 5001
rect 13634 4927 13690 4936
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13542 4176 13598 4185
rect 13542 4111 13598 4120
rect 13556 2650 13584 4111
rect 13648 3738 13676 4927
rect 13740 4690 13768 13110
rect 13924 12170 13952 15520
rect 14752 12442 14780 15520
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13726 4584 13782 4593
rect 13726 4519 13782 4528
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13740 3194 13768 4519
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 13832 2530 13860 9114
rect 13556 2502 13860 2530
rect 12992 1692 13044 1698
rect 12992 1634 13044 1640
rect 13452 1692 13504 1698
rect 13452 1634 13504 1640
rect 12452 1414 12848 1442
rect 12452 480 12480 1414
rect 12624 1352 12676 1358
rect 12624 1294 12676 1300
rect 11150 439 11206 448
rect 11334 0 11390 480
rect 11886 0 11942 480
rect 12438 0 12494 480
rect 12636 241 12664 1294
rect 13004 480 13032 1634
rect 13556 480 13584 2502
rect 14108 480 14136 12310
rect 15580 11626 15608 15520
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 14646 3632 14702 3641
rect 14646 3567 14702 3576
rect 14660 480 14688 3567
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 15212 480 15240 2518
rect 15764 480 15792 3062
rect 12622 232 12678 241
rect 12622 167 12678 176
rect 12990 0 13046 480
rect 13542 0 13598 480
rect 14094 0 14150 480
rect 14646 0 14702 480
rect 15198 0 15254 480
rect 15750 0 15806 480
<< via2 >>
rect 3330 15816 3386 15872
rect 1490 14592 1546 14648
rect 938 7928 994 7984
rect 846 6568 902 6624
rect 2594 15000 2650 15056
rect 1122 8200 1178 8256
rect 1490 7248 1546 7304
rect 1214 4528 1270 4584
rect 1030 3712 1086 3768
rect 1398 3032 1454 3088
rect 2134 12724 2136 12744
rect 2136 12724 2188 12744
rect 2188 12724 2190 12744
rect 2134 12688 2190 12724
rect 1766 9288 1822 9344
rect 1766 5888 1822 5944
rect 1674 5616 1730 5672
rect 1950 6024 2006 6080
rect 1950 5480 2006 5536
rect 1858 5344 1914 5400
rect 1674 3576 1730 3632
rect 1766 2624 1822 2680
rect 1582 1264 1638 1320
rect 2226 5072 2282 5128
rect 2134 3440 2190 3496
rect 2042 1672 2098 1728
rect 11610 15816 11666 15872
rect 4066 14204 4122 14240
rect 4066 14184 4068 14204
rect 4068 14184 4120 14204
rect 4120 14184 4122 14204
rect 4066 13812 4068 13832
rect 4068 13812 4120 13832
rect 4120 13812 4122 13832
rect 4066 13776 4122 13812
rect 3254 13082 3310 13084
rect 3334 13082 3390 13084
rect 3414 13082 3470 13084
rect 3494 13082 3550 13084
rect 3254 13030 3280 13082
rect 3280 13030 3310 13082
rect 3334 13030 3344 13082
rect 3344 13030 3390 13082
rect 3414 13030 3460 13082
rect 3460 13030 3470 13082
rect 3494 13030 3524 13082
rect 3524 13030 3550 13082
rect 3254 13028 3310 13030
rect 3334 13028 3390 13030
rect 3414 13028 3470 13030
rect 3494 13028 3550 13030
rect 3054 12960 3110 13016
rect 2686 11056 2742 11112
rect 2410 9968 2466 10024
rect 2686 9288 2742 9344
rect 3514 12588 3516 12608
rect 3516 12588 3568 12608
rect 3568 12588 3570 12608
rect 3514 12552 3570 12588
rect 3238 12436 3294 12472
rect 3238 12416 3240 12436
rect 3240 12416 3292 12436
rect 3292 12416 3294 12436
rect 3254 11994 3310 11996
rect 3334 11994 3390 11996
rect 3414 11994 3470 11996
rect 3494 11994 3550 11996
rect 3254 11942 3280 11994
rect 3280 11942 3310 11994
rect 3334 11942 3344 11994
rect 3344 11942 3390 11994
rect 3414 11942 3460 11994
rect 3460 11942 3470 11994
rect 3494 11942 3524 11994
rect 3524 11942 3550 11994
rect 3254 11940 3310 11942
rect 3334 11940 3390 11942
rect 3414 11940 3470 11942
rect 3494 11940 3550 11942
rect 3882 13368 3938 13424
rect 3054 10920 3110 10976
rect 2962 10240 3018 10296
rect 2778 9036 2834 9072
rect 2778 9016 2780 9036
rect 2780 9016 2832 9036
rect 2832 9016 2834 9036
rect 2594 4800 2650 4856
rect 2502 4664 2558 4720
rect 2318 856 2374 912
rect 3254 10906 3310 10908
rect 3334 10906 3390 10908
rect 3414 10906 3470 10908
rect 3494 10906 3550 10908
rect 3254 10854 3280 10906
rect 3280 10854 3310 10906
rect 3334 10854 3344 10906
rect 3344 10854 3390 10906
rect 3414 10854 3460 10906
rect 3460 10854 3470 10906
rect 3494 10854 3524 10906
rect 3524 10854 3550 10906
rect 3254 10852 3310 10854
rect 3334 10852 3390 10854
rect 3414 10852 3470 10854
rect 3494 10852 3550 10854
rect 3146 9968 3202 10024
rect 3254 9818 3310 9820
rect 3334 9818 3390 9820
rect 3414 9818 3470 9820
rect 3494 9818 3550 9820
rect 3254 9766 3280 9818
rect 3280 9766 3310 9818
rect 3334 9766 3344 9818
rect 3344 9766 3390 9818
rect 3414 9766 3460 9818
rect 3460 9766 3470 9818
rect 3494 9766 3524 9818
rect 3524 9766 3550 9818
rect 3254 9764 3310 9766
rect 3334 9764 3390 9766
rect 3414 9764 3470 9766
rect 3494 9764 3550 9766
rect 3606 9288 3662 9344
rect 3254 8730 3310 8732
rect 3334 8730 3390 8732
rect 3414 8730 3470 8732
rect 3494 8730 3550 8732
rect 3254 8678 3280 8730
rect 3280 8678 3310 8730
rect 3334 8678 3344 8730
rect 3344 8678 3390 8730
rect 3414 8678 3460 8730
rect 3460 8678 3470 8730
rect 3494 8678 3524 8730
rect 3524 8678 3550 8730
rect 3254 8676 3310 8678
rect 3334 8676 3390 8678
rect 3414 8676 3470 8678
rect 3494 8676 3550 8678
rect 3254 7642 3310 7644
rect 3334 7642 3390 7644
rect 3414 7642 3470 7644
rect 3494 7642 3550 7644
rect 3254 7590 3280 7642
rect 3280 7590 3310 7642
rect 3334 7590 3344 7642
rect 3344 7590 3390 7642
rect 3414 7590 3460 7642
rect 3460 7590 3470 7642
rect 3494 7590 3524 7642
rect 3524 7590 3550 7642
rect 3254 7588 3310 7590
rect 3334 7588 3390 7590
rect 3414 7588 3470 7590
rect 3494 7588 3550 7590
rect 3422 7384 3478 7440
rect 3254 6554 3310 6556
rect 3334 6554 3390 6556
rect 3414 6554 3470 6556
rect 3494 6554 3550 6556
rect 3254 6502 3280 6554
rect 3280 6502 3310 6554
rect 3334 6502 3344 6554
rect 3344 6502 3390 6554
rect 3414 6502 3460 6554
rect 3460 6502 3470 6554
rect 3494 6502 3524 6554
rect 3524 6502 3550 6554
rect 3254 6500 3310 6502
rect 3334 6500 3390 6502
rect 3414 6500 3470 6502
rect 3494 6500 3550 6502
rect 3254 5466 3310 5468
rect 3334 5466 3390 5468
rect 3414 5466 3470 5468
rect 3494 5466 3550 5468
rect 3254 5414 3280 5466
rect 3280 5414 3310 5466
rect 3334 5414 3344 5466
rect 3344 5414 3390 5466
rect 3414 5414 3460 5466
rect 3460 5414 3470 5466
rect 3494 5414 3524 5466
rect 3524 5414 3550 5466
rect 3254 5412 3310 5414
rect 3334 5412 3390 5414
rect 3414 5412 3470 5414
rect 3494 5412 3550 5414
rect 3514 5228 3570 5264
rect 3514 5208 3516 5228
rect 3516 5208 3568 5228
rect 3568 5208 3570 5228
rect 3146 4528 3202 4584
rect 2962 2488 3018 2544
rect 3254 4378 3310 4380
rect 3334 4378 3390 4380
rect 3414 4378 3470 4380
rect 3494 4378 3550 4380
rect 3254 4326 3280 4378
rect 3280 4326 3310 4378
rect 3334 4326 3344 4378
rect 3344 4326 3390 4378
rect 3414 4326 3460 4378
rect 3460 4326 3470 4378
rect 3494 4326 3524 4378
rect 3524 4326 3550 4378
rect 3254 4324 3310 4326
rect 3334 4324 3390 4326
rect 3414 4324 3470 4326
rect 3494 4324 3550 4326
rect 3882 11192 3938 11248
rect 3974 10956 3976 10976
rect 3976 10956 4028 10976
rect 4028 10956 4030 10976
rect 3974 10920 4030 10956
rect 3974 10104 4030 10160
rect 4250 12300 4306 12336
rect 4250 12280 4252 12300
rect 4252 12280 4304 12300
rect 4304 12280 4306 12300
rect 3974 7792 4030 7848
rect 3974 7112 4030 7168
rect 4066 6432 4122 6488
rect 4066 6160 4122 6216
rect 4710 12144 4766 12200
rect 4066 5752 4122 5808
rect 4066 4936 4122 4992
rect 3882 4392 3938 4448
rect 3606 4120 3662 4176
rect 3790 3884 3792 3904
rect 3792 3884 3844 3904
rect 3844 3884 3846 3904
rect 3790 3848 3846 3884
rect 3974 3848 4030 3904
rect 3974 3712 4030 3768
rect 3254 3290 3310 3292
rect 3334 3290 3390 3292
rect 3414 3290 3470 3292
rect 3494 3290 3550 3292
rect 3254 3238 3280 3290
rect 3280 3238 3310 3290
rect 3334 3238 3344 3290
rect 3344 3238 3390 3290
rect 3414 3238 3460 3290
rect 3460 3238 3470 3290
rect 3494 3238 3524 3290
rect 3524 3238 3550 3290
rect 3254 3236 3310 3238
rect 3334 3236 3390 3238
rect 3414 3236 3470 3238
rect 3494 3236 3550 3238
rect 4066 2896 4122 2952
rect 4342 4256 4398 4312
rect 4526 3168 4582 3224
rect 3698 2488 3754 2544
rect 2870 2352 2926 2408
rect 4618 2488 4674 2544
rect 3254 2202 3310 2204
rect 3334 2202 3390 2204
rect 3414 2202 3470 2204
rect 3494 2202 3550 2204
rect 3254 2150 3280 2202
rect 3280 2150 3310 2202
rect 3334 2150 3344 2202
rect 3344 2150 3390 2202
rect 3414 2150 3460 2202
rect 3460 2150 3470 2202
rect 3494 2150 3524 2202
rect 3524 2150 3550 2202
rect 3254 2148 3310 2150
rect 3334 2148 3390 2150
rect 3414 2148 3470 2150
rect 3494 2148 3550 2150
rect 3054 2080 3110 2136
rect 4618 2388 4620 2408
rect 4620 2388 4672 2408
rect 4672 2388 4674 2408
rect 4618 2352 4674 2388
rect 2778 448 2834 504
rect 4802 6432 4858 6488
rect 4894 2796 4896 2816
rect 4896 2796 4948 2816
rect 4948 2796 4950 2816
rect 4894 2760 4950 2796
rect 5170 12144 5226 12200
rect 5078 11756 5134 11792
rect 5078 11736 5080 11756
rect 5080 11736 5132 11756
rect 5132 11736 5134 11756
rect 5078 8880 5134 8936
rect 5078 8472 5134 8528
rect 5078 6704 5134 6760
rect 5553 13626 5609 13628
rect 5633 13626 5689 13628
rect 5713 13626 5769 13628
rect 5793 13626 5849 13628
rect 5553 13574 5579 13626
rect 5579 13574 5609 13626
rect 5633 13574 5643 13626
rect 5643 13574 5689 13626
rect 5713 13574 5759 13626
rect 5759 13574 5769 13626
rect 5793 13574 5823 13626
rect 5823 13574 5849 13626
rect 5553 13572 5609 13574
rect 5633 13572 5689 13574
rect 5713 13572 5769 13574
rect 5793 13572 5849 13574
rect 5553 12538 5609 12540
rect 5633 12538 5689 12540
rect 5713 12538 5769 12540
rect 5793 12538 5849 12540
rect 5553 12486 5579 12538
rect 5579 12486 5609 12538
rect 5633 12486 5643 12538
rect 5643 12486 5689 12538
rect 5713 12486 5759 12538
rect 5759 12486 5769 12538
rect 5793 12486 5823 12538
rect 5823 12486 5849 12538
rect 5553 12484 5609 12486
rect 5633 12484 5689 12486
rect 5713 12484 5769 12486
rect 5793 12484 5849 12486
rect 6458 15408 6514 15464
rect 5553 11450 5609 11452
rect 5633 11450 5689 11452
rect 5713 11450 5769 11452
rect 5793 11450 5849 11452
rect 5553 11398 5579 11450
rect 5579 11398 5609 11450
rect 5633 11398 5643 11450
rect 5643 11398 5689 11450
rect 5713 11398 5759 11450
rect 5759 11398 5769 11450
rect 5793 11398 5823 11450
rect 5823 11398 5849 11450
rect 5553 11396 5609 11398
rect 5633 11396 5689 11398
rect 5713 11396 5769 11398
rect 5793 11396 5849 11398
rect 6090 12280 6146 12336
rect 6458 11192 6514 11248
rect 5553 10362 5609 10364
rect 5633 10362 5689 10364
rect 5713 10362 5769 10364
rect 5793 10362 5849 10364
rect 5553 10310 5579 10362
rect 5579 10310 5609 10362
rect 5633 10310 5643 10362
rect 5643 10310 5689 10362
rect 5713 10310 5759 10362
rect 5759 10310 5769 10362
rect 5793 10310 5823 10362
rect 5823 10310 5849 10362
rect 5553 10308 5609 10310
rect 5633 10308 5689 10310
rect 5713 10308 5769 10310
rect 5793 10308 5849 10310
rect 5553 9274 5609 9276
rect 5633 9274 5689 9276
rect 5713 9274 5769 9276
rect 5793 9274 5849 9276
rect 5553 9222 5579 9274
rect 5579 9222 5609 9274
rect 5633 9222 5643 9274
rect 5643 9222 5689 9274
rect 5713 9222 5759 9274
rect 5759 9222 5769 9274
rect 5793 9222 5823 9274
rect 5823 9222 5849 9274
rect 5553 9220 5609 9222
rect 5633 9220 5689 9222
rect 5713 9220 5769 9222
rect 5793 9220 5849 9222
rect 5553 8186 5609 8188
rect 5633 8186 5689 8188
rect 5713 8186 5769 8188
rect 5793 8186 5849 8188
rect 5553 8134 5579 8186
rect 5579 8134 5609 8186
rect 5633 8134 5643 8186
rect 5643 8134 5689 8186
rect 5713 8134 5759 8186
rect 5759 8134 5769 8186
rect 5793 8134 5823 8186
rect 5823 8134 5849 8186
rect 5553 8132 5609 8134
rect 5633 8132 5689 8134
rect 5713 8132 5769 8134
rect 5793 8132 5849 8134
rect 5354 5752 5410 5808
rect 5262 4800 5318 4856
rect 5078 3032 5134 3088
rect 5262 4020 5264 4040
rect 5264 4020 5316 4040
rect 5316 4020 5318 4040
rect 5262 3984 5318 4020
rect 5553 7098 5609 7100
rect 5633 7098 5689 7100
rect 5713 7098 5769 7100
rect 5793 7098 5849 7100
rect 5553 7046 5579 7098
rect 5579 7046 5609 7098
rect 5633 7046 5643 7098
rect 5643 7046 5689 7098
rect 5713 7046 5759 7098
rect 5759 7046 5769 7098
rect 5793 7046 5823 7098
rect 5823 7046 5849 7098
rect 5553 7044 5609 7046
rect 5633 7044 5689 7046
rect 5713 7044 5769 7046
rect 5793 7044 5849 7046
rect 5553 6010 5609 6012
rect 5633 6010 5689 6012
rect 5713 6010 5769 6012
rect 5793 6010 5849 6012
rect 5553 5958 5579 6010
rect 5579 5958 5609 6010
rect 5633 5958 5643 6010
rect 5643 5958 5689 6010
rect 5713 5958 5759 6010
rect 5759 5958 5769 6010
rect 5793 5958 5823 6010
rect 5823 5958 5849 6010
rect 5553 5956 5609 5958
rect 5633 5956 5689 5958
rect 5713 5956 5769 5958
rect 5793 5956 5849 5958
rect 5553 4922 5609 4924
rect 5633 4922 5689 4924
rect 5713 4922 5769 4924
rect 5793 4922 5849 4924
rect 5553 4870 5579 4922
rect 5579 4870 5609 4922
rect 5633 4870 5643 4922
rect 5643 4870 5689 4922
rect 5713 4870 5759 4922
rect 5759 4870 5769 4922
rect 5793 4870 5823 4922
rect 5823 4870 5849 4922
rect 5553 4868 5609 4870
rect 5633 4868 5689 4870
rect 5713 4868 5769 4870
rect 5793 4868 5849 4870
rect 6090 5888 6146 5944
rect 5814 4564 5816 4584
rect 5816 4564 5868 4584
rect 5868 4564 5870 4584
rect 5814 4528 5870 4564
rect 5553 3834 5609 3836
rect 5633 3834 5689 3836
rect 5713 3834 5769 3836
rect 5793 3834 5849 3836
rect 5553 3782 5579 3834
rect 5579 3782 5609 3834
rect 5633 3782 5643 3834
rect 5643 3782 5689 3834
rect 5713 3782 5759 3834
rect 5759 3782 5769 3834
rect 5793 3782 5823 3834
rect 5823 3782 5849 3834
rect 5553 3780 5609 3782
rect 5633 3780 5689 3782
rect 5713 3780 5769 3782
rect 5793 3780 5849 3782
rect 5446 3440 5502 3496
rect 5553 2746 5609 2748
rect 5633 2746 5689 2748
rect 5713 2746 5769 2748
rect 5793 2746 5849 2748
rect 5553 2694 5579 2746
rect 5579 2694 5609 2746
rect 5633 2694 5643 2746
rect 5643 2694 5689 2746
rect 5713 2694 5759 2746
rect 5759 2694 5769 2746
rect 5793 2694 5823 2746
rect 5823 2694 5849 2746
rect 5553 2692 5609 2694
rect 5633 2692 5689 2694
rect 5713 2692 5769 2694
rect 5793 2692 5849 2694
rect 6274 5888 6330 5944
rect 6550 6296 6606 6352
rect 6458 5344 6514 5400
rect 7194 12688 7250 12744
rect 7102 10512 7158 10568
rect 7010 10240 7066 10296
rect 6734 4664 6790 4720
rect 7194 9424 7250 9480
rect 7562 9560 7618 9616
rect 7470 9424 7526 9480
rect 7470 9288 7526 9344
rect 7286 5616 7342 5672
rect 7286 5092 7342 5128
rect 7286 5072 7288 5092
rect 7288 5072 7340 5092
rect 7340 5072 7342 5092
rect 7852 13082 7908 13084
rect 7932 13082 7988 13084
rect 8012 13082 8068 13084
rect 8092 13082 8148 13084
rect 7852 13030 7878 13082
rect 7878 13030 7908 13082
rect 7932 13030 7942 13082
rect 7942 13030 7988 13082
rect 8012 13030 8058 13082
rect 8058 13030 8068 13082
rect 8092 13030 8122 13082
rect 8122 13030 8148 13082
rect 7852 13028 7908 13030
rect 7932 13028 7988 13030
rect 8012 13028 8068 13030
rect 8092 13028 8148 13030
rect 7852 11994 7908 11996
rect 7932 11994 7988 11996
rect 8012 11994 8068 11996
rect 8092 11994 8148 11996
rect 7852 11942 7878 11994
rect 7878 11942 7908 11994
rect 7932 11942 7942 11994
rect 7942 11942 7988 11994
rect 8012 11942 8058 11994
rect 8058 11942 8068 11994
rect 8092 11942 8122 11994
rect 8122 11942 8148 11994
rect 7852 11940 7908 11942
rect 7932 11940 7988 11942
rect 8012 11940 8068 11942
rect 8092 11940 8148 11942
rect 7852 10906 7908 10908
rect 7932 10906 7988 10908
rect 8012 10906 8068 10908
rect 8092 10906 8148 10908
rect 7852 10854 7878 10906
rect 7878 10854 7908 10906
rect 7932 10854 7942 10906
rect 7942 10854 7988 10906
rect 8012 10854 8058 10906
rect 8058 10854 8068 10906
rect 8092 10854 8122 10906
rect 8122 10854 8148 10906
rect 7852 10852 7908 10854
rect 7932 10852 7988 10854
rect 8012 10852 8068 10854
rect 8092 10852 8148 10854
rect 8206 10512 8262 10568
rect 8482 12280 8538 12336
rect 8942 12688 8998 12744
rect 7852 9818 7908 9820
rect 7932 9818 7988 9820
rect 8012 9818 8068 9820
rect 8092 9818 8148 9820
rect 7852 9766 7878 9818
rect 7878 9766 7908 9818
rect 7932 9766 7942 9818
rect 7942 9766 7988 9818
rect 8012 9766 8058 9818
rect 8058 9766 8068 9818
rect 8092 9766 8122 9818
rect 8122 9766 8148 9818
rect 7852 9764 7908 9766
rect 7932 9764 7988 9766
rect 8012 9764 8068 9766
rect 8092 9764 8148 9766
rect 7852 8730 7908 8732
rect 7932 8730 7988 8732
rect 8012 8730 8068 8732
rect 8092 8730 8148 8732
rect 7852 8678 7878 8730
rect 7878 8678 7908 8730
rect 7932 8678 7942 8730
rect 7942 8678 7988 8730
rect 8012 8678 8058 8730
rect 8058 8678 8068 8730
rect 8092 8678 8122 8730
rect 8122 8678 8148 8730
rect 7852 8676 7908 8678
rect 7932 8676 7988 8678
rect 8012 8676 8068 8678
rect 8092 8676 8148 8678
rect 7852 7642 7908 7644
rect 7932 7642 7988 7644
rect 8012 7642 8068 7644
rect 8092 7642 8148 7644
rect 7852 7590 7878 7642
rect 7878 7590 7908 7642
rect 7932 7590 7942 7642
rect 7942 7590 7988 7642
rect 8012 7590 8058 7642
rect 8058 7590 8068 7642
rect 8092 7590 8122 7642
rect 8122 7590 8148 7642
rect 7852 7588 7908 7590
rect 7932 7588 7988 7590
rect 8012 7588 8068 7590
rect 8092 7588 8148 7590
rect 7852 6554 7908 6556
rect 7932 6554 7988 6556
rect 8012 6554 8068 6556
rect 8092 6554 8148 6556
rect 7852 6502 7878 6554
rect 7878 6502 7908 6554
rect 7932 6502 7942 6554
rect 7942 6502 7988 6554
rect 8012 6502 8058 6554
rect 8058 6502 8068 6554
rect 8092 6502 8122 6554
rect 8122 6502 8148 6554
rect 7852 6500 7908 6502
rect 7932 6500 7988 6502
rect 8012 6500 8068 6502
rect 8092 6500 8148 6502
rect 7852 5466 7908 5468
rect 7932 5466 7988 5468
rect 8012 5466 8068 5468
rect 8092 5466 8148 5468
rect 7852 5414 7878 5466
rect 7878 5414 7908 5466
rect 7932 5414 7942 5466
rect 7942 5414 7988 5466
rect 8012 5414 8058 5466
rect 8058 5414 8068 5466
rect 8092 5414 8122 5466
rect 8122 5414 8148 5466
rect 7852 5412 7908 5414
rect 7932 5412 7988 5414
rect 8012 5412 8068 5414
rect 8092 5412 8148 5414
rect 7746 5072 7802 5128
rect 7852 4378 7908 4380
rect 7932 4378 7988 4380
rect 8012 4378 8068 4380
rect 8092 4378 8148 4380
rect 7852 4326 7878 4378
rect 7878 4326 7908 4378
rect 7932 4326 7942 4378
rect 7942 4326 7988 4378
rect 8012 4326 8058 4378
rect 8058 4326 8068 4378
rect 8092 4326 8122 4378
rect 8122 4326 8148 4378
rect 7852 4324 7908 4326
rect 7932 4324 7988 4326
rect 8012 4324 8068 4326
rect 8092 4324 8148 4326
rect 8574 9016 8630 9072
rect 8666 7928 8722 7984
rect 8666 6296 8722 6352
rect 8666 6024 8722 6080
rect 8666 4664 8722 4720
rect 7852 3290 7908 3292
rect 7932 3290 7988 3292
rect 8012 3290 8068 3292
rect 8092 3290 8148 3292
rect 7852 3238 7878 3290
rect 7878 3238 7908 3290
rect 7932 3238 7942 3290
rect 7942 3238 7988 3290
rect 8012 3238 8058 3290
rect 8058 3238 8068 3290
rect 8092 3238 8122 3290
rect 8122 3238 8148 3290
rect 7852 3236 7908 3238
rect 7932 3236 7988 3238
rect 8012 3236 8068 3238
rect 8092 3236 8148 3238
rect 7852 2202 7908 2204
rect 7932 2202 7988 2204
rect 8012 2202 8068 2204
rect 8092 2202 8148 2204
rect 7852 2150 7878 2202
rect 7878 2150 7908 2202
rect 7932 2150 7942 2202
rect 7942 2150 7988 2202
rect 8012 2150 8058 2202
rect 8058 2150 8068 2202
rect 8092 2150 8122 2202
rect 8122 2150 8148 2202
rect 7852 2148 7908 2150
rect 7932 2148 7988 2150
rect 8012 2148 8068 2150
rect 8092 2148 8148 2150
rect 8758 2896 8814 2952
rect 9770 12824 9826 12880
rect 9862 12708 9918 12744
rect 9862 12688 9864 12708
rect 9864 12688 9916 12708
rect 9916 12688 9918 12708
rect 9678 12008 9734 12064
rect 9126 10260 9182 10296
rect 9126 10240 9128 10260
rect 9128 10240 9180 10260
rect 9180 10240 9182 10260
rect 9310 9968 9366 10024
rect 9126 7248 9182 7304
rect 8942 6740 8944 6760
rect 8944 6740 8996 6760
rect 8996 6740 8998 6760
rect 8942 6704 8998 6740
rect 9034 5208 9090 5264
rect 8942 3440 8998 3496
rect 10690 13776 10746 13832
rect 10150 13626 10206 13628
rect 10230 13626 10286 13628
rect 10310 13626 10366 13628
rect 10390 13626 10446 13628
rect 10150 13574 10176 13626
rect 10176 13574 10206 13626
rect 10230 13574 10240 13626
rect 10240 13574 10286 13626
rect 10310 13574 10356 13626
rect 10356 13574 10366 13626
rect 10390 13574 10420 13626
rect 10420 13574 10446 13626
rect 10150 13572 10206 13574
rect 10230 13572 10286 13574
rect 10310 13572 10366 13574
rect 10390 13572 10446 13574
rect 10150 12538 10206 12540
rect 10230 12538 10286 12540
rect 10310 12538 10366 12540
rect 10390 12538 10446 12540
rect 10150 12486 10176 12538
rect 10176 12486 10206 12538
rect 10230 12486 10240 12538
rect 10240 12486 10286 12538
rect 10310 12486 10356 12538
rect 10356 12486 10366 12538
rect 10390 12486 10420 12538
rect 10420 12486 10446 12538
rect 10150 12484 10206 12486
rect 10230 12484 10286 12486
rect 10310 12484 10366 12486
rect 10390 12484 10446 12486
rect 10150 11450 10206 11452
rect 10230 11450 10286 11452
rect 10310 11450 10366 11452
rect 10390 11450 10446 11452
rect 10150 11398 10176 11450
rect 10176 11398 10206 11450
rect 10230 11398 10240 11450
rect 10240 11398 10286 11450
rect 10310 11398 10356 11450
rect 10356 11398 10366 11450
rect 10390 11398 10420 11450
rect 10420 11398 10446 11450
rect 10150 11396 10206 11398
rect 10230 11396 10286 11398
rect 10310 11396 10366 11398
rect 10390 11396 10446 11398
rect 9586 5888 9642 5944
rect 9586 5752 9642 5808
rect 9678 3712 9734 3768
rect 10150 10362 10206 10364
rect 10230 10362 10286 10364
rect 10310 10362 10366 10364
rect 10390 10362 10446 10364
rect 10150 10310 10176 10362
rect 10176 10310 10206 10362
rect 10230 10310 10240 10362
rect 10240 10310 10286 10362
rect 10310 10310 10356 10362
rect 10356 10310 10366 10362
rect 10390 10310 10420 10362
rect 10420 10310 10446 10362
rect 10150 10308 10206 10310
rect 10230 10308 10286 10310
rect 10310 10308 10366 10310
rect 10390 10308 10446 10310
rect 10046 10140 10048 10160
rect 10048 10140 10100 10160
rect 10100 10140 10102 10160
rect 10046 10104 10102 10140
rect 10046 9696 10102 9752
rect 10150 9274 10206 9276
rect 10230 9274 10286 9276
rect 10310 9274 10366 9276
rect 10390 9274 10446 9276
rect 10150 9222 10176 9274
rect 10176 9222 10206 9274
rect 10230 9222 10240 9274
rect 10240 9222 10286 9274
rect 10310 9222 10356 9274
rect 10356 9222 10366 9274
rect 10390 9222 10420 9274
rect 10420 9222 10446 9274
rect 10150 9220 10206 9222
rect 10230 9220 10286 9222
rect 10310 9220 10366 9222
rect 10390 9220 10446 9222
rect 10150 8186 10206 8188
rect 10230 8186 10286 8188
rect 10310 8186 10366 8188
rect 10390 8186 10446 8188
rect 10150 8134 10176 8186
rect 10176 8134 10206 8186
rect 10230 8134 10240 8186
rect 10240 8134 10286 8186
rect 10310 8134 10356 8186
rect 10356 8134 10366 8186
rect 10390 8134 10420 8186
rect 10420 8134 10446 8186
rect 10150 8132 10206 8134
rect 10230 8132 10286 8134
rect 10310 8132 10366 8134
rect 10390 8132 10446 8134
rect 10690 12144 10746 12200
rect 11058 15000 11114 15056
rect 11242 14592 11298 14648
rect 11150 14184 11206 14240
rect 11242 12824 11298 12880
rect 11058 12552 11114 12608
rect 11058 12144 11114 12200
rect 10966 12008 11022 12064
rect 11058 11756 11114 11792
rect 11058 11736 11060 11756
rect 11060 11736 11112 11756
rect 11112 11736 11114 11756
rect 11242 12280 11298 12336
rect 11058 11328 11114 11384
rect 10150 7098 10206 7100
rect 10230 7098 10286 7100
rect 10310 7098 10366 7100
rect 10390 7098 10446 7100
rect 10150 7046 10176 7098
rect 10176 7046 10206 7098
rect 10230 7046 10240 7098
rect 10240 7046 10286 7098
rect 10310 7046 10356 7098
rect 10356 7046 10366 7098
rect 10390 7046 10420 7098
rect 10420 7046 10446 7098
rect 10150 7044 10206 7046
rect 10230 7044 10286 7046
rect 10310 7044 10366 7046
rect 10390 7044 10446 7046
rect 10150 6010 10206 6012
rect 10230 6010 10286 6012
rect 10310 6010 10366 6012
rect 10390 6010 10446 6012
rect 10150 5958 10176 6010
rect 10176 5958 10206 6010
rect 10230 5958 10240 6010
rect 10240 5958 10286 6010
rect 10310 5958 10356 6010
rect 10356 5958 10366 6010
rect 10390 5958 10420 6010
rect 10420 5958 10446 6010
rect 10150 5956 10206 5958
rect 10230 5956 10286 5958
rect 10310 5956 10366 5958
rect 10390 5956 10446 5958
rect 10138 5208 10194 5264
rect 10230 5072 10286 5128
rect 10150 4922 10206 4924
rect 10230 4922 10286 4924
rect 10310 4922 10366 4924
rect 10390 4922 10446 4924
rect 10150 4870 10176 4922
rect 10176 4870 10206 4922
rect 10230 4870 10240 4922
rect 10240 4870 10286 4922
rect 10310 4870 10356 4922
rect 10356 4870 10366 4922
rect 10390 4870 10420 4922
rect 10420 4870 10446 4922
rect 10150 4868 10206 4870
rect 10230 4868 10286 4870
rect 10310 4868 10366 4870
rect 10390 4868 10446 4870
rect 10150 3834 10206 3836
rect 10230 3834 10286 3836
rect 10310 3834 10366 3836
rect 10390 3834 10446 3836
rect 10150 3782 10176 3834
rect 10176 3782 10206 3834
rect 10230 3782 10240 3834
rect 10240 3782 10286 3834
rect 10310 3782 10356 3834
rect 10356 3782 10366 3834
rect 10390 3782 10420 3834
rect 10420 3782 10446 3834
rect 10150 3780 10206 3782
rect 10230 3780 10286 3782
rect 10310 3780 10366 3782
rect 10390 3780 10446 3782
rect 9678 2896 9734 2952
rect 11058 10668 11114 10704
rect 11058 10648 11060 10668
rect 11060 10648 11112 10668
rect 11112 10648 11114 10668
rect 10966 9696 11022 9752
rect 11058 9288 11114 9344
rect 11702 9968 11758 10024
rect 11334 8608 11390 8664
rect 11426 8472 11482 8528
rect 11058 7792 11114 7848
rect 11058 7248 11114 7304
rect 11058 6840 11114 6896
rect 10874 6160 10930 6216
rect 10150 2746 10206 2748
rect 10230 2746 10286 2748
rect 10310 2746 10366 2748
rect 10390 2746 10446 2748
rect 10150 2694 10176 2746
rect 10176 2694 10206 2746
rect 10230 2694 10240 2746
rect 10240 2694 10286 2746
rect 10310 2694 10356 2746
rect 10356 2694 10366 2746
rect 10390 2694 10420 2746
rect 10420 2694 10446 2746
rect 10150 2692 10206 2694
rect 10230 2692 10286 2694
rect 10310 2692 10366 2694
rect 10390 2692 10446 2694
rect 11518 6976 11574 7032
rect 10966 2896 11022 2952
rect 11058 2352 11114 2408
rect 11426 3440 11482 3496
rect 11334 2760 11390 2816
rect 2870 176 2926 232
rect 11150 448 11206 504
rect 11426 1672 11482 1728
rect 11518 1264 11574 1320
rect 11794 8064 11850 8120
rect 11794 7112 11850 7168
rect 11978 15408 12034 15464
rect 12898 13368 12954 13424
rect 12449 13082 12505 13084
rect 12529 13082 12585 13084
rect 12609 13082 12665 13084
rect 12689 13082 12745 13084
rect 12449 13030 12475 13082
rect 12475 13030 12505 13082
rect 12529 13030 12539 13082
rect 12539 13030 12585 13082
rect 12609 13030 12655 13082
rect 12655 13030 12665 13082
rect 12689 13030 12719 13082
rect 12719 13030 12745 13082
rect 12449 13028 12505 13030
rect 12529 13028 12585 13030
rect 12609 13028 12665 13030
rect 12689 13028 12745 13030
rect 12898 12688 12954 12744
rect 12449 11994 12505 11996
rect 12529 11994 12585 11996
rect 12609 11994 12665 11996
rect 12689 11994 12745 11996
rect 12449 11942 12475 11994
rect 12475 11942 12505 11994
rect 12529 11942 12539 11994
rect 12539 11942 12585 11994
rect 12609 11942 12655 11994
rect 12655 11942 12665 11994
rect 12689 11942 12719 11994
rect 12719 11942 12745 11994
rect 12449 11940 12505 11942
rect 12529 11940 12585 11942
rect 12609 11940 12665 11942
rect 12689 11940 12745 11942
rect 12254 10512 12310 10568
rect 12070 4528 12126 4584
rect 12254 8880 12310 8936
rect 12449 10906 12505 10908
rect 12529 10906 12585 10908
rect 12609 10906 12665 10908
rect 12689 10906 12745 10908
rect 12449 10854 12475 10906
rect 12475 10854 12505 10906
rect 12529 10854 12539 10906
rect 12539 10854 12585 10906
rect 12609 10854 12655 10906
rect 12655 10854 12665 10906
rect 12689 10854 12719 10906
rect 12719 10854 12745 10906
rect 12449 10852 12505 10854
rect 12529 10852 12585 10854
rect 12609 10852 12665 10854
rect 12689 10852 12745 10854
rect 12449 9818 12505 9820
rect 12529 9818 12585 9820
rect 12609 9818 12665 9820
rect 12689 9818 12745 9820
rect 12449 9766 12475 9818
rect 12475 9766 12505 9818
rect 12529 9766 12539 9818
rect 12539 9766 12585 9818
rect 12609 9766 12655 9818
rect 12655 9766 12665 9818
rect 12689 9766 12719 9818
rect 12719 9766 12745 9818
rect 12449 9764 12505 9766
rect 12529 9764 12585 9766
rect 12609 9764 12665 9766
rect 12689 9764 12745 9766
rect 12449 8730 12505 8732
rect 12529 8730 12585 8732
rect 12609 8730 12665 8732
rect 12689 8730 12745 8732
rect 12449 8678 12475 8730
rect 12475 8678 12505 8730
rect 12529 8678 12539 8730
rect 12539 8678 12585 8730
rect 12609 8678 12655 8730
rect 12655 8678 12665 8730
rect 12689 8678 12719 8730
rect 12719 8678 12745 8730
rect 12449 8676 12505 8678
rect 12529 8676 12585 8678
rect 12609 8676 12665 8678
rect 12689 8676 12745 8678
rect 13174 8472 13230 8528
rect 12449 7642 12505 7644
rect 12529 7642 12585 7644
rect 12609 7642 12665 7644
rect 12689 7642 12745 7644
rect 12449 7590 12475 7642
rect 12475 7590 12505 7642
rect 12529 7590 12539 7642
rect 12539 7590 12585 7642
rect 12609 7590 12655 7642
rect 12655 7590 12665 7642
rect 12689 7590 12719 7642
rect 12719 7590 12745 7642
rect 12449 7588 12505 7590
rect 12529 7588 12585 7590
rect 12609 7588 12665 7590
rect 12689 7588 12745 7590
rect 12346 7384 12402 7440
rect 12449 6554 12505 6556
rect 12529 6554 12585 6556
rect 12609 6554 12665 6556
rect 12689 6554 12745 6556
rect 12449 6502 12475 6554
rect 12475 6502 12505 6554
rect 12529 6502 12539 6554
rect 12539 6502 12585 6554
rect 12609 6502 12655 6554
rect 12655 6502 12665 6554
rect 12689 6502 12719 6554
rect 12719 6502 12745 6554
rect 12449 6500 12505 6502
rect 12529 6500 12585 6502
rect 12609 6500 12665 6502
rect 12689 6500 12745 6502
rect 12449 5466 12505 5468
rect 12529 5466 12585 5468
rect 12609 5466 12665 5468
rect 12689 5466 12745 5468
rect 12449 5414 12475 5466
rect 12475 5414 12505 5466
rect 12529 5414 12539 5466
rect 12539 5414 12585 5466
rect 12609 5414 12655 5466
rect 12655 5414 12665 5466
rect 12689 5414 12719 5466
rect 12719 5414 12745 5466
rect 12449 5412 12505 5414
rect 12529 5412 12585 5414
rect 12609 5412 12665 5414
rect 12689 5412 12745 5414
rect 12438 5208 12494 5264
rect 12449 4378 12505 4380
rect 12529 4378 12585 4380
rect 12609 4378 12665 4380
rect 12689 4378 12745 4380
rect 12449 4326 12475 4378
rect 12475 4326 12505 4378
rect 12529 4326 12539 4378
rect 12539 4326 12585 4378
rect 12609 4326 12655 4378
rect 12655 4326 12665 4378
rect 12689 4326 12719 4378
rect 12719 4326 12745 4378
rect 12449 4324 12505 4326
rect 12529 4324 12585 4326
rect 12609 4324 12665 4326
rect 12689 4324 12745 4326
rect 12254 4120 12310 4176
rect 12162 2488 12218 2544
rect 12346 3732 12402 3768
rect 12346 3712 12348 3732
rect 12348 3712 12400 3732
rect 12400 3712 12402 3732
rect 12449 3290 12505 3292
rect 12529 3290 12585 3292
rect 12609 3290 12665 3292
rect 12689 3290 12745 3292
rect 12449 3238 12475 3290
rect 12475 3238 12505 3290
rect 12529 3238 12539 3290
rect 12539 3238 12585 3290
rect 12609 3238 12655 3290
rect 12655 3238 12665 3290
rect 12689 3238 12719 3290
rect 12719 3238 12745 3290
rect 12449 3236 12505 3238
rect 12529 3236 12585 3238
rect 12609 3236 12665 3238
rect 12689 3236 12745 3238
rect 12990 3032 13046 3088
rect 13358 5072 13414 5128
rect 11610 856 11666 912
rect 12449 2202 12505 2204
rect 12529 2202 12585 2204
rect 12609 2202 12665 2204
rect 12689 2202 12745 2204
rect 12449 2150 12475 2202
rect 12475 2150 12505 2202
rect 12529 2150 12539 2202
rect 12539 2150 12585 2202
rect 12609 2150 12655 2202
rect 12655 2150 12665 2202
rect 12689 2150 12719 2202
rect 12719 2150 12745 2202
rect 12449 2148 12505 2150
rect 12529 2148 12585 2150
rect 12609 2148 12665 2150
rect 12689 2148 12745 2150
rect 13634 8200 13690 8256
rect 13634 7248 13690 7304
rect 13542 5752 13598 5808
rect 13542 5344 13598 5400
rect 13634 4936 13690 4992
rect 13542 4120 13598 4176
rect 13726 4528 13782 4584
rect 14646 3576 14702 3632
rect 12622 176 12678 232
<< metal3 >>
rect 0 15874 480 15904
rect 3325 15874 3391 15877
rect 0 15872 3391 15874
rect 0 15816 3330 15872
rect 3386 15816 3391 15872
rect 0 15814 3391 15816
rect 0 15784 480 15814
rect 3325 15811 3391 15814
rect 11605 15874 11671 15877
rect 15520 15874 16000 15904
rect 11605 15872 16000 15874
rect 11605 15816 11610 15872
rect 11666 15816 16000 15872
rect 11605 15814 16000 15816
rect 11605 15811 11671 15814
rect 15520 15784 16000 15814
rect 0 15466 480 15496
rect 6453 15466 6519 15469
rect 0 15464 6519 15466
rect 0 15408 6458 15464
rect 6514 15408 6519 15464
rect 0 15406 6519 15408
rect 0 15376 480 15406
rect 6453 15403 6519 15406
rect 11973 15466 12039 15469
rect 15520 15466 16000 15496
rect 11973 15464 16000 15466
rect 11973 15408 11978 15464
rect 12034 15408 16000 15464
rect 11973 15406 16000 15408
rect 11973 15403 12039 15406
rect 15520 15376 16000 15406
rect 0 15058 480 15088
rect 2589 15058 2655 15061
rect 0 15056 2655 15058
rect 0 15000 2594 15056
rect 2650 15000 2655 15056
rect 0 14998 2655 15000
rect 0 14968 480 14998
rect 2589 14995 2655 14998
rect 11053 15058 11119 15061
rect 15520 15058 16000 15088
rect 11053 15056 16000 15058
rect 11053 15000 11058 15056
rect 11114 15000 16000 15056
rect 11053 14998 16000 15000
rect 11053 14995 11119 14998
rect 15520 14968 16000 14998
rect 0 14650 480 14680
rect 1485 14650 1551 14653
rect 0 14648 1551 14650
rect 0 14592 1490 14648
rect 1546 14592 1551 14648
rect 0 14590 1551 14592
rect 0 14560 480 14590
rect 1485 14587 1551 14590
rect 11237 14650 11303 14653
rect 15520 14650 16000 14680
rect 11237 14648 16000 14650
rect 11237 14592 11242 14648
rect 11298 14592 16000 14648
rect 11237 14590 16000 14592
rect 11237 14587 11303 14590
rect 15520 14560 16000 14590
rect 0 14242 480 14272
rect 4061 14242 4127 14245
rect 0 14240 4127 14242
rect 0 14184 4066 14240
rect 4122 14184 4127 14240
rect 0 14182 4127 14184
rect 0 14152 480 14182
rect 4061 14179 4127 14182
rect 11145 14242 11211 14245
rect 15520 14242 16000 14272
rect 11145 14240 16000 14242
rect 11145 14184 11150 14240
rect 11206 14184 16000 14240
rect 11145 14182 16000 14184
rect 11145 14179 11211 14182
rect 15520 14152 16000 14182
rect 0 13834 480 13864
rect 4061 13834 4127 13837
rect 0 13832 4127 13834
rect 0 13776 4066 13832
rect 4122 13776 4127 13832
rect 0 13774 4127 13776
rect 0 13744 480 13774
rect 4061 13771 4127 13774
rect 10685 13834 10751 13837
rect 15520 13834 16000 13864
rect 10685 13832 16000 13834
rect 10685 13776 10690 13832
rect 10746 13776 16000 13832
rect 10685 13774 16000 13776
rect 10685 13771 10751 13774
rect 15520 13744 16000 13774
rect 5541 13632 5861 13633
rect 5541 13568 5549 13632
rect 5613 13568 5629 13632
rect 5693 13568 5709 13632
rect 5773 13568 5789 13632
rect 5853 13568 5861 13632
rect 5541 13567 5861 13568
rect 10138 13632 10458 13633
rect 10138 13568 10146 13632
rect 10210 13568 10226 13632
rect 10290 13568 10306 13632
rect 10370 13568 10386 13632
rect 10450 13568 10458 13632
rect 10138 13567 10458 13568
rect 0 13426 480 13456
rect 3877 13426 3943 13429
rect 0 13424 3943 13426
rect 0 13368 3882 13424
rect 3938 13368 3943 13424
rect 0 13366 3943 13368
rect 0 13336 480 13366
rect 3877 13363 3943 13366
rect 12893 13426 12959 13429
rect 15520 13426 16000 13456
rect 12893 13424 16000 13426
rect 12893 13368 12898 13424
rect 12954 13368 16000 13424
rect 12893 13366 16000 13368
rect 12893 13363 12959 13366
rect 15520 13336 16000 13366
rect 3242 13088 3562 13089
rect 0 13018 480 13048
rect 3242 13024 3250 13088
rect 3314 13024 3330 13088
rect 3394 13024 3410 13088
rect 3474 13024 3490 13088
rect 3554 13024 3562 13088
rect 3242 13023 3562 13024
rect 7840 13088 8160 13089
rect 7840 13024 7848 13088
rect 7912 13024 7928 13088
rect 7992 13024 8008 13088
rect 8072 13024 8088 13088
rect 8152 13024 8160 13088
rect 7840 13023 8160 13024
rect 12437 13088 12757 13089
rect 12437 13024 12445 13088
rect 12509 13024 12525 13088
rect 12589 13024 12605 13088
rect 12669 13024 12685 13088
rect 12749 13024 12757 13088
rect 12437 13023 12757 13024
rect 3049 13018 3115 13021
rect 15520 13018 16000 13048
rect 0 13016 3115 13018
rect 0 12960 3054 13016
rect 3110 12960 3115 13016
rect 0 12958 3115 12960
rect 0 12928 480 12958
rect 3049 12955 3115 12958
rect 12942 12958 16000 13018
rect 9765 12884 9831 12885
rect 9765 12880 9812 12884
rect 9876 12882 9882 12884
rect 11237 12882 11303 12885
rect 12942 12882 13002 12958
rect 15520 12928 16000 12958
rect 9765 12824 9770 12880
rect 9765 12820 9812 12824
rect 9876 12822 9922 12882
rect 11237 12880 13002 12882
rect 11237 12824 11242 12880
rect 11298 12824 13002 12880
rect 11237 12822 13002 12824
rect 9876 12820 9882 12822
rect 9765 12819 9831 12820
rect 11237 12819 11303 12822
rect 2129 12746 2195 12749
rect 7189 12746 7255 12749
rect 8937 12746 9003 12749
rect 2129 12744 9003 12746
rect 2129 12688 2134 12744
rect 2190 12688 7194 12744
rect 7250 12688 8942 12744
rect 8998 12688 9003 12744
rect 2129 12686 9003 12688
rect 2129 12683 2195 12686
rect 7189 12683 7255 12686
rect 8937 12683 9003 12686
rect 9857 12746 9923 12749
rect 12893 12746 12959 12749
rect 9857 12744 12959 12746
rect 9857 12688 9862 12744
rect 9918 12688 12898 12744
rect 12954 12688 12959 12744
rect 9857 12686 12959 12688
rect 9857 12683 9923 12686
rect 12893 12683 12959 12686
rect 0 12610 480 12640
rect 3509 12610 3575 12613
rect 0 12608 3575 12610
rect 0 12552 3514 12608
rect 3570 12552 3575 12608
rect 0 12550 3575 12552
rect 0 12520 480 12550
rect 3509 12547 3575 12550
rect 11053 12610 11119 12613
rect 15520 12610 16000 12640
rect 11053 12608 16000 12610
rect 11053 12552 11058 12608
rect 11114 12552 16000 12608
rect 11053 12550 16000 12552
rect 11053 12547 11119 12550
rect 5541 12544 5861 12545
rect 5541 12480 5549 12544
rect 5613 12480 5629 12544
rect 5693 12480 5709 12544
rect 5773 12480 5789 12544
rect 5853 12480 5861 12544
rect 5541 12479 5861 12480
rect 10138 12544 10458 12545
rect 10138 12480 10146 12544
rect 10210 12480 10226 12544
rect 10290 12480 10306 12544
rect 10370 12480 10386 12544
rect 10450 12480 10458 12544
rect 15520 12520 16000 12550
rect 10138 12479 10458 12480
rect 2814 12412 2820 12476
rect 2884 12474 2890 12476
rect 3233 12474 3299 12477
rect 2884 12472 3299 12474
rect 2884 12416 3238 12472
rect 3294 12416 3299 12472
rect 2884 12414 3299 12416
rect 2884 12412 2890 12414
rect 3233 12411 3299 12414
rect 4245 12338 4311 12341
rect 6085 12338 6151 12341
rect 4245 12336 6151 12338
rect 4245 12280 4250 12336
rect 4306 12280 6090 12336
rect 6146 12280 6151 12336
rect 4245 12278 6151 12280
rect 4245 12275 4311 12278
rect 6085 12275 6151 12278
rect 8477 12338 8543 12341
rect 11237 12338 11303 12341
rect 8477 12336 11303 12338
rect 8477 12280 8482 12336
rect 8538 12280 11242 12336
rect 11298 12280 11303 12336
rect 8477 12278 11303 12280
rect 8477 12275 8543 12278
rect 11237 12275 11303 12278
rect 0 12202 480 12232
rect 4705 12202 4771 12205
rect 0 12200 4771 12202
rect 0 12144 4710 12200
rect 4766 12144 4771 12200
rect 0 12142 4771 12144
rect 0 12112 480 12142
rect 4705 12139 4771 12142
rect 5165 12202 5231 12205
rect 10685 12202 10751 12205
rect 5165 12200 10751 12202
rect 5165 12144 5170 12200
rect 5226 12144 10690 12200
rect 10746 12144 10751 12200
rect 5165 12142 10751 12144
rect 5165 12139 5231 12142
rect 10685 12139 10751 12142
rect 11053 12202 11119 12205
rect 15520 12202 16000 12232
rect 11053 12200 16000 12202
rect 11053 12144 11058 12200
rect 11114 12144 16000 12200
rect 11053 12142 16000 12144
rect 11053 12139 11119 12142
rect 15520 12112 16000 12142
rect 9673 12066 9739 12069
rect 10961 12066 11027 12069
rect 9673 12064 11027 12066
rect 9673 12008 9678 12064
rect 9734 12008 10966 12064
rect 11022 12008 11027 12064
rect 9673 12006 11027 12008
rect 9673 12003 9739 12006
rect 10961 12003 11027 12006
rect 3242 12000 3562 12001
rect 3242 11936 3250 12000
rect 3314 11936 3330 12000
rect 3394 11936 3410 12000
rect 3474 11936 3490 12000
rect 3554 11936 3562 12000
rect 3242 11935 3562 11936
rect 7840 12000 8160 12001
rect 7840 11936 7848 12000
rect 7912 11936 7928 12000
rect 7992 11936 8008 12000
rect 8072 11936 8088 12000
rect 8152 11936 8160 12000
rect 7840 11935 8160 11936
rect 12437 12000 12757 12001
rect 12437 11936 12445 12000
rect 12509 11936 12525 12000
rect 12589 11936 12605 12000
rect 12669 11936 12685 12000
rect 12749 11936 12757 12000
rect 12437 11935 12757 11936
rect 0 11794 480 11824
rect 5073 11794 5139 11797
rect 0 11792 5139 11794
rect 0 11736 5078 11792
rect 5134 11736 5139 11792
rect 0 11734 5139 11736
rect 0 11704 480 11734
rect 5073 11731 5139 11734
rect 11053 11794 11119 11797
rect 15520 11794 16000 11824
rect 11053 11792 16000 11794
rect 11053 11736 11058 11792
rect 11114 11736 16000 11792
rect 11053 11734 16000 11736
rect 11053 11731 11119 11734
rect 15520 11704 16000 11734
rect 5541 11456 5861 11457
rect 0 11386 480 11416
rect 5541 11392 5549 11456
rect 5613 11392 5629 11456
rect 5693 11392 5709 11456
rect 5773 11392 5789 11456
rect 5853 11392 5861 11456
rect 5541 11391 5861 11392
rect 10138 11456 10458 11457
rect 10138 11392 10146 11456
rect 10210 11392 10226 11456
rect 10290 11392 10306 11456
rect 10370 11392 10386 11456
rect 10450 11392 10458 11456
rect 10138 11391 10458 11392
rect 11053 11386 11119 11389
rect 15520 11386 16000 11416
rect 0 11326 5458 11386
rect 0 11296 480 11326
rect 3734 11188 3740 11252
rect 3804 11250 3810 11252
rect 3877 11250 3943 11253
rect 3804 11248 3943 11250
rect 3804 11192 3882 11248
rect 3938 11192 3943 11248
rect 3804 11190 3943 11192
rect 5398 11250 5458 11326
rect 11053 11384 16000 11386
rect 11053 11328 11058 11384
rect 11114 11328 16000 11384
rect 11053 11326 16000 11328
rect 11053 11323 11119 11326
rect 15520 11296 16000 11326
rect 6453 11250 6519 11253
rect 5398 11248 6519 11250
rect 5398 11192 6458 11248
rect 6514 11192 6519 11248
rect 5398 11190 6519 11192
rect 3804 11188 3810 11190
rect 3877 11187 3943 11190
rect 6453 11187 6519 11190
rect 2681 11114 2747 11117
rect 4102 11114 4108 11116
rect 2681 11112 4108 11114
rect 2681 11056 2686 11112
rect 2742 11056 4108 11112
rect 2681 11054 4108 11056
rect 2681 11051 2747 11054
rect 4102 11052 4108 11054
rect 4172 11052 4178 11116
rect 0 10978 480 11008
rect 3049 10978 3115 10981
rect 3969 10980 4035 10981
rect 3918 10978 3924 10980
rect 0 10976 3115 10978
rect 0 10920 3054 10976
rect 3110 10920 3115 10976
rect 0 10918 3115 10920
rect 3878 10918 3924 10978
rect 3988 10976 4035 10980
rect 15520 10978 16000 11008
rect 4030 10920 4035 10976
rect 0 10888 480 10918
rect 3049 10915 3115 10918
rect 3918 10916 3924 10918
rect 3988 10916 4035 10920
rect 3969 10915 4035 10916
rect 13862 10918 16000 10978
rect 3242 10912 3562 10913
rect 3242 10848 3250 10912
rect 3314 10848 3330 10912
rect 3394 10848 3410 10912
rect 3474 10848 3490 10912
rect 3554 10848 3562 10912
rect 3242 10847 3562 10848
rect 7840 10912 8160 10913
rect 7840 10848 7848 10912
rect 7912 10848 7928 10912
rect 7992 10848 8008 10912
rect 8072 10848 8088 10912
rect 8152 10848 8160 10912
rect 7840 10847 8160 10848
rect 12437 10912 12757 10913
rect 12437 10848 12445 10912
rect 12509 10848 12525 10912
rect 12589 10848 12605 10912
rect 12669 10848 12685 10912
rect 12749 10848 12757 10912
rect 12437 10847 12757 10848
rect 11053 10706 11119 10709
rect 13862 10706 13922 10918
rect 15520 10888 16000 10918
rect 11053 10704 13922 10706
rect 11053 10648 11058 10704
rect 11114 10648 13922 10704
rect 11053 10646 13922 10648
rect 11053 10643 11119 10646
rect 0 10570 480 10600
rect 7097 10570 7163 10573
rect 8201 10570 8267 10573
rect 0 10568 8267 10570
rect 0 10512 7102 10568
rect 7158 10512 8206 10568
rect 8262 10512 8267 10568
rect 0 10510 8267 10512
rect 0 10480 480 10510
rect 7097 10507 7163 10510
rect 8201 10507 8267 10510
rect 12249 10570 12315 10573
rect 15520 10570 16000 10600
rect 12249 10568 16000 10570
rect 12249 10512 12254 10568
rect 12310 10512 16000 10568
rect 12249 10510 16000 10512
rect 12249 10507 12315 10510
rect 15520 10480 16000 10510
rect 5541 10368 5861 10369
rect 5541 10304 5549 10368
rect 5613 10304 5629 10368
rect 5693 10304 5709 10368
rect 5773 10304 5789 10368
rect 5853 10304 5861 10368
rect 5541 10303 5861 10304
rect 10138 10368 10458 10369
rect 10138 10304 10146 10368
rect 10210 10304 10226 10368
rect 10290 10304 10306 10368
rect 10370 10304 10386 10368
rect 10450 10304 10458 10368
rect 10138 10303 10458 10304
rect 2957 10300 3023 10301
rect 2957 10298 3004 10300
rect 2912 10296 3004 10298
rect 2912 10240 2962 10296
rect 2912 10238 3004 10240
rect 2957 10236 3004 10238
rect 3068 10236 3074 10300
rect 7005 10298 7071 10301
rect 9121 10298 9187 10301
rect 7005 10296 9187 10298
rect 7005 10240 7010 10296
rect 7066 10240 9126 10296
rect 9182 10240 9187 10296
rect 7005 10238 9187 10240
rect 2957 10235 3023 10236
rect 7005 10235 7071 10238
rect 9121 10235 9187 10238
rect 0 10162 480 10192
rect 3969 10162 4035 10165
rect 0 10160 4035 10162
rect 0 10104 3974 10160
rect 4030 10104 4035 10160
rect 0 10102 4035 10104
rect 0 10072 480 10102
rect 3969 10099 4035 10102
rect 10041 10162 10107 10165
rect 15520 10162 16000 10192
rect 10041 10160 16000 10162
rect 10041 10104 10046 10160
rect 10102 10104 16000 10160
rect 10041 10102 16000 10104
rect 10041 10099 10107 10102
rect 15520 10072 16000 10102
rect 2405 10026 2471 10029
rect 3141 10026 3207 10029
rect 2405 10024 3207 10026
rect 2405 9968 2410 10024
rect 2466 9968 3146 10024
rect 3202 9968 3207 10024
rect 2405 9966 3207 9968
rect 2405 9963 2471 9966
rect 3141 9963 3207 9966
rect 9305 10026 9371 10029
rect 11697 10026 11763 10029
rect 9305 10024 11763 10026
rect 9305 9968 9310 10024
rect 9366 9968 11702 10024
rect 11758 9968 11763 10024
rect 9305 9966 11763 9968
rect 9305 9963 9371 9966
rect 11697 9963 11763 9966
rect 12198 9964 12204 10028
rect 12268 10026 12274 10028
rect 12268 9966 13922 10026
rect 12268 9964 12274 9966
rect 3242 9824 3562 9825
rect 0 9754 480 9784
rect 3242 9760 3250 9824
rect 3314 9760 3330 9824
rect 3394 9760 3410 9824
rect 3474 9760 3490 9824
rect 3554 9760 3562 9824
rect 3242 9759 3562 9760
rect 7840 9824 8160 9825
rect 7840 9760 7848 9824
rect 7912 9760 7928 9824
rect 7992 9760 8008 9824
rect 8072 9760 8088 9824
rect 8152 9760 8160 9824
rect 7840 9759 8160 9760
rect 12437 9824 12757 9825
rect 12437 9760 12445 9824
rect 12509 9760 12525 9824
rect 12589 9760 12605 9824
rect 12669 9760 12685 9824
rect 12749 9760 12757 9824
rect 12437 9759 12757 9760
rect 10041 9754 10107 9757
rect 10961 9754 11027 9757
rect 0 9694 3066 9754
rect 0 9664 480 9694
rect 3006 9618 3066 9694
rect 10041 9752 11027 9754
rect 10041 9696 10046 9752
rect 10102 9696 10966 9752
rect 11022 9696 11027 9752
rect 10041 9694 11027 9696
rect 13862 9754 13922 9966
rect 15520 9754 16000 9784
rect 13862 9694 16000 9754
rect 10041 9691 10107 9694
rect 10961 9691 11027 9694
rect 15520 9664 16000 9694
rect 4470 9618 4476 9620
rect 3006 9558 4476 9618
rect 4470 9556 4476 9558
rect 4540 9556 4546 9620
rect 7557 9618 7623 9621
rect 7557 9616 7666 9618
rect 7557 9560 7562 9616
rect 7618 9560 7666 9616
rect 7557 9555 7666 9560
rect 7189 9482 7255 9485
rect 7465 9482 7531 9485
rect 7189 9480 7531 9482
rect 7189 9424 7194 9480
rect 7250 9424 7470 9480
rect 7526 9424 7531 9480
rect 7189 9422 7531 9424
rect 7189 9419 7255 9422
rect 7465 9419 7531 9422
rect 0 9346 480 9376
rect 1761 9346 1827 9349
rect 2681 9346 2747 9349
rect 0 9344 2747 9346
rect 0 9288 1766 9344
rect 1822 9288 2686 9344
rect 2742 9288 2747 9344
rect 0 9286 2747 9288
rect 0 9256 480 9286
rect 1761 9283 1827 9286
rect 2681 9283 2747 9286
rect 2814 9284 2820 9348
rect 2884 9346 2890 9348
rect 3601 9346 3667 9349
rect 2884 9344 3667 9346
rect 2884 9288 3606 9344
rect 3662 9288 3667 9344
rect 2884 9286 3667 9288
rect 2884 9284 2890 9286
rect 3601 9283 3667 9286
rect 7465 9346 7531 9349
rect 7606 9346 7666 9555
rect 7465 9344 7666 9346
rect 7465 9288 7470 9344
rect 7526 9288 7666 9344
rect 7465 9286 7666 9288
rect 11053 9346 11119 9349
rect 15520 9346 16000 9376
rect 11053 9344 16000 9346
rect 11053 9288 11058 9344
rect 11114 9288 16000 9344
rect 11053 9286 16000 9288
rect 7465 9283 7531 9286
rect 11053 9283 11119 9286
rect 5541 9280 5861 9281
rect 5541 9216 5549 9280
rect 5613 9216 5629 9280
rect 5693 9216 5709 9280
rect 5773 9216 5789 9280
rect 5853 9216 5861 9280
rect 5541 9215 5861 9216
rect 10138 9280 10458 9281
rect 10138 9216 10146 9280
rect 10210 9216 10226 9280
rect 10290 9216 10306 9280
rect 10370 9216 10386 9280
rect 10450 9216 10458 9280
rect 15520 9256 16000 9286
rect 10138 9215 10458 9216
rect 2773 9074 2839 9077
rect 8569 9074 8635 9077
rect 2773 9072 8635 9074
rect 2773 9016 2778 9072
rect 2834 9016 8574 9072
rect 8630 9016 8635 9072
rect 2773 9014 8635 9016
rect 2773 9011 2839 9014
rect 8569 9011 8635 9014
rect 0 8938 480 8968
rect 4286 8938 4292 8940
rect 0 8878 4292 8938
rect 0 8848 480 8878
rect 4286 8876 4292 8878
rect 4356 8938 4362 8940
rect 5073 8938 5139 8941
rect 4356 8936 5139 8938
rect 4356 8880 5078 8936
rect 5134 8880 5139 8936
rect 4356 8878 5139 8880
rect 4356 8876 4362 8878
rect 5073 8875 5139 8878
rect 12249 8938 12315 8941
rect 15520 8938 16000 8968
rect 12249 8936 16000 8938
rect 12249 8880 12254 8936
rect 12310 8880 16000 8936
rect 12249 8878 16000 8880
rect 12249 8875 12315 8878
rect 15520 8848 16000 8878
rect 3242 8736 3562 8737
rect 3242 8672 3250 8736
rect 3314 8672 3330 8736
rect 3394 8672 3410 8736
rect 3474 8672 3490 8736
rect 3554 8672 3562 8736
rect 3242 8671 3562 8672
rect 7840 8736 8160 8737
rect 7840 8672 7848 8736
rect 7912 8672 7928 8736
rect 7992 8672 8008 8736
rect 8072 8672 8088 8736
rect 8152 8672 8160 8736
rect 7840 8671 8160 8672
rect 12437 8736 12757 8737
rect 12437 8672 12445 8736
rect 12509 8672 12525 8736
rect 12589 8672 12605 8736
rect 12669 8672 12685 8736
rect 12749 8672 12757 8736
rect 12437 8671 12757 8672
rect 11329 8668 11395 8669
rect 11278 8666 11284 8668
rect 11238 8606 11284 8666
rect 11348 8664 11395 8668
rect 11390 8608 11395 8664
rect 11278 8604 11284 8606
rect 11348 8604 11395 8608
rect 11329 8603 11395 8604
rect 0 8530 480 8560
rect 5073 8530 5139 8533
rect 0 8528 5139 8530
rect 0 8472 5078 8528
rect 5134 8472 5139 8528
rect 0 8470 5139 8472
rect 0 8440 480 8470
rect 5073 8467 5139 8470
rect 11421 8530 11487 8533
rect 13169 8530 13235 8533
rect 15520 8530 16000 8560
rect 11421 8528 16000 8530
rect 11421 8472 11426 8528
rect 11482 8472 13174 8528
rect 13230 8472 16000 8528
rect 11421 8470 16000 8472
rect 11421 8467 11487 8470
rect 13169 8467 13235 8470
rect 15520 8440 16000 8470
rect 0 8258 480 8288
rect 1117 8258 1183 8261
rect 0 8256 1183 8258
rect 0 8200 1122 8256
rect 1178 8200 1183 8256
rect 0 8198 1183 8200
rect 0 8168 480 8198
rect 1117 8195 1183 8198
rect 13629 8258 13695 8261
rect 15520 8258 16000 8288
rect 13629 8256 16000 8258
rect 13629 8200 13634 8256
rect 13690 8200 16000 8256
rect 13629 8198 16000 8200
rect 13629 8195 13695 8198
rect 5541 8192 5861 8193
rect 5541 8128 5549 8192
rect 5613 8128 5629 8192
rect 5693 8128 5709 8192
rect 5773 8128 5789 8192
rect 5853 8128 5861 8192
rect 5541 8127 5861 8128
rect 10138 8192 10458 8193
rect 10138 8128 10146 8192
rect 10210 8128 10226 8192
rect 10290 8128 10306 8192
rect 10370 8128 10386 8192
rect 10450 8128 10458 8192
rect 15520 8168 16000 8198
rect 10138 8127 10458 8128
rect 11789 8124 11855 8125
rect 11789 8120 11836 8124
rect 11900 8122 11906 8124
rect 11789 8064 11794 8120
rect 11789 8060 11836 8064
rect 11900 8062 11946 8122
rect 11900 8060 11906 8062
rect 11789 8059 11855 8060
rect 933 7986 999 7989
rect 8661 7986 8727 7989
rect 933 7984 8727 7986
rect 933 7928 938 7984
rect 994 7928 8666 7984
rect 8722 7928 8727 7984
rect 933 7926 8727 7928
rect 933 7923 999 7926
rect 8661 7923 8727 7926
rect 0 7850 480 7880
rect 3969 7850 4035 7853
rect 0 7848 4035 7850
rect 0 7792 3974 7848
rect 4030 7792 4035 7848
rect 0 7790 4035 7792
rect 0 7760 480 7790
rect 3969 7787 4035 7790
rect 11053 7850 11119 7853
rect 15520 7850 16000 7880
rect 11053 7848 16000 7850
rect 11053 7792 11058 7848
rect 11114 7792 16000 7848
rect 11053 7790 16000 7792
rect 11053 7787 11119 7790
rect 15520 7760 16000 7790
rect 3242 7648 3562 7649
rect 3242 7584 3250 7648
rect 3314 7584 3330 7648
rect 3394 7584 3410 7648
rect 3474 7584 3490 7648
rect 3554 7584 3562 7648
rect 3242 7583 3562 7584
rect 7840 7648 8160 7649
rect 7840 7584 7848 7648
rect 7912 7584 7928 7648
rect 7992 7584 8008 7648
rect 8072 7584 8088 7648
rect 8152 7584 8160 7648
rect 7840 7583 8160 7584
rect 12437 7648 12757 7649
rect 12437 7584 12445 7648
rect 12509 7584 12525 7648
rect 12589 7584 12605 7648
rect 12669 7584 12685 7648
rect 12749 7584 12757 7648
rect 12437 7583 12757 7584
rect 0 7442 480 7472
rect 3417 7442 3483 7445
rect 0 7440 3483 7442
rect 0 7384 3422 7440
rect 3478 7384 3483 7440
rect 0 7382 3483 7384
rect 0 7352 480 7382
rect 3417 7379 3483 7382
rect 12341 7442 12407 7445
rect 15520 7442 16000 7472
rect 12341 7440 16000 7442
rect 12341 7384 12346 7440
rect 12402 7384 16000 7440
rect 12341 7382 16000 7384
rect 12341 7379 12407 7382
rect 15520 7352 16000 7382
rect 1485 7306 1551 7309
rect 9121 7306 9187 7309
rect 1485 7304 9187 7306
rect 1485 7248 1490 7304
rect 1546 7248 9126 7304
rect 9182 7248 9187 7304
rect 1485 7246 9187 7248
rect 1485 7243 1551 7246
rect 9121 7243 9187 7246
rect 11053 7306 11119 7309
rect 13629 7306 13695 7309
rect 11053 7304 13695 7306
rect 11053 7248 11058 7304
rect 11114 7248 13634 7304
rect 13690 7248 13695 7304
rect 11053 7246 13695 7248
rect 11053 7243 11119 7246
rect 13629 7243 13695 7246
rect 3969 7170 4035 7173
rect 11789 7172 11855 7173
rect 11789 7170 11836 7172
rect 1350 7168 4035 7170
rect 1350 7112 3974 7168
rect 4030 7112 4035 7168
rect 1350 7110 4035 7112
rect 11744 7168 11836 7170
rect 11744 7112 11794 7168
rect 11744 7110 11836 7112
rect 0 7034 480 7064
rect 1350 7034 1410 7110
rect 3969 7107 4035 7110
rect 11789 7108 11836 7110
rect 11900 7108 11906 7172
rect 11789 7107 11855 7108
rect 5541 7104 5861 7105
rect 5541 7040 5549 7104
rect 5613 7040 5629 7104
rect 5693 7040 5709 7104
rect 5773 7040 5789 7104
rect 5853 7040 5861 7104
rect 5541 7039 5861 7040
rect 10138 7104 10458 7105
rect 10138 7040 10146 7104
rect 10210 7040 10226 7104
rect 10290 7040 10306 7104
rect 10370 7040 10386 7104
rect 10450 7040 10458 7104
rect 10138 7039 10458 7040
rect 0 6974 1410 7034
rect 11513 7034 11579 7037
rect 15520 7034 16000 7064
rect 11513 7032 16000 7034
rect 11513 6976 11518 7032
rect 11574 6976 16000 7032
rect 11513 6974 16000 6976
rect 0 6944 480 6974
rect 11513 6971 11579 6974
rect 15520 6944 16000 6974
rect 11053 6898 11119 6901
rect 11053 6896 13922 6898
rect 11053 6840 11058 6896
rect 11114 6840 13922 6896
rect 11053 6838 13922 6840
rect 11053 6835 11119 6838
rect 5073 6762 5139 6765
rect 7230 6762 7236 6764
rect 5073 6760 7236 6762
rect 5073 6704 5078 6760
rect 5134 6704 7236 6760
rect 5073 6702 7236 6704
rect 5073 6699 5139 6702
rect 7230 6700 7236 6702
rect 7300 6762 7306 6764
rect 8937 6762 9003 6765
rect 7300 6760 9003 6762
rect 7300 6704 8942 6760
rect 8998 6704 9003 6760
rect 7300 6702 9003 6704
rect 7300 6700 7306 6702
rect 8937 6699 9003 6702
rect 0 6626 480 6656
rect 841 6626 907 6629
rect 0 6624 907 6626
rect 0 6568 846 6624
rect 902 6568 907 6624
rect 0 6566 907 6568
rect 13862 6626 13922 6838
rect 15520 6626 16000 6656
rect 13862 6566 16000 6626
rect 0 6536 480 6566
rect 841 6563 907 6566
rect 3242 6560 3562 6561
rect 3242 6496 3250 6560
rect 3314 6496 3330 6560
rect 3394 6496 3410 6560
rect 3474 6496 3490 6560
rect 3554 6496 3562 6560
rect 3242 6495 3562 6496
rect 7840 6560 8160 6561
rect 7840 6496 7848 6560
rect 7912 6496 7928 6560
rect 7992 6496 8008 6560
rect 8072 6496 8088 6560
rect 8152 6496 8160 6560
rect 7840 6495 8160 6496
rect 12437 6560 12757 6561
rect 12437 6496 12445 6560
rect 12509 6496 12525 6560
rect 12589 6496 12605 6560
rect 12669 6496 12685 6560
rect 12749 6496 12757 6560
rect 15520 6536 16000 6566
rect 12437 6495 12757 6496
rect 4061 6490 4127 6493
rect 4797 6490 4863 6493
rect 4061 6488 4863 6490
rect 4061 6432 4066 6488
rect 4122 6432 4802 6488
rect 4858 6432 4863 6488
rect 4061 6430 4863 6432
rect 4061 6427 4127 6430
rect 4797 6427 4863 6430
rect 6545 6354 6611 6357
rect 8661 6354 8727 6357
rect 6545 6352 8727 6354
rect 6545 6296 6550 6352
rect 6606 6296 8666 6352
rect 8722 6296 8727 6352
rect 6545 6294 8727 6296
rect 6545 6291 6611 6294
rect 8661 6291 8727 6294
rect 0 6218 480 6248
rect 4061 6218 4127 6221
rect 10869 6218 10935 6221
rect 15520 6218 16000 6248
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 480 6158
rect 4061 6155 4127 6158
rect 5398 6158 6010 6218
rect 1945 6082 2011 6085
rect 5398 6082 5458 6158
rect 1945 6080 5458 6082
rect 1945 6024 1950 6080
rect 2006 6024 5458 6080
rect 1945 6022 5458 6024
rect 5950 6082 6010 6158
rect 10869 6216 16000 6218
rect 10869 6160 10874 6216
rect 10930 6160 16000 6216
rect 10869 6158 16000 6160
rect 10869 6155 10935 6158
rect 15520 6128 16000 6158
rect 8661 6082 8727 6085
rect 5950 6080 8727 6082
rect 5950 6024 8666 6080
rect 8722 6024 8727 6080
rect 5950 6022 8727 6024
rect 1945 6019 2011 6022
rect 8661 6019 8727 6022
rect 5541 6016 5861 6017
rect 5541 5952 5549 6016
rect 5613 5952 5629 6016
rect 5693 5952 5709 6016
rect 5773 5952 5789 6016
rect 5853 5952 5861 6016
rect 5541 5951 5861 5952
rect 10138 6016 10458 6017
rect 10138 5952 10146 6016
rect 10210 5952 10226 6016
rect 10290 5952 10306 6016
rect 10370 5952 10386 6016
rect 10450 5952 10458 6016
rect 10138 5951 10458 5952
rect 1761 5946 1827 5949
rect 6085 5946 6151 5949
rect 6269 5946 6335 5949
rect 9581 5946 9647 5949
rect 1761 5944 5274 5946
rect 1761 5888 1766 5944
rect 1822 5888 5274 5944
rect 1761 5886 5274 5888
rect 1761 5883 1827 5886
rect 0 5810 480 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 480 5750
rect 4061 5747 4127 5750
rect 1669 5674 1735 5677
rect 5214 5674 5274 5886
rect 6085 5944 9647 5946
rect 6085 5888 6090 5944
rect 6146 5888 6274 5944
rect 6330 5888 9586 5944
rect 9642 5888 9647 5944
rect 6085 5886 9647 5888
rect 6085 5883 6151 5886
rect 6269 5883 6335 5886
rect 9581 5883 9647 5886
rect 5349 5810 5415 5813
rect 9581 5810 9647 5813
rect 5349 5808 9647 5810
rect 5349 5752 5354 5808
rect 5410 5752 9586 5808
rect 9642 5752 9647 5808
rect 5349 5750 9647 5752
rect 5349 5747 5415 5750
rect 9581 5747 9647 5750
rect 13537 5810 13603 5813
rect 15520 5810 16000 5840
rect 13537 5808 16000 5810
rect 13537 5752 13542 5808
rect 13598 5752 16000 5808
rect 13537 5750 16000 5752
rect 13537 5747 13603 5750
rect 15520 5720 16000 5750
rect 7281 5674 7347 5677
rect 1669 5672 1962 5674
rect 1669 5616 1674 5672
rect 1730 5616 1962 5672
rect 1669 5614 1962 5616
rect 5214 5672 7347 5674
rect 5214 5616 7286 5672
rect 7342 5616 7347 5672
rect 5214 5614 7347 5616
rect 1669 5611 1735 5614
rect 1902 5541 1962 5614
rect 7281 5611 7347 5614
rect 1902 5536 2011 5541
rect 1902 5480 1950 5536
rect 2006 5480 2011 5536
rect 1902 5478 2011 5480
rect 1945 5475 2011 5478
rect 3242 5472 3562 5473
rect 0 5402 480 5432
rect 3242 5408 3250 5472
rect 3314 5408 3330 5472
rect 3394 5408 3410 5472
rect 3474 5408 3490 5472
rect 3554 5408 3562 5472
rect 3242 5407 3562 5408
rect 7840 5472 8160 5473
rect 7840 5408 7848 5472
rect 7912 5408 7928 5472
rect 7992 5408 8008 5472
rect 8072 5408 8088 5472
rect 8152 5408 8160 5472
rect 7840 5407 8160 5408
rect 12437 5472 12757 5473
rect 12437 5408 12445 5472
rect 12509 5408 12525 5472
rect 12589 5408 12605 5472
rect 12669 5408 12685 5472
rect 12749 5408 12757 5472
rect 12437 5407 12757 5408
rect 1853 5402 1919 5405
rect 0 5400 1919 5402
rect 0 5344 1858 5400
rect 1914 5344 1919 5400
rect 0 5342 1919 5344
rect 0 5312 480 5342
rect 1853 5339 1919 5342
rect 4102 5340 4108 5404
rect 4172 5402 4178 5404
rect 6453 5402 6519 5405
rect 4172 5400 6519 5402
rect 4172 5344 6458 5400
rect 6514 5344 6519 5400
rect 4172 5342 6519 5344
rect 4172 5340 4178 5342
rect 6453 5339 6519 5342
rect 13537 5402 13603 5405
rect 15520 5402 16000 5432
rect 13537 5400 16000 5402
rect 13537 5344 13542 5400
rect 13598 5344 16000 5400
rect 13537 5342 16000 5344
rect 13537 5339 13603 5342
rect 15520 5312 16000 5342
rect 3509 5266 3575 5269
rect 3734 5266 3740 5268
rect 3509 5264 3740 5266
rect 3509 5208 3514 5264
rect 3570 5208 3740 5264
rect 3509 5206 3740 5208
rect 3509 5203 3575 5206
rect 3734 5204 3740 5206
rect 3804 5266 3810 5268
rect 9029 5266 9095 5269
rect 3804 5264 9095 5266
rect 3804 5208 9034 5264
rect 9090 5208 9095 5264
rect 3804 5206 9095 5208
rect 3804 5204 3810 5206
rect 9029 5203 9095 5206
rect 10133 5266 10199 5269
rect 12198 5266 12204 5268
rect 10133 5264 12204 5266
rect 10133 5208 10138 5264
rect 10194 5208 12204 5264
rect 10133 5206 12204 5208
rect 10133 5203 10199 5206
rect 12198 5204 12204 5206
rect 12268 5266 12274 5268
rect 12433 5266 12499 5269
rect 12268 5264 12499 5266
rect 12268 5208 12438 5264
rect 12494 5208 12499 5264
rect 12268 5206 12499 5208
rect 12268 5204 12274 5206
rect 12433 5203 12499 5206
rect 2221 5130 2287 5133
rect 7281 5132 7347 5133
rect 2221 5128 6010 5130
rect 2221 5072 2226 5128
rect 2282 5072 6010 5128
rect 2221 5070 6010 5072
rect 2221 5067 2287 5070
rect 0 4994 480 5024
rect 4061 4994 4127 4997
rect 0 4992 4127 4994
rect 0 4936 4066 4992
rect 4122 4936 4127 4992
rect 0 4934 4127 4936
rect 5950 4994 6010 5070
rect 7230 5068 7236 5132
rect 7300 5130 7347 5132
rect 7741 5130 7807 5133
rect 7300 5128 7392 5130
rect 7342 5072 7392 5128
rect 7300 5070 7392 5072
rect 7468 5128 7807 5130
rect 7468 5072 7746 5128
rect 7802 5072 7807 5128
rect 7468 5070 7807 5072
rect 7300 5068 7347 5070
rect 7281 5067 7347 5068
rect 7468 4994 7528 5070
rect 7741 5067 7807 5070
rect 10225 5130 10291 5133
rect 13353 5130 13419 5133
rect 10225 5128 13419 5130
rect 10225 5072 10230 5128
rect 10286 5072 13358 5128
rect 13414 5072 13419 5128
rect 10225 5070 13419 5072
rect 10225 5067 10291 5070
rect 13353 5067 13419 5070
rect 5950 4934 7528 4994
rect 13629 4994 13695 4997
rect 15520 4994 16000 5024
rect 13629 4992 16000 4994
rect 13629 4936 13634 4992
rect 13690 4936 16000 4992
rect 13629 4934 16000 4936
rect 0 4904 480 4934
rect 4061 4931 4127 4934
rect 13629 4931 13695 4934
rect 5541 4928 5861 4929
rect 5541 4864 5549 4928
rect 5613 4864 5629 4928
rect 5693 4864 5709 4928
rect 5773 4864 5789 4928
rect 5853 4864 5861 4928
rect 5541 4863 5861 4864
rect 10138 4928 10458 4929
rect 10138 4864 10146 4928
rect 10210 4864 10226 4928
rect 10290 4864 10306 4928
rect 10370 4864 10386 4928
rect 10450 4864 10458 4928
rect 15520 4904 16000 4934
rect 10138 4863 10458 4864
rect 2589 4858 2655 4861
rect 5257 4858 5323 4861
rect 2589 4856 5323 4858
rect 2589 4800 2594 4856
rect 2650 4800 5262 4856
rect 5318 4800 5323 4856
rect 2589 4798 5323 4800
rect 2589 4795 2655 4798
rect 5257 4795 5323 4798
rect 2497 4722 2563 4725
rect 6729 4722 6795 4725
rect 8661 4722 8727 4725
rect 2497 4720 4124 4722
rect 2497 4664 2502 4720
rect 2558 4664 4124 4720
rect 2497 4662 4124 4664
rect 2497 4659 2563 4662
rect 0 4586 480 4616
rect 1209 4586 1275 4589
rect 0 4584 1275 4586
rect 0 4528 1214 4584
rect 1270 4528 1275 4584
rect 0 4526 1275 4528
rect 0 4496 480 4526
rect 1209 4523 1275 4526
rect 3141 4586 3207 4589
rect 3918 4586 3924 4588
rect 3141 4584 3924 4586
rect 3141 4528 3146 4584
rect 3202 4528 3924 4584
rect 3141 4526 3924 4528
rect 3141 4523 3207 4526
rect 3918 4524 3924 4526
rect 3988 4524 3994 4588
rect 3877 4450 3943 4453
rect 4064 4450 4124 4662
rect 6729 4720 8727 4722
rect 6729 4664 6734 4720
rect 6790 4664 8666 4720
rect 8722 4664 8727 4720
rect 6729 4662 8727 4664
rect 6729 4659 6795 4662
rect 8661 4659 8727 4662
rect 4470 4524 4476 4588
rect 4540 4586 4546 4588
rect 5809 4586 5875 4589
rect 12065 4586 12131 4589
rect 4540 4584 5875 4586
rect 4540 4528 5814 4584
rect 5870 4528 5875 4584
rect 4540 4526 5875 4528
rect 4540 4524 4546 4526
rect 5809 4523 5875 4526
rect 5950 4584 12131 4586
rect 5950 4528 12070 4584
rect 12126 4528 12131 4584
rect 5950 4526 12131 4528
rect 5950 4450 6010 4526
rect 12065 4523 12131 4526
rect 13721 4586 13787 4589
rect 15520 4586 16000 4616
rect 13721 4584 16000 4586
rect 13721 4528 13726 4584
rect 13782 4528 16000 4584
rect 13721 4526 16000 4528
rect 13721 4523 13787 4526
rect 15520 4496 16000 4526
rect 3877 4448 6010 4450
rect 3877 4392 3882 4448
rect 3938 4392 6010 4448
rect 3877 4390 6010 4392
rect 3877 4387 3943 4390
rect 3242 4384 3562 4385
rect 3242 4320 3250 4384
rect 3314 4320 3330 4384
rect 3394 4320 3410 4384
rect 3474 4320 3490 4384
rect 3554 4320 3562 4384
rect 3242 4319 3562 4320
rect 7840 4384 8160 4385
rect 7840 4320 7848 4384
rect 7912 4320 7928 4384
rect 7992 4320 8008 4384
rect 8072 4320 8088 4384
rect 8152 4320 8160 4384
rect 7840 4319 8160 4320
rect 12437 4384 12757 4385
rect 12437 4320 12445 4384
rect 12509 4320 12525 4384
rect 12589 4320 12605 4384
rect 12669 4320 12685 4384
rect 12749 4320 12757 4384
rect 12437 4319 12757 4320
rect 4337 4316 4403 4317
rect 4286 4314 4292 4316
rect 4210 4254 4292 4314
rect 4356 4314 4403 4316
rect 4356 4312 7666 4314
rect 4398 4256 7666 4312
rect 4286 4252 4292 4254
rect 4356 4254 7666 4256
rect 4356 4252 4403 4254
rect 4337 4251 4403 4252
rect 0 4178 480 4208
rect 3601 4178 3667 4181
rect 0 4176 3667 4178
rect 0 4120 3606 4176
rect 3662 4120 3667 4176
rect 0 4118 3667 4120
rect 7606 4178 7666 4254
rect 12249 4178 12315 4181
rect 7606 4176 12315 4178
rect 7606 4120 12254 4176
rect 12310 4120 12315 4176
rect 7606 4118 12315 4120
rect 0 4088 480 4118
rect 3601 4115 3667 4118
rect 12249 4115 12315 4118
rect 13537 4178 13603 4181
rect 15520 4178 16000 4208
rect 13537 4176 16000 4178
rect 13537 4120 13542 4176
rect 13598 4120 16000 4176
rect 13537 4118 16000 4120
rect 13537 4115 13603 4118
rect 15520 4088 16000 4118
rect 5257 4042 5323 4045
rect 9806 4042 9812 4044
rect 5257 4040 9812 4042
rect 5257 3984 5262 4040
rect 5318 3984 9812 4040
rect 5257 3982 9812 3984
rect 5257 3979 5323 3982
rect 9806 3980 9812 3982
rect 9876 3980 9882 4044
rect 2998 3844 3004 3908
rect 3068 3906 3074 3908
rect 3785 3906 3851 3909
rect 3969 3908 4035 3909
rect 3068 3904 3851 3906
rect 3068 3848 3790 3904
rect 3846 3848 3851 3904
rect 3068 3846 3851 3848
rect 3068 3844 3074 3846
rect 3785 3843 3851 3846
rect 3918 3844 3924 3908
rect 3988 3906 4035 3908
rect 3988 3904 4080 3906
rect 4030 3848 4080 3904
rect 3988 3846 4080 3848
rect 3988 3844 4035 3846
rect 3969 3843 4035 3844
rect 5541 3840 5861 3841
rect 0 3770 480 3800
rect 5541 3776 5549 3840
rect 5613 3776 5629 3840
rect 5693 3776 5709 3840
rect 5773 3776 5789 3840
rect 5853 3776 5861 3840
rect 5541 3775 5861 3776
rect 10138 3840 10458 3841
rect 10138 3776 10146 3840
rect 10210 3776 10226 3840
rect 10290 3776 10306 3840
rect 10370 3776 10386 3840
rect 10450 3776 10458 3840
rect 10138 3775 10458 3776
rect 1025 3770 1091 3773
rect 3969 3770 4035 3773
rect 9673 3772 9739 3773
rect 0 3768 1091 3770
rect 0 3712 1030 3768
rect 1086 3712 1091 3768
rect 0 3710 1091 3712
rect 0 3680 480 3710
rect 1025 3707 1091 3710
rect 1350 3768 4035 3770
rect 1350 3712 3974 3768
rect 4030 3712 4035 3768
rect 1350 3710 4035 3712
rect 0 3362 480 3392
rect 1350 3362 1410 3710
rect 3969 3707 4035 3710
rect 9622 3708 9628 3772
rect 9692 3770 9739 3772
rect 12341 3770 12407 3773
rect 15520 3770 16000 3800
rect 9692 3768 9784 3770
rect 9734 3712 9784 3768
rect 9692 3710 9784 3712
rect 12341 3768 16000 3770
rect 12341 3712 12346 3768
rect 12402 3712 16000 3768
rect 12341 3710 16000 3712
rect 9692 3708 9739 3710
rect 9673 3707 9739 3708
rect 12341 3707 12407 3710
rect 15520 3680 16000 3710
rect 1669 3634 1735 3637
rect 14641 3634 14707 3637
rect 1669 3632 14707 3634
rect 1669 3576 1674 3632
rect 1730 3576 14646 3632
rect 14702 3576 14707 3632
rect 1669 3574 14707 3576
rect 1669 3571 1735 3574
rect 14641 3571 14707 3574
rect 2129 3498 2195 3501
rect 5441 3498 5507 3501
rect 8937 3498 9003 3501
rect 2129 3496 3756 3498
rect 2129 3440 2134 3496
rect 2190 3440 3756 3496
rect 2129 3438 3756 3440
rect 2129 3435 2195 3438
rect 0 3302 1410 3362
rect 3696 3362 3756 3438
rect 5030 3496 9003 3498
rect 5030 3440 5446 3496
rect 5502 3440 8942 3496
rect 8998 3440 9003 3496
rect 5030 3438 9003 3440
rect 5030 3362 5090 3438
rect 5441 3435 5507 3438
rect 8937 3435 9003 3438
rect 11421 3498 11487 3501
rect 11421 3496 13922 3498
rect 11421 3440 11426 3496
rect 11482 3440 13922 3496
rect 11421 3438 13922 3440
rect 11421 3435 11487 3438
rect 3696 3302 5090 3362
rect 13862 3362 13922 3438
rect 15520 3362 16000 3392
rect 13862 3302 16000 3362
rect 0 3272 480 3302
rect 3242 3296 3562 3297
rect 3242 3232 3250 3296
rect 3314 3232 3330 3296
rect 3394 3232 3410 3296
rect 3474 3232 3490 3296
rect 3554 3232 3562 3296
rect 3242 3231 3562 3232
rect 7840 3296 8160 3297
rect 7840 3232 7848 3296
rect 7912 3232 7928 3296
rect 7992 3232 8008 3296
rect 8072 3232 8088 3296
rect 8152 3232 8160 3296
rect 7840 3231 8160 3232
rect 12437 3296 12757 3297
rect 12437 3232 12445 3296
rect 12509 3232 12525 3296
rect 12589 3232 12605 3296
rect 12669 3232 12685 3296
rect 12749 3232 12757 3296
rect 15520 3272 16000 3302
rect 12437 3231 12757 3232
rect 4521 3228 4587 3229
rect 4470 3164 4476 3228
rect 4540 3226 4587 3228
rect 4540 3224 4632 3226
rect 4582 3168 4632 3224
rect 4540 3166 4632 3168
rect 4540 3164 4587 3166
rect 4521 3163 4587 3164
rect 1393 3090 1459 3093
rect 5073 3090 5139 3093
rect 12985 3090 13051 3093
rect 1393 3088 4906 3090
rect 1393 3032 1398 3088
rect 1454 3032 4906 3088
rect 1393 3030 4906 3032
rect 1393 3027 1459 3030
rect 0 2954 480 2984
rect 4061 2954 4127 2957
rect 0 2952 4127 2954
rect 0 2896 4066 2952
rect 4122 2896 4127 2952
rect 0 2894 4127 2896
rect 4846 2954 4906 3030
rect 5073 3088 13051 3090
rect 5073 3032 5078 3088
rect 5134 3032 12990 3088
rect 13046 3032 13051 3088
rect 5073 3030 13051 3032
rect 5073 3027 5139 3030
rect 12985 3027 13051 3030
rect 8753 2954 8819 2957
rect 9673 2956 9739 2957
rect 4846 2952 8819 2954
rect 4846 2896 8758 2952
rect 8814 2896 8819 2952
rect 4846 2894 8819 2896
rect 0 2864 480 2894
rect 4061 2891 4127 2894
rect 8753 2891 8819 2894
rect 9622 2892 9628 2956
rect 9692 2954 9739 2956
rect 10961 2954 11027 2957
rect 15520 2954 16000 2984
rect 9692 2952 9784 2954
rect 9734 2896 9784 2952
rect 9692 2894 9784 2896
rect 10961 2952 16000 2954
rect 10961 2896 10966 2952
rect 11022 2896 16000 2952
rect 10961 2894 16000 2896
rect 9692 2892 9739 2894
rect 9673 2891 9739 2892
rect 10961 2891 11027 2894
rect 15520 2864 16000 2894
rect 4102 2756 4108 2820
rect 4172 2818 4178 2820
rect 4889 2818 4955 2821
rect 11329 2820 11395 2821
rect 4172 2816 4955 2818
rect 4172 2760 4894 2816
rect 4950 2760 4955 2816
rect 4172 2758 4955 2760
rect 4172 2756 4178 2758
rect 4889 2755 4955 2758
rect 11278 2756 11284 2820
rect 11348 2818 11395 2820
rect 11348 2816 11440 2818
rect 11390 2760 11440 2816
rect 11348 2758 11440 2760
rect 11348 2756 11395 2758
rect 11329 2755 11395 2756
rect 5541 2752 5861 2753
rect 5541 2688 5549 2752
rect 5613 2688 5629 2752
rect 5693 2688 5709 2752
rect 5773 2688 5789 2752
rect 5853 2688 5861 2752
rect 5541 2687 5861 2688
rect 10138 2752 10458 2753
rect 10138 2688 10146 2752
rect 10210 2688 10226 2752
rect 10290 2688 10306 2752
rect 10370 2688 10386 2752
rect 10450 2688 10458 2752
rect 10138 2687 10458 2688
rect 1761 2682 1827 2685
rect 1761 2680 3250 2682
rect 1761 2624 1766 2680
rect 1822 2624 3250 2680
rect 1761 2622 3250 2624
rect 1761 2619 1827 2622
rect 0 2546 480 2576
rect 2957 2546 3023 2549
rect 0 2544 3023 2546
rect 0 2488 2962 2544
rect 3018 2488 3023 2544
rect 0 2486 3023 2488
rect 3190 2546 3250 2622
rect 3693 2546 3759 2549
rect 4613 2546 4679 2549
rect 3190 2544 4679 2546
rect 3190 2488 3698 2544
rect 3754 2488 4618 2544
rect 4674 2488 4679 2544
rect 3190 2486 4679 2488
rect 0 2456 480 2486
rect 2957 2483 3023 2486
rect 3693 2483 3759 2486
rect 4613 2483 4679 2486
rect 12157 2546 12223 2549
rect 15520 2546 16000 2576
rect 12157 2544 16000 2546
rect 12157 2488 12162 2544
rect 12218 2488 16000 2544
rect 12157 2486 16000 2488
rect 12157 2483 12223 2486
rect 15520 2456 16000 2486
rect 2865 2410 2931 2413
rect 3918 2410 3924 2412
rect 2865 2408 3924 2410
rect 2865 2352 2870 2408
rect 2926 2352 3924 2408
rect 2865 2350 3924 2352
rect 2865 2347 2931 2350
rect 3918 2348 3924 2350
rect 3988 2410 3994 2412
rect 4613 2410 4679 2413
rect 3988 2408 4679 2410
rect 3988 2352 4618 2408
rect 4674 2352 4679 2408
rect 3988 2350 4679 2352
rect 3988 2348 3994 2350
rect 4613 2347 4679 2350
rect 11053 2410 11119 2413
rect 11053 2408 13922 2410
rect 11053 2352 11058 2408
rect 11114 2352 13922 2408
rect 11053 2350 13922 2352
rect 11053 2347 11119 2350
rect 3242 2208 3562 2209
rect 0 2138 480 2168
rect 3242 2144 3250 2208
rect 3314 2144 3330 2208
rect 3394 2144 3410 2208
rect 3474 2144 3490 2208
rect 3554 2144 3562 2208
rect 3242 2143 3562 2144
rect 7840 2208 8160 2209
rect 7840 2144 7848 2208
rect 7912 2144 7928 2208
rect 7992 2144 8008 2208
rect 8072 2144 8088 2208
rect 8152 2144 8160 2208
rect 7840 2143 8160 2144
rect 12437 2208 12757 2209
rect 12437 2144 12445 2208
rect 12509 2144 12525 2208
rect 12589 2144 12605 2208
rect 12669 2144 12685 2208
rect 12749 2144 12757 2208
rect 12437 2143 12757 2144
rect 3049 2138 3115 2141
rect 0 2136 3115 2138
rect 0 2080 3054 2136
rect 3110 2080 3115 2136
rect 0 2078 3115 2080
rect 13862 2138 13922 2350
rect 15520 2138 16000 2168
rect 13862 2078 16000 2138
rect 0 2048 480 2078
rect 3049 2075 3115 2078
rect 15520 2048 16000 2078
rect 0 1730 480 1760
rect 2037 1730 2103 1733
rect 0 1728 2103 1730
rect 0 1672 2042 1728
rect 2098 1672 2103 1728
rect 0 1670 2103 1672
rect 0 1640 480 1670
rect 2037 1667 2103 1670
rect 11421 1730 11487 1733
rect 15520 1730 16000 1760
rect 11421 1728 16000 1730
rect 11421 1672 11426 1728
rect 11482 1672 16000 1728
rect 11421 1670 16000 1672
rect 11421 1667 11487 1670
rect 15520 1640 16000 1670
rect 0 1322 480 1352
rect 1577 1322 1643 1325
rect 0 1320 1643 1322
rect 0 1264 1582 1320
rect 1638 1264 1643 1320
rect 0 1262 1643 1264
rect 0 1232 480 1262
rect 1577 1259 1643 1262
rect 11513 1322 11579 1325
rect 15520 1322 16000 1352
rect 11513 1320 16000 1322
rect 11513 1264 11518 1320
rect 11574 1264 16000 1320
rect 11513 1262 16000 1264
rect 11513 1259 11579 1262
rect 15520 1232 16000 1262
rect 0 914 480 944
rect 2313 914 2379 917
rect 0 912 2379 914
rect 0 856 2318 912
rect 2374 856 2379 912
rect 0 854 2379 856
rect 0 824 480 854
rect 2313 851 2379 854
rect 11605 914 11671 917
rect 15520 914 16000 944
rect 11605 912 16000 914
rect 11605 856 11610 912
rect 11666 856 16000 912
rect 11605 854 16000 856
rect 11605 851 11671 854
rect 15520 824 16000 854
rect 0 506 480 536
rect 2773 506 2839 509
rect 0 504 2839 506
rect 0 448 2778 504
rect 2834 448 2839 504
rect 0 446 2839 448
rect 0 416 480 446
rect 2773 443 2839 446
rect 11145 506 11211 509
rect 15520 506 16000 536
rect 11145 504 16000 506
rect 11145 448 11150 504
rect 11206 448 16000 504
rect 11145 446 16000 448
rect 11145 443 11211 446
rect 15520 416 16000 446
rect 0 234 480 264
rect 2865 234 2931 237
rect 0 232 2931 234
rect 0 176 2870 232
rect 2926 176 2931 232
rect 0 174 2931 176
rect 0 144 480 174
rect 2865 171 2931 174
rect 12617 234 12683 237
rect 15520 234 16000 264
rect 12617 232 16000 234
rect 12617 176 12622 232
rect 12678 176 16000 232
rect 12617 174 16000 176
rect 12617 171 12683 174
rect 15520 144 16000 174
<< via3 >>
rect 5549 13628 5613 13632
rect 5549 13572 5553 13628
rect 5553 13572 5609 13628
rect 5609 13572 5613 13628
rect 5549 13568 5613 13572
rect 5629 13628 5693 13632
rect 5629 13572 5633 13628
rect 5633 13572 5689 13628
rect 5689 13572 5693 13628
rect 5629 13568 5693 13572
rect 5709 13628 5773 13632
rect 5709 13572 5713 13628
rect 5713 13572 5769 13628
rect 5769 13572 5773 13628
rect 5709 13568 5773 13572
rect 5789 13628 5853 13632
rect 5789 13572 5793 13628
rect 5793 13572 5849 13628
rect 5849 13572 5853 13628
rect 5789 13568 5853 13572
rect 10146 13628 10210 13632
rect 10146 13572 10150 13628
rect 10150 13572 10206 13628
rect 10206 13572 10210 13628
rect 10146 13568 10210 13572
rect 10226 13628 10290 13632
rect 10226 13572 10230 13628
rect 10230 13572 10286 13628
rect 10286 13572 10290 13628
rect 10226 13568 10290 13572
rect 10306 13628 10370 13632
rect 10306 13572 10310 13628
rect 10310 13572 10366 13628
rect 10366 13572 10370 13628
rect 10306 13568 10370 13572
rect 10386 13628 10450 13632
rect 10386 13572 10390 13628
rect 10390 13572 10446 13628
rect 10446 13572 10450 13628
rect 10386 13568 10450 13572
rect 3250 13084 3314 13088
rect 3250 13028 3254 13084
rect 3254 13028 3310 13084
rect 3310 13028 3314 13084
rect 3250 13024 3314 13028
rect 3330 13084 3394 13088
rect 3330 13028 3334 13084
rect 3334 13028 3390 13084
rect 3390 13028 3394 13084
rect 3330 13024 3394 13028
rect 3410 13084 3474 13088
rect 3410 13028 3414 13084
rect 3414 13028 3470 13084
rect 3470 13028 3474 13084
rect 3410 13024 3474 13028
rect 3490 13084 3554 13088
rect 3490 13028 3494 13084
rect 3494 13028 3550 13084
rect 3550 13028 3554 13084
rect 3490 13024 3554 13028
rect 7848 13084 7912 13088
rect 7848 13028 7852 13084
rect 7852 13028 7908 13084
rect 7908 13028 7912 13084
rect 7848 13024 7912 13028
rect 7928 13084 7992 13088
rect 7928 13028 7932 13084
rect 7932 13028 7988 13084
rect 7988 13028 7992 13084
rect 7928 13024 7992 13028
rect 8008 13084 8072 13088
rect 8008 13028 8012 13084
rect 8012 13028 8068 13084
rect 8068 13028 8072 13084
rect 8008 13024 8072 13028
rect 8088 13084 8152 13088
rect 8088 13028 8092 13084
rect 8092 13028 8148 13084
rect 8148 13028 8152 13084
rect 8088 13024 8152 13028
rect 12445 13084 12509 13088
rect 12445 13028 12449 13084
rect 12449 13028 12505 13084
rect 12505 13028 12509 13084
rect 12445 13024 12509 13028
rect 12525 13084 12589 13088
rect 12525 13028 12529 13084
rect 12529 13028 12585 13084
rect 12585 13028 12589 13084
rect 12525 13024 12589 13028
rect 12605 13084 12669 13088
rect 12605 13028 12609 13084
rect 12609 13028 12665 13084
rect 12665 13028 12669 13084
rect 12605 13024 12669 13028
rect 12685 13084 12749 13088
rect 12685 13028 12689 13084
rect 12689 13028 12745 13084
rect 12745 13028 12749 13084
rect 12685 13024 12749 13028
rect 9812 12880 9876 12884
rect 9812 12824 9826 12880
rect 9826 12824 9876 12880
rect 9812 12820 9876 12824
rect 5549 12540 5613 12544
rect 5549 12484 5553 12540
rect 5553 12484 5609 12540
rect 5609 12484 5613 12540
rect 5549 12480 5613 12484
rect 5629 12540 5693 12544
rect 5629 12484 5633 12540
rect 5633 12484 5689 12540
rect 5689 12484 5693 12540
rect 5629 12480 5693 12484
rect 5709 12540 5773 12544
rect 5709 12484 5713 12540
rect 5713 12484 5769 12540
rect 5769 12484 5773 12540
rect 5709 12480 5773 12484
rect 5789 12540 5853 12544
rect 5789 12484 5793 12540
rect 5793 12484 5849 12540
rect 5849 12484 5853 12540
rect 5789 12480 5853 12484
rect 10146 12540 10210 12544
rect 10146 12484 10150 12540
rect 10150 12484 10206 12540
rect 10206 12484 10210 12540
rect 10146 12480 10210 12484
rect 10226 12540 10290 12544
rect 10226 12484 10230 12540
rect 10230 12484 10286 12540
rect 10286 12484 10290 12540
rect 10226 12480 10290 12484
rect 10306 12540 10370 12544
rect 10306 12484 10310 12540
rect 10310 12484 10366 12540
rect 10366 12484 10370 12540
rect 10306 12480 10370 12484
rect 10386 12540 10450 12544
rect 10386 12484 10390 12540
rect 10390 12484 10446 12540
rect 10446 12484 10450 12540
rect 10386 12480 10450 12484
rect 2820 12412 2884 12476
rect 3250 11996 3314 12000
rect 3250 11940 3254 11996
rect 3254 11940 3310 11996
rect 3310 11940 3314 11996
rect 3250 11936 3314 11940
rect 3330 11996 3394 12000
rect 3330 11940 3334 11996
rect 3334 11940 3390 11996
rect 3390 11940 3394 11996
rect 3330 11936 3394 11940
rect 3410 11996 3474 12000
rect 3410 11940 3414 11996
rect 3414 11940 3470 11996
rect 3470 11940 3474 11996
rect 3410 11936 3474 11940
rect 3490 11996 3554 12000
rect 3490 11940 3494 11996
rect 3494 11940 3550 11996
rect 3550 11940 3554 11996
rect 3490 11936 3554 11940
rect 7848 11996 7912 12000
rect 7848 11940 7852 11996
rect 7852 11940 7908 11996
rect 7908 11940 7912 11996
rect 7848 11936 7912 11940
rect 7928 11996 7992 12000
rect 7928 11940 7932 11996
rect 7932 11940 7988 11996
rect 7988 11940 7992 11996
rect 7928 11936 7992 11940
rect 8008 11996 8072 12000
rect 8008 11940 8012 11996
rect 8012 11940 8068 11996
rect 8068 11940 8072 11996
rect 8008 11936 8072 11940
rect 8088 11996 8152 12000
rect 8088 11940 8092 11996
rect 8092 11940 8148 11996
rect 8148 11940 8152 11996
rect 8088 11936 8152 11940
rect 12445 11996 12509 12000
rect 12445 11940 12449 11996
rect 12449 11940 12505 11996
rect 12505 11940 12509 11996
rect 12445 11936 12509 11940
rect 12525 11996 12589 12000
rect 12525 11940 12529 11996
rect 12529 11940 12585 11996
rect 12585 11940 12589 11996
rect 12525 11936 12589 11940
rect 12605 11996 12669 12000
rect 12605 11940 12609 11996
rect 12609 11940 12665 11996
rect 12665 11940 12669 11996
rect 12605 11936 12669 11940
rect 12685 11996 12749 12000
rect 12685 11940 12689 11996
rect 12689 11940 12745 11996
rect 12745 11940 12749 11996
rect 12685 11936 12749 11940
rect 5549 11452 5613 11456
rect 5549 11396 5553 11452
rect 5553 11396 5609 11452
rect 5609 11396 5613 11452
rect 5549 11392 5613 11396
rect 5629 11452 5693 11456
rect 5629 11396 5633 11452
rect 5633 11396 5689 11452
rect 5689 11396 5693 11452
rect 5629 11392 5693 11396
rect 5709 11452 5773 11456
rect 5709 11396 5713 11452
rect 5713 11396 5769 11452
rect 5769 11396 5773 11452
rect 5709 11392 5773 11396
rect 5789 11452 5853 11456
rect 5789 11396 5793 11452
rect 5793 11396 5849 11452
rect 5849 11396 5853 11452
rect 5789 11392 5853 11396
rect 10146 11452 10210 11456
rect 10146 11396 10150 11452
rect 10150 11396 10206 11452
rect 10206 11396 10210 11452
rect 10146 11392 10210 11396
rect 10226 11452 10290 11456
rect 10226 11396 10230 11452
rect 10230 11396 10286 11452
rect 10286 11396 10290 11452
rect 10226 11392 10290 11396
rect 10306 11452 10370 11456
rect 10306 11396 10310 11452
rect 10310 11396 10366 11452
rect 10366 11396 10370 11452
rect 10306 11392 10370 11396
rect 10386 11452 10450 11456
rect 10386 11396 10390 11452
rect 10390 11396 10446 11452
rect 10446 11396 10450 11452
rect 10386 11392 10450 11396
rect 3740 11188 3804 11252
rect 4108 11052 4172 11116
rect 3924 10976 3988 10980
rect 3924 10920 3974 10976
rect 3974 10920 3988 10976
rect 3924 10916 3988 10920
rect 3250 10908 3314 10912
rect 3250 10852 3254 10908
rect 3254 10852 3310 10908
rect 3310 10852 3314 10908
rect 3250 10848 3314 10852
rect 3330 10908 3394 10912
rect 3330 10852 3334 10908
rect 3334 10852 3390 10908
rect 3390 10852 3394 10908
rect 3330 10848 3394 10852
rect 3410 10908 3474 10912
rect 3410 10852 3414 10908
rect 3414 10852 3470 10908
rect 3470 10852 3474 10908
rect 3410 10848 3474 10852
rect 3490 10908 3554 10912
rect 3490 10852 3494 10908
rect 3494 10852 3550 10908
rect 3550 10852 3554 10908
rect 3490 10848 3554 10852
rect 7848 10908 7912 10912
rect 7848 10852 7852 10908
rect 7852 10852 7908 10908
rect 7908 10852 7912 10908
rect 7848 10848 7912 10852
rect 7928 10908 7992 10912
rect 7928 10852 7932 10908
rect 7932 10852 7988 10908
rect 7988 10852 7992 10908
rect 7928 10848 7992 10852
rect 8008 10908 8072 10912
rect 8008 10852 8012 10908
rect 8012 10852 8068 10908
rect 8068 10852 8072 10908
rect 8008 10848 8072 10852
rect 8088 10908 8152 10912
rect 8088 10852 8092 10908
rect 8092 10852 8148 10908
rect 8148 10852 8152 10908
rect 8088 10848 8152 10852
rect 12445 10908 12509 10912
rect 12445 10852 12449 10908
rect 12449 10852 12505 10908
rect 12505 10852 12509 10908
rect 12445 10848 12509 10852
rect 12525 10908 12589 10912
rect 12525 10852 12529 10908
rect 12529 10852 12585 10908
rect 12585 10852 12589 10908
rect 12525 10848 12589 10852
rect 12605 10908 12669 10912
rect 12605 10852 12609 10908
rect 12609 10852 12665 10908
rect 12665 10852 12669 10908
rect 12605 10848 12669 10852
rect 12685 10908 12749 10912
rect 12685 10852 12689 10908
rect 12689 10852 12745 10908
rect 12745 10852 12749 10908
rect 12685 10848 12749 10852
rect 5549 10364 5613 10368
rect 5549 10308 5553 10364
rect 5553 10308 5609 10364
rect 5609 10308 5613 10364
rect 5549 10304 5613 10308
rect 5629 10364 5693 10368
rect 5629 10308 5633 10364
rect 5633 10308 5689 10364
rect 5689 10308 5693 10364
rect 5629 10304 5693 10308
rect 5709 10364 5773 10368
rect 5709 10308 5713 10364
rect 5713 10308 5769 10364
rect 5769 10308 5773 10364
rect 5709 10304 5773 10308
rect 5789 10364 5853 10368
rect 5789 10308 5793 10364
rect 5793 10308 5849 10364
rect 5849 10308 5853 10364
rect 5789 10304 5853 10308
rect 10146 10364 10210 10368
rect 10146 10308 10150 10364
rect 10150 10308 10206 10364
rect 10206 10308 10210 10364
rect 10146 10304 10210 10308
rect 10226 10364 10290 10368
rect 10226 10308 10230 10364
rect 10230 10308 10286 10364
rect 10286 10308 10290 10364
rect 10226 10304 10290 10308
rect 10306 10364 10370 10368
rect 10306 10308 10310 10364
rect 10310 10308 10366 10364
rect 10366 10308 10370 10364
rect 10306 10304 10370 10308
rect 10386 10364 10450 10368
rect 10386 10308 10390 10364
rect 10390 10308 10446 10364
rect 10446 10308 10450 10364
rect 10386 10304 10450 10308
rect 3004 10296 3068 10300
rect 3004 10240 3018 10296
rect 3018 10240 3068 10296
rect 3004 10236 3068 10240
rect 12204 9964 12268 10028
rect 3250 9820 3314 9824
rect 3250 9764 3254 9820
rect 3254 9764 3310 9820
rect 3310 9764 3314 9820
rect 3250 9760 3314 9764
rect 3330 9820 3394 9824
rect 3330 9764 3334 9820
rect 3334 9764 3390 9820
rect 3390 9764 3394 9820
rect 3330 9760 3394 9764
rect 3410 9820 3474 9824
rect 3410 9764 3414 9820
rect 3414 9764 3470 9820
rect 3470 9764 3474 9820
rect 3410 9760 3474 9764
rect 3490 9820 3554 9824
rect 3490 9764 3494 9820
rect 3494 9764 3550 9820
rect 3550 9764 3554 9820
rect 3490 9760 3554 9764
rect 7848 9820 7912 9824
rect 7848 9764 7852 9820
rect 7852 9764 7908 9820
rect 7908 9764 7912 9820
rect 7848 9760 7912 9764
rect 7928 9820 7992 9824
rect 7928 9764 7932 9820
rect 7932 9764 7988 9820
rect 7988 9764 7992 9820
rect 7928 9760 7992 9764
rect 8008 9820 8072 9824
rect 8008 9764 8012 9820
rect 8012 9764 8068 9820
rect 8068 9764 8072 9820
rect 8008 9760 8072 9764
rect 8088 9820 8152 9824
rect 8088 9764 8092 9820
rect 8092 9764 8148 9820
rect 8148 9764 8152 9820
rect 8088 9760 8152 9764
rect 12445 9820 12509 9824
rect 12445 9764 12449 9820
rect 12449 9764 12505 9820
rect 12505 9764 12509 9820
rect 12445 9760 12509 9764
rect 12525 9820 12589 9824
rect 12525 9764 12529 9820
rect 12529 9764 12585 9820
rect 12585 9764 12589 9820
rect 12525 9760 12589 9764
rect 12605 9820 12669 9824
rect 12605 9764 12609 9820
rect 12609 9764 12665 9820
rect 12665 9764 12669 9820
rect 12605 9760 12669 9764
rect 12685 9820 12749 9824
rect 12685 9764 12689 9820
rect 12689 9764 12745 9820
rect 12745 9764 12749 9820
rect 12685 9760 12749 9764
rect 4476 9556 4540 9620
rect 2820 9284 2884 9348
rect 5549 9276 5613 9280
rect 5549 9220 5553 9276
rect 5553 9220 5609 9276
rect 5609 9220 5613 9276
rect 5549 9216 5613 9220
rect 5629 9276 5693 9280
rect 5629 9220 5633 9276
rect 5633 9220 5689 9276
rect 5689 9220 5693 9276
rect 5629 9216 5693 9220
rect 5709 9276 5773 9280
rect 5709 9220 5713 9276
rect 5713 9220 5769 9276
rect 5769 9220 5773 9276
rect 5709 9216 5773 9220
rect 5789 9276 5853 9280
rect 5789 9220 5793 9276
rect 5793 9220 5849 9276
rect 5849 9220 5853 9276
rect 5789 9216 5853 9220
rect 10146 9276 10210 9280
rect 10146 9220 10150 9276
rect 10150 9220 10206 9276
rect 10206 9220 10210 9276
rect 10146 9216 10210 9220
rect 10226 9276 10290 9280
rect 10226 9220 10230 9276
rect 10230 9220 10286 9276
rect 10286 9220 10290 9276
rect 10226 9216 10290 9220
rect 10306 9276 10370 9280
rect 10306 9220 10310 9276
rect 10310 9220 10366 9276
rect 10366 9220 10370 9276
rect 10306 9216 10370 9220
rect 10386 9276 10450 9280
rect 10386 9220 10390 9276
rect 10390 9220 10446 9276
rect 10446 9220 10450 9276
rect 10386 9216 10450 9220
rect 4292 8876 4356 8940
rect 3250 8732 3314 8736
rect 3250 8676 3254 8732
rect 3254 8676 3310 8732
rect 3310 8676 3314 8732
rect 3250 8672 3314 8676
rect 3330 8732 3394 8736
rect 3330 8676 3334 8732
rect 3334 8676 3390 8732
rect 3390 8676 3394 8732
rect 3330 8672 3394 8676
rect 3410 8732 3474 8736
rect 3410 8676 3414 8732
rect 3414 8676 3470 8732
rect 3470 8676 3474 8732
rect 3410 8672 3474 8676
rect 3490 8732 3554 8736
rect 3490 8676 3494 8732
rect 3494 8676 3550 8732
rect 3550 8676 3554 8732
rect 3490 8672 3554 8676
rect 7848 8732 7912 8736
rect 7848 8676 7852 8732
rect 7852 8676 7908 8732
rect 7908 8676 7912 8732
rect 7848 8672 7912 8676
rect 7928 8732 7992 8736
rect 7928 8676 7932 8732
rect 7932 8676 7988 8732
rect 7988 8676 7992 8732
rect 7928 8672 7992 8676
rect 8008 8732 8072 8736
rect 8008 8676 8012 8732
rect 8012 8676 8068 8732
rect 8068 8676 8072 8732
rect 8008 8672 8072 8676
rect 8088 8732 8152 8736
rect 8088 8676 8092 8732
rect 8092 8676 8148 8732
rect 8148 8676 8152 8732
rect 8088 8672 8152 8676
rect 12445 8732 12509 8736
rect 12445 8676 12449 8732
rect 12449 8676 12505 8732
rect 12505 8676 12509 8732
rect 12445 8672 12509 8676
rect 12525 8732 12589 8736
rect 12525 8676 12529 8732
rect 12529 8676 12585 8732
rect 12585 8676 12589 8732
rect 12525 8672 12589 8676
rect 12605 8732 12669 8736
rect 12605 8676 12609 8732
rect 12609 8676 12665 8732
rect 12665 8676 12669 8732
rect 12605 8672 12669 8676
rect 12685 8732 12749 8736
rect 12685 8676 12689 8732
rect 12689 8676 12745 8732
rect 12745 8676 12749 8732
rect 12685 8672 12749 8676
rect 11284 8664 11348 8668
rect 11284 8608 11334 8664
rect 11334 8608 11348 8664
rect 11284 8604 11348 8608
rect 5549 8188 5613 8192
rect 5549 8132 5553 8188
rect 5553 8132 5609 8188
rect 5609 8132 5613 8188
rect 5549 8128 5613 8132
rect 5629 8188 5693 8192
rect 5629 8132 5633 8188
rect 5633 8132 5689 8188
rect 5689 8132 5693 8188
rect 5629 8128 5693 8132
rect 5709 8188 5773 8192
rect 5709 8132 5713 8188
rect 5713 8132 5769 8188
rect 5769 8132 5773 8188
rect 5709 8128 5773 8132
rect 5789 8188 5853 8192
rect 5789 8132 5793 8188
rect 5793 8132 5849 8188
rect 5849 8132 5853 8188
rect 5789 8128 5853 8132
rect 10146 8188 10210 8192
rect 10146 8132 10150 8188
rect 10150 8132 10206 8188
rect 10206 8132 10210 8188
rect 10146 8128 10210 8132
rect 10226 8188 10290 8192
rect 10226 8132 10230 8188
rect 10230 8132 10286 8188
rect 10286 8132 10290 8188
rect 10226 8128 10290 8132
rect 10306 8188 10370 8192
rect 10306 8132 10310 8188
rect 10310 8132 10366 8188
rect 10366 8132 10370 8188
rect 10306 8128 10370 8132
rect 10386 8188 10450 8192
rect 10386 8132 10390 8188
rect 10390 8132 10446 8188
rect 10446 8132 10450 8188
rect 10386 8128 10450 8132
rect 11836 8120 11900 8124
rect 11836 8064 11850 8120
rect 11850 8064 11900 8120
rect 11836 8060 11900 8064
rect 3250 7644 3314 7648
rect 3250 7588 3254 7644
rect 3254 7588 3310 7644
rect 3310 7588 3314 7644
rect 3250 7584 3314 7588
rect 3330 7644 3394 7648
rect 3330 7588 3334 7644
rect 3334 7588 3390 7644
rect 3390 7588 3394 7644
rect 3330 7584 3394 7588
rect 3410 7644 3474 7648
rect 3410 7588 3414 7644
rect 3414 7588 3470 7644
rect 3470 7588 3474 7644
rect 3410 7584 3474 7588
rect 3490 7644 3554 7648
rect 3490 7588 3494 7644
rect 3494 7588 3550 7644
rect 3550 7588 3554 7644
rect 3490 7584 3554 7588
rect 7848 7644 7912 7648
rect 7848 7588 7852 7644
rect 7852 7588 7908 7644
rect 7908 7588 7912 7644
rect 7848 7584 7912 7588
rect 7928 7644 7992 7648
rect 7928 7588 7932 7644
rect 7932 7588 7988 7644
rect 7988 7588 7992 7644
rect 7928 7584 7992 7588
rect 8008 7644 8072 7648
rect 8008 7588 8012 7644
rect 8012 7588 8068 7644
rect 8068 7588 8072 7644
rect 8008 7584 8072 7588
rect 8088 7644 8152 7648
rect 8088 7588 8092 7644
rect 8092 7588 8148 7644
rect 8148 7588 8152 7644
rect 8088 7584 8152 7588
rect 12445 7644 12509 7648
rect 12445 7588 12449 7644
rect 12449 7588 12505 7644
rect 12505 7588 12509 7644
rect 12445 7584 12509 7588
rect 12525 7644 12589 7648
rect 12525 7588 12529 7644
rect 12529 7588 12585 7644
rect 12585 7588 12589 7644
rect 12525 7584 12589 7588
rect 12605 7644 12669 7648
rect 12605 7588 12609 7644
rect 12609 7588 12665 7644
rect 12665 7588 12669 7644
rect 12605 7584 12669 7588
rect 12685 7644 12749 7648
rect 12685 7588 12689 7644
rect 12689 7588 12745 7644
rect 12745 7588 12749 7644
rect 12685 7584 12749 7588
rect 11836 7168 11900 7172
rect 11836 7112 11850 7168
rect 11850 7112 11900 7168
rect 11836 7108 11900 7112
rect 5549 7100 5613 7104
rect 5549 7044 5553 7100
rect 5553 7044 5609 7100
rect 5609 7044 5613 7100
rect 5549 7040 5613 7044
rect 5629 7100 5693 7104
rect 5629 7044 5633 7100
rect 5633 7044 5689 7100
rect 5689 7044 5693 7100
rect 5629 7040 5693 7044
rect 5709 7100 5773 7104
rect 5709 7044 5713 7100
rect 5713 7044 5769 7100
rect 5769 7044 5773 7100
rect 5709 7040 5773 7044
rect 5789 7100 5853 7104
rect 5789 7044 5793 7100
rect 5793 7044 5849 7100
rect 5849 7044 5853 7100
rect 5789 7040 5853 7044
rect 10146 7100 10210 7104
rect 10146 7044 10150 7100
rect 10150 7044 10206 7100
rect 10206 7044 10210 7100
rect 10146 7040 10210 7044
rect 10226 7100 10290 7104
rect 10226 7044 10230 7100
rect 10230 7044 10286 7100
rect 10286 7044 10290 7100
rect 10226 7040 10290 7044
rect 10306 7100 10370 7104
rect 10306 7044 10310 7100
rect 10310 7044 10366 7100
rect 10366 7044 10370 7100
rect 10306 7040 10370 7044
rect 10386 7100 10450 7104
rect 10386 7044 10390 7100
rect 10390 7044 10446 7100
rect 10446 7044 10450 7100
rect 10386 7040 10450 7044
rect 7236 6700 7300 6764
rect 3250 6556 3314 6560
rect 3250 6500 3254 6556
rect 3254 6500 3310 6556
rect 3310 6500 3314 6556
rect 3250 6496 3314 6500
rect 3330 6556 3394 6560
rect 3330 6500 3334 6556
rect 3334 6500 3390 6556
rect 3390 6500 3394 6556
rect 3330 6496 3394 6500
rect 3410 6556 3474 6560
rect 3410 6500 3414 6556
rect 3414 6500 3470 6556
rect 3470 6500 3474 6556
rect 3410 6496 3474 6500
rect 3490 6556 3554 6560
rect 3490 6500 3494 6556
rect 3494 6500 3550 6556
rect 3550 6500 3554 6556
rect 3490 6496 3554 6500
rect 7848 6556 7912 6560
rect 7848 6500 7852 6556
rect 7852 6500 7908 6556
rect 7908 6500 7912 6556
rect 7848 6496 7912 6500
rect 7928 6556 7992 6560
rect 7928 6500 7932 6556
rect 7932 6500 7988 6556
rect 7988 6500 7992 6556
rect 7928 6496 7992 6500
rect 8008 6556 8072 6560
rect 8008 6500 8012 6556
rect 8012 6500 8068 6556
rect 8068 6500 8072 6556
rect 8008 6496 8072 6500
rect 8088 6556 8152 6560
rect 8088 6500 8092 6556
rect 8092 6500 8148 6556
rect 8148 6500 8152 6556
rect 8088 6496 8152 6500
rect 12445 6556 12509 6560
rect 12445 6500 12449 6556
rect 12449 6500 12505 6556
rect 12505 6500 12509 6556
rect 12445 6496 12509 6500
rect 12525 6556 12589 6560
rect 12525 6500 12529 6556
rect 12529 6500 12585 6556
rect 12585 6500 12589 6556
rect 12525 6496 12589 6500
rect 12605 6556 12669 6560
rect 12605 6500 12609 6556
rect 12609 6500 12665 6556
rect 12665 6500 12669 6556
rect 12605 6496 12669 6500
rect 12685 6556 12749 6560
rect 12685 6500 12689 6556
rect 12689 6500 12745 6556
rect 12745 6500 12749 6556
rect 12685 6496 12749 6500
rect 5549 6012 5613 6016
rect 5549 5956 5553 6012
rect 5553 5956 5609 6012
rect 5609 5956 5613 6012
rect 5549 5952 5613 5956
rect 5629 6012 5693 6016
rect 5629 5956 5633 6012
rect 5633 5956 5689 6012
rect 5689 5956 5693 6012
rect 5629 5952 5693 5956
rect 5709 6012 5773 6016
rect 5709 5956 5713 6012
rect 5713 5956 5769 6012
rect 5769 5956 5773 6012
rect 5709 5952 5773 5956
rect 5789 6012 5853 6016
rect 5789 5956 5793 6012
rect 5793 5956 5849 6012
rect 5849 5956 5853 6012
rect 5789 5952 5853 5956
rect 10146 6012 10210 6016
rect 10146 5956 10150 6012
rect 10150 5956 10206 6012
rect 10206 5956 10210 6012
rect 10146 5952 10210 5956
rect 10226 6012 10290 6016
rect 10226 5956 10230 6012
rect 10230 5956 10286 6012
rect 10286 5956 10290 6012
rect 10226 5952 10290 5956
rect 10306 6012 10370 6016
rect 10306 5956 10310 6012
rect 10310 5956 10366 6012
rect 10366 5956 10370 6012
rect 10306 5952 10370 5956
rect 10386 6012 10450 6016
rect 10386 5956 10390 6012
rect 10390 5956 10446 6012
rect 10446 5956 10450 6012
rect 10386 5952 10450 5956
rect 3250 5468 3314 5472
rect 3250 5412 3254 5468
rect 3254 5412 3310 5468
rect 3310 5412 3314 5468
rect 3250 5408 3314 5412
rect 3330 5468 3394 5472
rect 3330 5412 3334 5468
rect 3334 5412 3390 5468
rect 3390 5412 3394 5468
rect 3330 5408 3394 5412
rect 3410 5468 3474 5472
rect 3410 5412 3414 5468
rect 3414 5412 3470 5468
rect 3470 5412 3474 5468
rect 3410 5408 3474 5412
rect 3490 5468 3554 5472
rect 3490 5412 3494 5468
rect 3494 5412 3550 5468
rect 3550 5412 3554 5468
rect 3490 5408 3554 5412
rect 7848 5468 7912 5472
rect 7848 5412 7852 5468
rect 7852 5412 7908 5468
rect 7908 5412 7912 5468
rect 7848 5408 7912 5412
rect 7928 5468 7992 5472
rect 7928 5412 7932 5468
rect 7932 5412 7988 5468
rect 7988 5412 7992 5468
rect 7928 5408 7992 5412
rect 8008 5468 8072 5472
rect 8008 5412 8012 5468
rect 8012 5412 8068 5468
rect 8068 5412 8072 5468
rect 8008 5408 8072 5412
rect 8088 5468 8152 5472
rect 8088 5412 8092 5468
rect 8092 5412 8148 5468
rect 8148 5412 8152 5468
rect 8088 5408 8152 5412
rect 12445 5468 12509 5472
rect 12445 5412 12449 5468
rect 12449 5412 12505 5468
rect 12505 5412 12509 5468
rect 12445 5408 12509 5412
rect 12525 5468 12589 5472
rect 12525 5412 12529 5468
rect 12529 5412 12585 5468
rect 12585 5412 12589 5468
rect 12525 5408 12589 5412
rect 12605 5468 12669 5472
rect 12605 5412 12609 5468
rect 12609 5412 12665 5468
rect 12665 5412 12669 5468
rect 12605 5408 12669 5412
rect 12685 5468 12749 5472
rect 12685 5412 12689 5468
rect 12689 5412 12745 5468
rect 12745 5412 12749 5468
rect 12685 5408 12749 5412
rect 4108 5340 4172 5404
rect 3740 5204 3804 5268
rect 12204 5204 12268 5268
rect 7236 5128 7300 5132
rect 7236 5072 7286 5128
rect 7286 5072 7300 5128
rect 7236 5068 7300 5072
rect 5549 4924 5613 4928
rect 5549 4868 5553 4924
rect 5553 4868 5609 4924
rect 5609 4868 5613 4924
rect 5549 4864 5613 4868
rect 5629 4924 5693 4928
rect 5629 4868 5633 4924
rect 5633 4868 5689 4924
rect 5689 4868 5693 4924
rect 5629 4864 5693 4868
rect 5709 4924 5773 4928
rect 5709 4868 5713 4924
rect 5713 4868 5769 4924
rect 5769 4868 5773 4924
rect 5709 4864 5773 4868
rect 5789 4924 5853 4928
rect 5789 4868 5793 4924
rect 5793 4868 5849 4924
rect 5849 4868 5853 4924
rect 5789 4864 5853 4868
rect 10146 4924 10210 4928
rect 10146 4868 10150 4924
rect 10150 4868 10206 4924
rect 10206 4868 10210 4924
rect 10146 4864 10210 4868
rect 10226 4924 10290 4928
rect 10226 4868 10230 4924
rect 10230 4868 10286 4924
rect 10286 4868 10290 4924
rect 10226 4864 10290 4868
rect 10306 4924 10370 4928
rect 10306 4868 10310 4924
rect 10310 4868 10366 4924
rect 10366 4868 10370 4924
rect 10306 4864 10370 4868
rect 10386 4924 10450 4928
rect 10386 4868 10390 4924
rect 10390 4868 10446 4924
rect 10446 4868 10450 4924
rect 10386 4864 10450 4868
rect 3924 4524 3988 4588
rect 4476 4524 4540 4588
rect 3250 4380 3314 4384
rect 3250 4324 3254 4380
rect 3254 4324 3310 4380
rect 3310 4324 3314 4380
rect 3250 4320 3314 4324
rect 3330 4380 3394 4384
rect 3330 4324 3334 4380
rect 3334 4324 3390 4380
rect 3390 4324 3394 4380
rect 3330 4320 3394 4324
rect 3410 4380 3474 4384
rect 3410 4324 3414 4380
rect 3414 4324 3470 4380
rect 3470 4324 3474 4380
rect 3410 4320 3474 4324
rect 3490 4380 3554 4384
rect 3490 4324 3494 4380
rect 3494 4324 3550 4380
rect 3550 4324 3554 4380
rect 3490 4320 3554 4324
rect 7848 4380 7912 4384
rect 7848 4324 7852 4380
rect 7852 4324 7908 4380
rect 7908 4324 7912 4380
rect 7848 4320 7912 4324
rect 7928 4380 7992 4384
rect 7928 4324 7932 4380
rect 7932 4324 7988 4380
rect 7988 4324 7992 4380
rect 7928 4320 7992 4324
rect 8008 4380 8072 4384
rect 8008 4324 8012 4380
rect 8012 4324 8068 4380
rect 8068 4324 8072 4380
rect 8008 4320 8072 4324
rect 8088 4380 8152 4384
rect 8088 4324 8092 4380
rect 8092 4324 8148 4380
rect 8148 4324 8152 4380
rect 8088 4320 8152 4324
rect 12445 4380 12509 4384
rect 12445 4324 12449 4380
rect 12449 4324 12505 4380
rect 12505 4324 12509 4380
rect 12445 4320 12509 4324
rect 12525 4380 12589 4384
rect 12525 4324 12529 4380
rect 12529 4324 12585 4380
rect 12585 4324 12589 4380
rect 12525 4320 12589 4324
rect 12605 4380 12669 4384
rect 12605 4324 12609 4380
rect 12609 4324 12665 4380
rect 12665 4324 12669 4380
rect 12605 4320 12669 4324
rect 12685 4380 12749 4384
rect 12685 4324 12689 4380
rect 12689 4324 12745 4380
rect 12745 4324 12749 4380
rect 12685 4320 12749 4324
rect 4292 4312 4356 4316
rect 4292 4256 4342 4312
rect 4342 4256 4356 4312
rect 4292 4252 4356 4256
rect 9812 3980 9876 4044
rect 3004 3844 3068 3908
rect 3924 3904 3988 3908
rect 3924 3848 3974 3904
rect 3974 3848 3988 3904
rect 3924 3844 3988 3848
rect 5549 3836 5613 3840
rect 5549 3780 5553 3836
rect 5553 3780 5609 3836
rect 5609 3780 5613 3836
rect 5549 3776 5613 3780
rect 5629 3836 5693 3840
rect 5629 3780 5633 3836
rect 5633 3780 5689 3836
rect 5689 3780 5693 3836
rect 5629 3776 5693 3780
rect 5709 3836 5773 3840
rect 5709 3780 5713 3836
rect 5713 3780 5769 3836
rect 5769 3780 5773 3836
rect 5709 3776 5773 3780
rect 5789 3836 5853 3840
rect 5789 3780 5793 3836
rect 5793 3780 5849 3836
rect 5849 3780 5853 3836
rect 5789 3776 5853 3780
rect 10146 3836 10210 3840
rect 10146 3780 10150 3836
rect 10150 3780 10206 3836
rect 10206 3780 10210 3836
rect 10146 3776 10210 3780
rect 10226 3836 10290 3840
rect 10226 3780 10230 3836
rect 10230 3780 10286 3836
rect 10286 3780 10290 3836
rect 10226 3776 10290 3780
rect 10306 3836 10370 3840
rect 10306 3780 10310 3836
rect 10310 3780 10366 3836
rect 10366 3780 10370 3836
rect 10306 3776 10370 3780
rect 10386 3836 10450 3840
rect 10386 3780 10390 3836
rect 10390 3780 10446 3836
rect 10446 3780 10450 3836
rect 10386 3776 10450 3780
rect 9628 3768 9692 3772
rect 9628 3712 9678 3768
rect 9678 3712 9692 3768
rect 9628 3708 9692 3712
rect 3250 3292 3314 3296
rect 3250 3236 3254 3292
rect 3254 3236 3310 3292
rect 3310 3236 3314 3292
rect 3250 3232 3314 3236
rect 3330 3292 3394 3296
rect 3330 3236 3334 3292
rect 3334 3236 3390 3292
rect 3390 3236 3394 3292
rect 3330 3232 3394 3236
rect 3410 3292 3474 3296
rect 3410 3236 3414 3292
rect 3414 3236 3470 3292
rect 3470 3236 3474 3292
rect 3410 3232 3474 3236
rect 3490 3292 3554 3296
rect 3490 3236 3494 3292
rect 3494 3236 3550 3292
rect 3550 3236 3554 3292
rect 3490 3232 3554 3236
rect 7848 3292 7912 3296
rect 7848 3236 7852 3292
rect 7852 3236 7908 3292
rect 7908 3236 7912 3292
rect 7848 3232 7912 3236
rect 7928 3292 7992 3296
rect 7928 3236 7932 3292
rect 7932 3236 7988 3292
rect 7988 3236 7992 3292
rect 7928 3232 7992 3236
rect 8008 3292 8072 3296
rect 8008 3236 8012 3292
rect 8012 3236 8068 3292
rect 8068 3236 8072 3292
rect 8008 3232 8072 3236
rect 8088 3292 8152 3296
rect 8088 3236 8092 3292
rect 8092 3236 8148 3292
rect 8148 3236 8152 3292
rect 8088 3232 8152 3236
rect 12445 3292 12509 3296
rect 12445 3236 12449 3292
rect 12449 3236 12505 3292
rect 12505 3236 12509 3292
rect 12445 3232 12509 3236
rect 12525 3292 12589 3296
rect 12525 3236 12529 3292
rect 12529 3236 12585 3292
rect 12585 3236 12589 3292
rect 12525 3232 12589 3236
rect 12605 3292 12669 3296
rect 12605 3236 12609 3292
rect 12609 3236 12665 3292
rect 12665 3236 12669 3292
rect 12605 3232 12669 3236
rect 12685 3292 12749 3296
rect 12685 3236 12689 3292
rect 12689 3236 12745 3292
rect 12745 3236 12749 3292
rect 12685 3232 12749 3236
rect 4476 3224 4540 3228
rect 4476 3168 4526 3224
rect 4526 3168 4540 3224
rect 4476 3164 4540 3168
rect 9628 2952 9692 2956
rect 9628 2896 9678 2952
rect 9678 2896 9692 2952
rect 9628 2892 9692 2896
rect 4108 2756 4172 2820
rect 11284 2816 11348 2820
rect 11284 2760 11334 2816
rect 11334 2760 11348 2816
rect 11284 2756 11348 2760
rect 5549 2748 5613 2752
rect 5549 2692 5553 2748
rect 5553 2692 5609 2748
rect 5609 2692 5613 2748
rect 5549 2688 5613 2692
rect 5629 2748 5693 2752
rect 5629 2692 5633 2748
rect 5633 2692 5689 2748
rect 5689 2692 5693 2748
rect 5629 2688 5693 2692
rect 5709 2748 5773 2752
rect 5709 2692 5713 2748
rect 5713 2692 5769 2748
rect 5769 2692 5773 2748
rect 5709 2688 5773 2692
rect 5789 2748 5853 2752
rect 5789 2692 5793 2748
rect 5793 2692 5849 2748
rect 5849 2692 5853 2748
rect 5789 2688 5853 2692
rect 10146 2748 10210 2752
rect 10146 2692 10150 2748
rect 10150 2692 10206 2748
rect 10206 2692 10210 2748
rect 10146 2688 10210 2692
rect 10226 2748 10290 2752
rect 10226 2692 10230 2748
rect 10230 2692 10286 2748
rect 10286 2692 10290 2748
rect 10226 2688 10290 2692
rect 10306 2748 10370 2752
rect 10306 2692 10310 2748
rect 10310 2692 10366 2748
rect 10366 2692 10370 2748
rect 10306 2688 10370 2692
rect 10386 2748 10450 2752
rect 10386 2692 10390 2748
rect 10390 2692 10446 2748
rect 10446 2692 10450 2748
rect 10386 2688 10450 2692
rect 3924 2348 3988 2412
rect 3250 2204 3314 2208
rect 3250 2148 3254 2204
rect 3254 2148 3310 2204
rect 3310 2148 3314 2204
rect 3250 2144 3314 2148
rect 3330 2204 3394 2208
rect 3330 2148 3334 2204
rect 3334 2148 3390 2204
rect 3390 2148 3394 2204
rect 3330 2144 3394 2148
rect 3410 2204 3474 2208
rect 3410 2148 3414 2204
rect 3414 2148 3470 2204
rect 3470 2148 3474 2204
rect 3410 2144 3474 2148
rect 3490 2204 3554 2208
rect 3490 2148 3494 2204
rect 3494 2148 3550 2204
rect 3550 2148 3554 2204
rect 3490 2144 3554 2148
rect 7848 2204 7912 2208
rect 7848 2148 7852 2204
rect 7852 2148 7908 2204
rect 7908 2148 7912 2204
rect 7848 2144 7912 2148
rect 7928 2204 7992 2208
rect 7928 2148 7932 2204
rect 7932 2148 7988 2204
rect 7988 2148 7992 2204
rect 7928 2144 7992 2148
rect 8008 2204 8072 2208
rect 8008 2148 8012 2204
rect 8012 2148 8068 2204
rect 8068 2148 8072 2204
rect 8008 2144 8072 2148
rect 8088 2204 8152 2208
rect 8088 2148 8092 2204
rect 8092 2148 8148 2204
rect 8148 2148 8152 2204
rect 8088 2144 8152 2148
rect 12445 2204 12509 2208
rect 12445 2148 12449 2204
rect 12449 2148 12505 2204
rect 12505 2148 12509 2204
rect 12445 2144 12509 2148
rect 12525 2204 12589 2208
rect 12525 2148 12529 2204
rect 12529 2148 12585 2204
rect 12585 2148 12589 2204
rect 12525 2144 12589 2148
rect 12605 2204 12669 2208
rect 12605 2148 12609 2204
rect 12609 2148 12665 2204
rect 12665 2148 12669 2204
rect 12605 2144 12669 2148
rect 12685 2204 12749 2208
rect 12685 2148 12689 2204
rect 12689 2148 12745 2204
rect 12745 2148 12749 2204
rect 12685 2144 12749 2148
<< metal4 >>
rect 3242 13088 3563 13648
rect 3242 13024 3250 13088
rect 3314 13024 3330 13088
rect 3394 13024 3410 13088
rect 3474 13024 3490 13088
rect 3554 13024 3563 13088
rect 2819 12476 2885 12477
rect 2819 12412 2820 12476
rect 2884 12412 2885 12476
rect 2819 12411 2885 12412
rect 2822 9349 2882 12411
rect 3242 12000 3563 13024
rect 3242 11936 3250 12000
rect 3314 11936 3330 12000
rect 3394 11936 3410 12000
rect 3474 11936 3490 12000
rect 3554 11936 3563 12000
rect 3242 10912 3563 11936
rect 5541 13632 5861 13648
rect 5541 13568 5549 13632
rect 5613 13568 5629 13632
rect 5693 13568 5709 13632
rect 5773 13568 5789 13632
rect 5853 13568 5861 13632
rect 5541 12544 5861 13568
rect 5541 12480 5549 12544
rect 5613 12480 5629 12544
rect 5693 12480 5709 12544
rect 5773 12480 5789 12544
rect 5853 12480 5861 12544
rect 5541 11456 5861 12480
rect 5541 11392 5549 11456
rect 5613 11392 5629 11456
rect 5693 11392 5709 11456
rect 5773 11392 5789 11456
rect 5853 11392 5861 11456
rect 3739 11252 3805 11253
rect 3739 11188 3740 11252
rect 3804 11188 3805 11252
rect 3739 11187 3805 11188
rect 3242 10848 3250 10912
rect 3314 10848 3330 10912
rect 3394 10848 3410 10912
rect 3474 10848 3490 10912
rect 3554 10848 3563 10912
rect 3003 10300 3069 10301
rect 3003 10236 3004 10300
rect 3068 10236 3069 10300
rect 3003 10235 3069 10236
rect 2819 9348 2885 9349
rect 2819 9284 2820 9348
rect 2884 9284 2885 9348
rect 2819 9283 2885 9284
rect 3006 3909 3066 10235
rect 3242 9824 3563 10848
rect 3242 9760 3250 9824
rect 3314 9760 3330 9824
rect 3394 9760 3410 9824
rect 3474 9760 3490 9824
rect 3554 9760 3563 9824
rect 3242 8736 3563 9760
rect 3242 8672 3250 8736
rect 3314 8672 3330 8736
rect 3394 8672 3410 8736
rect 3474 8672 3490 8736
rect 3554 8672 3563 8736
rect 3242 7648 3563 8672
rect 3242 7584 3250 7648
rect 3314 7584 3330 7648
rect 3394 7584 3410 7648
rect 3474 7584 3490 7648
rect 3554 7584 3563 7648
rect 3242 6560 3563 7584
rect 3242 6496 3250 6560
rect 3314 6496 3330 6560
rect 3394 6496 3410 6560
rect 3474 6496 3490 6560
rect 3554 6496 3563 6560
rect 3242 5472 3563 6496
rect 3242 5408 3250 5472
rect 3314 5408 3330 5472
rect 3394 5408 3410 5472
rect 3474 5408 3490 5472
rect 3554 5408 3563 5472
rect 3242 4384 3563 5408
rect 3742 5269 3802 11187
rect 4107 11116 4173 11117
rect 4107 11052 4108 11116
rect 4172 11052 4173 11116
rect 4107 11051 4173 11052
rect 3923 10980 3989 10981
rect 3923 10916 3924 10980
rect 3988 10916 3989 10980
rect 3923 10915 3989 10916
rect 3739 5268 3805 5269
rect 3739 5204 3740 5268
rect 3804 5204 3805 5268
rect 3739 5203 3805 5204
rect 3926 4589 3986 10915
rect 4110 5405 4170 11051
rect 5541 10368 5861 11392
rect 5541 10304 5549 10368
rect 5613 10304 5629 10368
rect 5693 10304 5709 10368
rect 5773 10304 5789 10368
rect 5853 10304 5861 10368
rect 4475 9620 4541 9621
rect 4475 9556 4476 9620
rect 4540 9556 4541 9620
rect 4475 9555 4541 9556
rect 4291 8940 4357 8941
rect 4291 8876 4292 8940
rect 4356 8876 4357 8940
rect 4291 8875 4357 8876
rect 4107 5404 4173 5405
rect 4107 5340 4108 5404
rect 4172 5340 4173 5404
rect 4107 5339 4173 5340
rect 3923 4588 3989 4589
rect 3923 4524 3924 4588
rect 3988 4524 3989 4588
rect 3923 4523 3989 4524
rect 3242 4320 3250 4384
rect 3314 4320 3330 4384
rect 3394 4320 3410 4384
rect 3474 4320 3490 4384
rect 3554 4320 3563 4384
rect 3003 3908 3069 3909
rect 3003 3844 3004 3908
rect 3068 3844 3069 3908
rect 3003 3843 3069 3844
rect 3242 3296 3563 4320
rect 3923 3908 3989 3909
rect 3923 3844 3924 3908
rect 3988 3844 3989 3908
rect 3923 3843 3989 3844
rect 3242 3232 3250 3296
rect 3314 3232 3330 3296
rect 3394 3232 3410 3296
rect 3474 3232 3490 3296
rect 3554 3232 3563 3296
rect 3242 2208 3563 3232
rect 3926 2413 3986 3843
rect 4110 2821 4170 5339
rect 4294 4317 4354 8875
rect 4478 4589 4538 9555
rect 5541 9280 5861 10304
rect 5541 9216 5549 9280
rect 5613 9216 5629 9280
rect 5693 9216 5709 9280
rect 5773 9216 5789 9280
rect 5853 9216 5861 9280
rect 5541 8192 5861 9216
rect 5541 8128 5549 8192
rect 5613 8128 5629 8192
rect 5693 8128 5709 8192
rect 5773 8128 5789 8192
rect 5853 8128 5861 8192
rect 5541 7104 5861 8128
rect 5541 7040 5549 7104
rect 5613 7040 5629 7104
rect 5693 7040 5709 7104
rect 5773 7040 5789 7104
rect 5853 7040 5861 7104
rect 5541 6016 5861 7040
rect 7840 13088 8160 13648
rect 7840 13024 7848 13088
rect 7912 13024 7928 13088
rect 7992 13024 8008 13088
rect 8072 13024 8088 13088
rect 8152 13024 8160 13088
rect 7840 12000 8160 13024
rect 10138 13632 10458 13648
rect 10138 13568 10146 13632
rect 10210 13568 10226 13632
rect 10290 13568 10306 13632
rect 10370 13568 10386 13632
rect 10450 13568 10458 13632
rect 9811 12884 9877 12885
rect 9811 12820 9812 12884
rect 9876 12820 9877 12884
rect 9811 12819 9877 12820
rect 7840 11936 7848 12000
rect 7912 11936 7928 12000
rect 7992 11936 8008 12000
rect 8072 11936 8088 12000
rect 8152 11936 8160 12000
rect 7840 10912 8160 11936
rect 7840 10848 7848 10912
rect 7912 10848 7928 10912
rect 7992 10848 8008 10912
rect 8072 10848 8088 10912
rect 8152 10848 8160 10912
rect 7840 9824 8160 10848
rect 7840 9760 7848 9824
rect 7912 9760 7928 9824
rect 7992 9760 8008 9824
rect 8072 9760 8088 9824
rect 8152 9760 8160 9824
rect 7840 8736 8160 9760
rect 7840 8672 7848 8736
rect 7912 8672 7928 8736
rect 7992 8672 8008 8736
rect 8072 8672 8088 8736
rect 8152 8672 8160 8736
rect 7840 7648 8160 8672
rect 7840 7584 7848 7648
rect 7912 7584 7928 7648
rect 7992 7584 8008 7648
rect 8072 7584 8088 7648
rect 8152 7584 8160 7648
rect 7235 6764 7301 6765
rect 7235 6700 7236 6764
rect 7300 6700 7301 6764
rect 7235 6699 7301 6700
rect 5541 5952 5549 6016
rect 5613 5952 5629 6016
rect 5693 5952 5709 6016
rect 5773 5952 5789 6016
rect 5853 5952 5861 6016
rect 5541 4928 5861 5952
rect 7238 5133 7298 6699
rect 7840 6560 8160 7584
rect 7840 6496 7848 6560
rect 7912 6496 7928 6560
rect 7992 6496 8008 6560
rect 8072 6496 8088 6560
rect 8152 6496 8160 6560
rect 7840 5472 8160 6496
rect 7840 5408 7848 5472
rect 7912 5408 7928 5472
rect 7992 5408 8008 5472
rect 8072 5408 8088 5472
rect 8152 5408 8160 5472
rect 7235 5132 7301 5133
rect 7235 5068 7236 5132
rect 7300 5068 7301 5132
rect 7235 5067 7301 5068
rect 5541 4864 5549 4928
rect 5613 4864 5629 4928
rect 5693 4864 5709 4928
rect 5773 4864 5789 4928
rect 5853 4864 5861 4928
rect 4475 4588 4541 4589
rect 4475 4524 4476 4588
rect 4540 4524 4541 4588
rect 4475 4523 4541 4524
rect 4291 4316 4357 4317
rect 4291 4252 4292 4316
rect 4356 4252 4357 4316
rect 4291 4251 4357 4252
rect 4478 3229 4538 4523
rect 5541 3840 5861 4864
rect 5541 3776 5549 3840
rect 5613 3776 5629 3840
rect 5693 3776 5709 3840
rect 5773 3776 5789 3840
rect 5853 3776 5861 3840
rect 4475 3228 4541 3229
rect 4475 3164 4476 3228
rect 4540 3164 4541 3228
rect 4475 3163 4541 3164
rect 4107 2820 4173 2821
rect 4107 2756 4108 2820
rect 4172 2756 4173 2820
rect 4107 2755 4173 2756
rect 5541 2752 5861 3776
rect 5541 2688 5549 2752
rect 5613 2688 5629 2752
rect 5693 2688 5709 2752
rect 5773 2688 5789 2752
rect 5853 2688 5861 2752
rect 3923 2412 3989 2413
rect 3923 2348 3924 2412
rect 3988 2348 3989 2412
rect 3923 2347 3989 2348
rect 3242 2144 3250 2208
rect 3314 2144 3330 2208
rect 3394 2144 3410 2208
rect 3474 2144 3490 2208
rect 3554 2144 3563 2208
rect 3242 2128 3563 2144
rect 5541 2128 5861 2688
rect 7840 4384 8160 5408
rect 7840 4320 7848 4384
rect 7912 4320 7928 4384
rect 7992 4320 8008 4384
rect 8072 4320 8088 4384
rect 8152 4320 8160 4384
rect 7840 3296 8160 4320
rect 9814 4045 9874 12819
rect 10138 12544 10458 13568
rect 10138 12480 10146 12544
rect 10210 12480 10226 12544
rect 10290 12480 10306 12544
rect 10370 12480 10386 12544
rect 10450 12480 10458 12544
rect 10138 11456 10458 12480
rect 10138 11392 10146 11456
rect 10210 11392 10226 11456
rect 10290 11392 10306 11456
rect 10370 11392 10386 11456
rect 10450 11392 10458 11456
rect 10138 10368 10458 11392
rect 10138 10304 10146 10368
rect 10210 10304 10226 10368
rect 10290 10304 10306 10368
rect 10370 10304 10386 10368
rect 10450 10304 10458 10368
rect 10138 9280 10458 10304
rect 12437 13088 12757 13648
rect 12437 13024 12445 13088
rect 12509 13024 12525 13088
rect 12589 13024 12605 13088
rect 12669 13024 12685 13088
rect 12749 13024 12757 13088
rect 12437 12000 12757 13024
rect 12437 11936 12445 12000
rect 12509 11936 12525 12000
rect 12589 11936 12605 12000
rect 12669 11936 12685 12000
rect 12749 11936 12757 12000
rect 12437 10912 12757 11936
rect 12437 10848 12445 10912
rect 12509 10848 12525 10912
rect 12589 10848 12605 10912
rect 12669 10848 12685 10912
rect 12749 10848 12757 10912
rect 12203 10028 12269 10029
rect 12203 9964 12204 10028
rect 12268 9964 12269 10028
rect 12203 9963 12269 9964
rect 10138 9216 10146 9280
rect 10210 9216 10226 9280
rect 10290 9216 10306 9280
rect 10370 9216 10386 9280
rect 10450 9216 10458 9280
rect 10138 8192 10458 9216
rect 11283 8668 11349 8669
rect 11283 8604 11284 8668
rect 11348 8604 11349 8668
rect 11283 8603 11349 8604
rect 10138 8128 10146 8192
rect 10210 8128 10226 8192
rect 10290 8128 10306 8192
rect 10370 8128 10386 8192
rect 10450 8128 10458 8192
rect 10138 7104 10458 8128
rect 10138 7040 10146 7104
rect 10210 7040 10226 7104
rect 10290 7040 10306 7104
rect 10370 7040 10386 7104
rect 10450 7040 10458 7104
rect 10138 6016 10458 7040
rect 10138 5952 10146 6016
rect 10210 5952 10226 6016
rect 10290 5952 10306 6016
rect 10370 5952 10386 6016
rect 10450 5952 10458 6016
rect 10138 4928 10458 5952
rect 10138 4864 10146 4928
rect 10210 4864 10226 4928
rect 10290 4864 10306 4928
rect 10370 4864 10386 4928
rect 10450 4864 10458 4928
rect 9811 4044 9877 4045
rect 9811 3980 9812 4044
rect 9876 3980 9877 4044
rect 9811 3979 9877 3980
rect 10138 3840 10458 4864
rect 10138 3776 10146 3840
rect 10210 3776 10226 3840
rect 10290 3776 10306 3840
rect 10370 3776 10386 3840
rect 10450 3776 10458 3840
rect 9627 3772 9693 3773
rect 9627 3708 9628 3772
rect 9692 3708 9693 3772
rect 9627 3707 9693 3708
rect 7840 3232 7848 3296
rect 7912 3232 7928 3296
rect 7992 3232 8008 3296
rect 8072 3232 8088 3296
rect 8152 3232 8160 3296
rect 7840 2208 8160 3232
rect 9630 2957 9690 3707
rect 9627 2956 9693 2957
rect 9627 2892 9628 2956
rect 9692 2892 9693 2956
rect 9627 2891 9693 2892
rect 7840 2144 7848 2208
rect 7912 2144 7928 2208
rect 7992 2144 8008 2208
rect 8072 2144 8088 2208
rect 8152 2144 8160 2208
rect 7840 2128 8160 2144
rect 10138 2752 10458 3776
rect 11286 2821 11346 8603
rect 11835 8124 11901 8125
rect 11835 8060 11836 8124
rect 11900 8060 11901 8124
rect 11835 8059 11901 8060
rect 11838 7173 11898 8059
rect 11835 7172 11901 7173
rect 11835 7108 11836 7172
rect 11900 7108 11901 7172
rect 11835 7107 11901 7108
rect 12206 5269 12266 9963
rect 12437 9824 12757 10848
rect 12437 9760 12445 9824
rect 12509 9760 12525 9824
rect 12589 9760 12605 9824
rect 12669 9760 12685 9824
rect 12749 9760 12757 9824
rect 12437 8736 12757 9760
rect 12437 8672 12445 8736
rect 12509 8672 12525 8736
rect 12589 8672 12605 8736
rect 12669 8672 12685 8736
rect 12749 8672 12757 8736
rect 12437 7648 12757 8672
rect 12437 7584 12445 7648
rect 12509 7584 12525 7648
rect 12589 7584 12605 7648
rect 12669 7584 12685 7648
rect 12749 7584 12757 7648
rect 12437 6560 12757 7584
rect 12437 6496 12445 6560
rect 12509 6496 12525 6560
rect 12589 6496 12605 6560
rect 12669 6496 12685 6560
rect 12749 6496 12757 6560
rect 12437 5472 12757 6496
rect 12437 5408 12445 5472
rect 12509 5408 12525 5472
rect 12589 5408 12605 5472
rect 12669 5408 12685 5472
rect 12749 5408 12757 5472
rect 12203 5268 12269 5269
rect 12203 5204 12204 5268
rect 12268 5204 12269 5268
rect 12203 5203 12269 5204
rect 12437 4384 12757 5408
rect 12437 4320 12445 4384
rect 12509 4320 12525 4384
rect 12589 4320 12605 4384
rect 12669 4320 12685 4384
rect 12749 4320 12757 4384
rect 12437 3296 12757 4320
rect 12437 3232 12445 3296
rect 12509 3232 12525 3296
rect 12589 3232 12605 3296
rect 12669 3232 12685 3296
rect 12749 3232 12757 3296
rect 11283 2820 11349 2821
rect 11283 2756 11284 2820
rect 11348 2756 11349 2820
rect 11283 2755 11349 2756
rect 10138 2688 10146 2752
rect 10210 2688 10226 2752
rect 10290 2688 10306 2752
rect 10370 2688 10386 2752
rect 10450 2688 10458 2752
rect 10138 2128 10458 2688
rect 12437 2208 12757 3232
rect 12437 2144 12445 2208
rect 12509 2144 12525 2208
rect 12589 2144 12605 2208
rect 12669 2144 12685 2208
rect 12749 2144 12757 2208
rect 12437 2128 12757 2144
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__3.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__4.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2852 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__5.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4600 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28
timestamp 1604681595
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _24_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5704 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5152 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_54 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6072 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__1.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_0_79 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8372 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_78
timestamp 1604681595
transform 1 0 8280 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_98
timestamp 1604681595
transform 1 0 10120 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_90
timestamp 1604681595
transform 1 0 9384 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1604681595
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604681595
transform 1 0 13340 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1604681595
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_131
timestamp 1604681595
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_137
timestamp 1604681595
transform 1 0 13708 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1604681595
transform 1 0 14444 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 4876 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1604681595
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 5612 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__2.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6716 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_53
timestamp 1604681595
transform 1 0 5980 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_77
timestamp 1604681595
transform 1 0 8188 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1604681595
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_99
timestamp 1604681595
transform 1 0 10212 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 12236 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp 1604681595
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_113
timestamp 1604681595
transform 1 0 11500 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_125
timestamp 1604681595
transform 1 0 12604 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604681595
transform 1 0 13340 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_137
timestamp 1604681595
transform 1 0 13708 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2208 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 4508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 3680 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 3036 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_41
timestamp 1604681595
transform 1 0 4876 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5428 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8372 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_95
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_107
timestamp 1604681595
transform 1 0 10948 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1604681595
transform 1 0 13340 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1604681595
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_137
timestamp 1604681595
transform 1 0 13708 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_145
timestamp 1604681595
transform 1 0 14444 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_12
timestamp 1604681595
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_48
timestamp 1604681595
transform 1 0 5520 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_60
timestamp 1604681595
transform 1 0 6624 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_77
timestamp 1604681595
transform 1 0 8188 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10304 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1604681595
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_99
timestamp 1604681595
transform 1 0 10212 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_109
timestamp 1604681595
transform 1 0 11132 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_128
timestamp 1604681595
transform 1 0 12880 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_140
timestamp 1604681595
transform 1 0 13984 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2208 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4876 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 3312 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_21
timestamp 1604681595
transform 1 0 3036 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_33
timestamp 1604681595
transform 1 0 4140 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_50
timestamp 1604681595
transform 1 0 5704 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 6900 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8004 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_67
timestamp 1604681595
transform 1 0 7268 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9936 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 9568 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_84
timestamp 1604681595
transform 1 0 8832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1604681595
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12512 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_105
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_117 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1604681595
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_133
timestamp 1604681595
transform 1 0 13340 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_145
timestamp 1604681595
transform 1 0 14444 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _06_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _13_
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2392 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_6
timestamp 1604681595
transform 1 0 1656 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4416 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_30
timestamp 1604681595
transform 1 0 3864 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5244 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 5336 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1604681595
transform 1 0 6808 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7268 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_74
timestamp 1604681595
transform 1 0 7912 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_66
timestamp 1604681595
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_83
timestamp 1604681595
transform 1 0 8740 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9476 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12604 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12604 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1604681595
transform 1 0 11132 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1604681595
transform 1 0 12236 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_107
timestamp 1604681595
transform 1 0 10948 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp 1604681595
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_134
timestamp 1604681595
transform 1 0 13432 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_134
timestamp 1604681595
transform 1 0 13432 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_6
timestamp 1604681595
transform 1 0 1656 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6624 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_47
timestamp 1604681595
transform 1 0 5428 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_59
timestamp 1604681595
transform 1 0 6532 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9936 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1604681595
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12144 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_8_112
timestamp 1604681595
transform 1 0 11408 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_136
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1604681595
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1604681595
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4508 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_29
timestamp 1604681595
transform 1 0 3772 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_46
timestamp 1604681595
transform 1 0 5336 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1604681595
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_70
timestamp 1604681595
transform 1 0 7544 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_80
timestamp 1604681595
transform 1 0 8464 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10304 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_92
timestamp 1604681595
transform 1 0 9568 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_109
timestamp 1604681595
transform 1 0 11132 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1604681595
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_144
timestamp 1604681595
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_48
timestamp 1604681595
transform 1 0 5520 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_60
timestamp 1604681595
transform 1 0 6624 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6900 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_72
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_101
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_125
timestamp 1604681595
transform 1 0 12604 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_137
timestamp 1604681595
transform 1 0 13708 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_20
timestamp 1604681595
transform 1 0 2944 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3772 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_28
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_38
timestamp 1604681595
transform 1 0 4600 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1604681595
transform 1 0 5612 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 5336 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_53
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_71
timestamp 1604681595
transform 1 0 7636 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 9936 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_88
timestamp 1604681595
transform 1 0 9200 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_99
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_132
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_144
timestamp 1604681595
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _07_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_6
timestamp 1604681595
transform 1 0 1656 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_58
timestamp 1604681595
transform 1 0 6440 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7176 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 8740 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 1604681595
transform 1 0 8004 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10120 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_86
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1604681595
transform 1 0 10028 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12328 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_114
timestamp 1604681595
transform 1 0 11592 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_131
timestamp 1604681595
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_143
timestamp 1604681595
transform 1 0 14260 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2208 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_11
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3864 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4692 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_21
timestamp 1604681595
transform 1 0 3036 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_29
timestamp 1604681595
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_38
timestamp 1604681595
transform 1 0 4600 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_46
timestamp 1604681595
transform 1 0 5336 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_58
timestamp 1604681595
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_55
timestamp 1604681595
transform 1 0 6164 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7176 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_13_66
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_63
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_82
timestamp 1604681595
transform 1 0 8648 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1604681595
transform 1 0 9936 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_90
timestamp 1604681595
transform 1 0 9384 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_100
timestamp 1604681595
transform 1 0 10304 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11040 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_124
timestamp 1604681595
transform 1 0 12512 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 13340 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_132
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_144
timestamp 1604681595
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_132
timestamp 1604681595
transform 1 0 13248 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_137
timestamp 1604681595
transform 1 0 13708 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_11
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_35
timestamp 1604681595
transform 1 0 4324 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 5060 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_47
timestamp 1604681595
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_72
timestamp 1604681595
transform 1 0 7728 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 10028 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_89
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_101
timestamp 1604681595
transform 1 0 10396 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_109
timestamp 1604681595
transform 1 0 11132 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_144
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_28
timestamp 1604681595
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1604681595
transform 1 0 5980 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_61
timestamp 1604681595
transform 1 0 6716 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _08_
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_67
timestamp 1604681595
transform 1 0 7268 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _10_
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_109
timestamp 1604681595
transform 1 0 11132 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_120
timestamp 1604681595
transform 1 0 12144 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1604681595
transform 1 0 13340 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_132
timestamp 1604681595
transform 1 0 13248 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_137
timestamp 1604681595
transform 1 0 13708 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_13
timestamp 1604681595
transform 1 0 2300 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3036 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _12_
timestamp 1604681595
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_42
timestamp 1604681595
transform 1 0 4968 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_71
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_88
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_100
timestamp 1604681595
transform 1 0 10304 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_104
timestamp 1604681595
transform 1 0 10672 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_144
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1604681595
transform 1 0 2116 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_48
timestamp 1604681595
transform 1 0 5520 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_60
timestamp 1604681595
transform 1 0 6624 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6900 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_72
timestamp 1604681595
transform 1 0 7728 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 11224 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 12328 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_109
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_114
timestamp 1604681595
transform 1 0 11592 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 13432 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_126
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_138
timestamp 1604681595
transform 1 0 13800 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1604681595
transform 1 0 2116 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1604681595
transform 1 0 2116 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1604681595
transform 1 0 3220 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 4324 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_36
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 5428 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_48
timestamp 1604681595
transform 1 0 5520 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1604681595
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 8556 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_66
timestamp 1604681595
transform 1 0 7176 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_78
timestamp 1604681595
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_83
timestamp 1604681595
transform 1 0 8740 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_63
timestamp 1604681595
transform 1 0 6900 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_73
timestamp 1604681595
transform 1 0 7820 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_95
timestamp 1604681595
transform 1 0 9844 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_102
timestamp 1604681595
transform 1 0 10488 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1604681595
transform 1 0 8924 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_103
timestamp 1604681595
transform 1 0 10580 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 11316 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_115
timestamp 1604681595
transform 1 0 11684 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_125
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _09_
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_127
timestamp 1604681595
transform 1 0 12788 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_138
timestamp 1604681595
transform 1 0 13800 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_137
timestamp 1604681595
transform 1 0 13708 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5262 0 5318 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 5170 15520 5226 16000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 5814 0 5870 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 5906 15520 5962 16000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 294 0 350 480 6 bottom_grid_pin_0_
port 4 nsew default tristate
rlabel metal2 s 3054 0 3110 480 6 bottom_grid_pin_10_
port 5 nsew default tristate
rlabel metal2 s 846 0 902 480 6 bottom_grid_pin_2_
port 6 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 bottom_grid_pin_4_
port 7 nsew default tristate
rlabel metal2 s 1950 0 2006 480 6 bottom_grid_pin_6_
port 8 nsew default tristate
rlabel metal2 s 2502 0 2558 480 6 bottom_grid_pin_8_
port 9 nsew default tristate
rlabel metal2 s 3606 0 3662 480 6 ccff_head
port 10 nsew default input
rlabel metal2 s 4158 0 4214 480 6 ccff_tail
port 11 nsew default tristate
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[0]
port 12 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_left_in[10]
port 13 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[11]
port 14 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[12]
port 15 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[13]
port 16 nsew default input
rlabel metal3 s 0 13744 480 13864 6 chanx_left_in[14]
port 17 nsew default input
rlabel metal3 s 0 14152 480 14272 6 chanx_left_in[15]
port 18 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[16]
port 19 nsew default input
rlabel metal3 s 0 14968 480 15088 6 chanx_left_in[17]
port 20 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[18]
port 21 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[19]
port 22 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[1]
port 23 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[2]
port 24 nsew default input
rlabel metal3 s 0 9256 480 9376 6 chanx_left_in[3]
port 25 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[4]
port 26 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[5]
port 27 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[6]
port 28 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[7]
port 29 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[8]
port 30 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[9]
port 31 nsew default input
rlabel metal3 s 0 144 480 264 6 chanx_left_out[0]
port 32 nsew default tristate
rlabel metal3 s 0 4088 480 4208 6 chanx_left_out[10]
port 33 nsew default tristate
rlabel metal3 s 0 4496 480 4616 6 chanx_left_out[11]
port 34 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 chanx_left_out[12]
port 35 nsew default tristate
rlabel metal3 s 0 5312 480 5432 6 chanx_left_out[13]
port 36 nsew default tristate
rlabel metal3 s 0 5720 480 5840 6 chanx_left_out[14]
port 37 nsew default tristate
rlabel metal3 s 0 6128 480 6248 6 chanx_left_out[15]
port 38 nsew default tristate
rlabel metal3 s 0 6536 480 6656 6 chanx_left_out[16]
port 39 nsew default tristate
rlabel metal3 s 0 6944 480 7064 6 chanx_left_out[17]
port 40 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[18]
port 41 nsew default tristate
rlabel metal3 s 0 7760 480 7880 6 chanx_left_out[19]
port 42 nsew default tristate
rlabel metal3 s 0 416 480 536 6 chanx_left_out[1]
port 43 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[2]
port 44 nsew default tristate
rlabel metal3 s 0 1232 480 1352 6 chanx_left_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 1640 480 1760 6 chanx_left_out[4]
port 46 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 chanx_left_out[6]
port 48 nsew default tristate
rlabel metal3 s 0 2864 480 2984 6 chanx_left_out[7]
port 49 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[8]
port 50 nsew default tristate
rlabel metal3 s 0 3680 480 3800 6 chanx_left_out[9]
port 51 nsew default tristate
rlabel metal3 s 15520 8168 16000 8288 6 chanx_right_in[0]
port 52 nsew default input
rlabel metal3 s 15520 12112 16000 12232 6 chanx_right_in[10]
port 53 nsew default input
rlabel metal3 s 15520 12520 16000 12640 6 chanx_right_in[11]
port 54 nsew default input
rlabel metal3 s 15520 12928 16000 13048 6 chanx_right_in[12]
port 55 nsew default input
rlabel metal3 s 15520 13336 16000 13456 6 chanx_right_in[13]
port 56 nsew default input
rlabel metal3 s 15520 13744 16000 13864 6 chanx_right_in[14]
port 57 nsew default input
rlabel metal3 s 15520 14152 16000 14272 6 chanx_right_in[15]
port 58 nsew default input
rlabel metal3 s 15520 14560 16000 14680 6 chanx_right_in[16]
port 59 nsew default input
rlabel metal3 s 15520 14968 16000 15088 6 chanx_right_in[17]
port 60 nsew default input
rlabel metal3 s 15520 15376 16000 15496 6 chanx_right_in[18]
port 61 nsew default input
rlabel metal3 s 15520 15784 16000 15904 6 chanx_right_in[19]
port 62 nsew default input
rlabel metal3 s 15520 8440 16000 8560 6 chanx_right_in[1]
port 63 nsew default input
rlabel metal3 s 15520 8848 16000 8968 6 chanx_right_in[2]
port 64 nsew default input
rlabel metal3 s 15520 9256 16000 9376 6 chanx_right_in[3]
port 65 nsew default input
rlabel metal3 s 15520 9664 16000 9784 6 chanx_right_in[4]
port 66 nsew default input
rlabel metal3 s 15520 10072 16000 10192 6 chanx_right_in[5]
port 67 nsew default input
rlabel metal3 s 15520 10480 16000 10600 6 chanx_right_in[6]
port 68 nsew default input
rlabel metal3 s 15520 10888 16000 11008 6 chanx_right_in[7]
port 69 nsew default input
rlabel metal3 s 15520 11296 16000 11416 6 chanx_right_in[8]
port 70 nsew default input
rlabel metal3 s 15520 11704 16000 11824 6 chanx_right_in[9]
port 71 nsew default input
rlabel metal3 s 15520 144 16000 264 6 chanx_right_out[0]
port 72 nsew default tristate
rlabel metal3 s 15520 4088 16000 4208 6 chanx_right_out[10]
port 73 nsew default tristate
rlabel metal3 s 15520 4496 16000 4616 6 chanx_right_out[11]
port 74 nsew default tristate
rlabel metal3 s 15520 4904 16000 5024 6 chanx_right_out[12]
port 75 nsew default tristate
rlabel metal3 s 15520 5312 16000 5432 6 chanx_right_out[13]
port 76 nsew default tristate
rlabel metal3 s 15520 5720 16000 5840 6 chanx_right_out[14]
port 77 nsew default tristate
rlabel metal3 s 15520 6128 16000 6248 6 chanx_right_out[15]
port 78 nsew default tristate
rlabel metal3 s 15520 6536 16000 6656 6 chanx_right_out[16]
port 79 nsew default tristate
rlabel metal3 s 15520 6944 16000 7064 6 chanx_right_out[17]
port 80 nsew default tristate
rlabel metal3 s 15520 7352 16000 7472 6 chanx_right_out[18]
port 81 nsew default tristate
rlabel metal3 s 15520 7760 16000 7880 6 chanx_right_out[19]
port 82 nsew default tristate
rlabel metal3 s 15520 416 16000 536 6 chanx_right_out[1]
port 83 nsew default tristate
rlabel metal3 s 15520 824 16000 944 6 chanx_right_out[2]
port 84 nsew default tristate
rlabel metal3 s 15520 1232 16000 1352 6 chanx_right_out[3]
port 85 nsew default tristate
rlabel metal3 s 15520 1640 16000 1760 6 chanx_right_out[4]
port 86 nsew default tristate
rlabel metal3 s 15520 2048 16000 2168 6 chanx_right_out[5]
port 87 nsew default tristate
rlabel metal3 s 15520 2456 16000 2576 6 chanx_right_out[6]
port 88 nsew default tristate
rlabel metal3 s 15520 2864 16000 2984 6 chanx_right_out[7]
port 89 nsew default tristate
rlabel metal3 s 15520 3272 16000 3392 6 chanx_right_out[8]
port 90 nsew default tristate
rlabel metal3 s 15520 3680 16000 3800 6 chanx_right_out[9]
port 91 nsew default tristate
rlabel metal2 s 6366 0 6422 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
port 92 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
port 93 nsew default tristate
rlabel metal2 s 7470 0 7526 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
port 94 nsew default tristate
rlabel metal2 s 8022 0 8078 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
port 95 nsew default tristate
rlabel metal2 s 8574 0 8630 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
port 96 nsew default tristate
rlabel metal2 s 9126 0 9182 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
port 97 nsew default tristate
rlabel metal2 s 9678 0 9734 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[0]
port 98 nsew default input
rlabel metal2 s 10230 0 10286 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[1]
port 99 nsew default input
rlabel metal2 s 10782 0 10838 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[2]
port 100 nsew default input
rlabel metal2 s 11334 0 11390 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[3]
port 101 nsew default input
rlabel metal2 s 11886 0 11942 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[4]
port 102 nsew default input
rlabel metal2 s 12438 0 12494 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[5]
port 103 nsew default input
rlabel metal2 s 12990 0 13046 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
port 104 nsew default tristate
rlabel metal2 s 13542 0 13598 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
port 105 nsew default tristate
rlabel metal2 s 14094 0 14150 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
port 106 nsew default tristate
rlabel metal2 s 14646 0 14702 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
port 107 nsew default tristate
rlabel metal2 s 15198 0 15254 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
port 108 nsew default tristate
rlabel metal2 s 15750 0 15806 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
port 109 nsew default tristate
rlabel metal2 s 4710 0 4766 480 6 prog_clk
port 110 nsew default input
rlabel metal2 s 6734 15520 6790 16000 6 top_width_0_height_0__pin_0_
port 111 nsew default input
rlabel metal2 s 10782 15520 10838 16000 6 top_width_0_height_0__pin_10_
port 112 nsew default input
rlabel metal2 s 15566 15520 15622 16000 6 top_width_0_height_0__pin_11_lower
port 113 nsew default tristate
rlabel metal2 s 4342 15520 4398 16000 6 top_width_0_height_0__pin_11_upper
port 114 nsew default tristate
rlabel metal2 s 11518 15520 11574 16000 6 top_width_0_height_0__pin_1_lower
port 115 nsew default tristate
rlabel metal2 s 386 15520 442 16000 6 top_width_0_height_0__pin_1_upper
port 116 nsew default tristate
rlabel metal2 s 7562 15520 7618 16000 6 top_width_0_height_0__pin_2_
port 117 nsew default input
rlabel metal2 s 12346 15520 12402 16000 6 top_width_0_height_0__pin_3_lower
port 118 nsew default tristate
rlabel metal2 s 1122 15520 1178 16000 6 top_width_0_height_0__pin_3_upper
port 119 nsew default tristate
rlabel metal2 s 8390 15520 8446 16000 6 top_width_0_height_0__pin_4_
port 120 nsew default input
rlabel metal2 s 13174 15520 13230 16000 6 top_width_0_height_0__pin_5_lower
port 121 nsew default tristate
rlabel metal2 s 1950 15520 2006 16000 6 top_width_0_height_0__pin_5_upper
port 122 nsew default tristate
rlabel metal2 s 9126 15520 9182 16000 6 top_width_0_height_0__pin_6_
port 123 nsew default input
rlabel metal2 s 13910 15520 13966 16000 6 top_width_0_height_0__pin_7_lower
port 124 nsew default tristate
rlabel metal2 s 2778 15520 2834 16000 6 top_width_0_height_0__pin_7_upper
port 125 nsew default tristate
rlabel metal2 s 9954 15520 10010 16000 6 top_width_0_height_0__pin_8_
port 126 nsew default input
rlabel metal2 s 14738 15520 14794 16000 6 top_width_0_height_0__pin_9_lower
port 127 nsew default tristate
rlabel metal2 s 3514 15520 3570 16000 6 top_width_0_height_0__pin_9_upper
port 128 nsew default tristate
rlabel metal4 s 3243 2128 3563 13648 6 VPWR
port 129 nsew default input
rlabel metal4 s 5541 2128 5861 13648 6 VGND
port 130 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 16000
<< end >>
