VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__1_
  CLASS BLOCK ;
  FOREIGN sb_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.000 BY 114.000 ;
  PIN Test_en_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 110.000 92.370 114.000 ;
    END
  END Test_en_N_out
  PIN Test_en_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END Test_en_S_in
  PIN bottom_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END bottom_left_grid_pin_42_
  PIN bottom_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END bottom_left_grid_pin_43_
  PIN bottom_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END bottom_left_grid_pin_44_
  PIN bottom_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END bottom_left_grid_pin_45_
  PIN bottom_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END bottom_left_grid_pin_46_
  PIN bottom_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END bottom_left_grid_pin_47_
  PIN bottom_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END bottom_left_grid_pin_48_
  PIN bottom_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END bottom_left_grid_pin_49_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 16.360 114.000 16.960 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 36.080 114.000 36.680 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 38.120 114.000 38.720 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 39.480 114.000 40.080 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 41.520 114.000 42.120 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 43.560 114.000 44.160 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 45.600 114.000 46.200 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 47.640 114.000 48.240 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 49.680 114.000 50.280 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 51.720 114.000 52.320 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 53.760 114.000 54.360 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 18.400 114.000 19.000 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 19.760 114.000 20.360 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 21.800 114.000 22.400 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 23.840 114.000 24.440 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 25.880 114.000 26.480 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 27.920 114.000 28.520 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 29.960 114.000 30.560 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 32.000 114.000 32.600 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 34.040 114.000 34.640 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 55.800 114.000 56.400 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 75.520 114.000 76.120 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 76.880 114.000 77.480 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 78.920 114.000 79.520 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 80.960 114.000 81.560 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 83.000 114.000 83.600 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 85.040 114.000 85.640 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 87.080 114.000 87.680 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 89.120 114.000 89.720 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 91.160 114.000 91.760 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 93.200 114.000 93.800 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 57.840 114.000 58.440 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 59.200 114.000 59.800 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 61.240 114.000 61.840 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 63.280 114.000 63.880 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 65.320 114.000 65.920 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 67.360 114.000 67.960 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 69.400 114.000 70.000 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 71.440 114.000 72.040 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 73.480 114.000 74.080 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.190 110.000 16.470 114.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 110.000 35.330 114.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 110.000 37.170 114.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 110.000 39.010 114.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 110.000 40.850 114.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 110.000 42.690 114.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.710 110.000 44.990 114.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 110.000 46.830 114.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 110.000 48.670 114.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 110.000 50.510 114.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 110.000 52.350 114.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 110.000 18.310 114.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 110.000 20.150 114.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 110.000 21.990 114.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 110.000 23.830 114.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 110.000 25.670 114.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.230 110.000 27.510 114.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 110.000 29.810 114.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 110.000 31.650 114.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 110.000 33.490 114.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.910 110.000 54.190 114.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.230 110.000 73.510 114.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.070 110.000 75.350 114.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 110.000 77.190 114.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.750 110.000 79.030 114.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.590 110.000 80.870 114.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.430 110.000 82.710 114.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.270 110.000 84.550 114.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 110.000 86.850 114.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 110.000 88.690 114.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 110.000 90.530 114.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.750 110.000 56.030 114.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.050 110.000 58.330 114.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 110.000 60.170 114.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.730 110.000 62.010 114.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.570 110.000 63.850 114.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 110.000 65.690 114.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.250 110.000 67.530 114.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 110.000 69.370 114.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.930 110.000 71.210 114.000 ;
    END
  END chany_top_out[9]
  PIN clk_1_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 102.720 114.000 103.320 ;
    END
  END clk_1_E_out
  PIN clk_1_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 110.000 94.210 114.000 ;
    END
  END clk_1_N_in
  PIN clk_1_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END clk_1_S_in
  PIN clk_1_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END clk_1_W_out
  PIN clk_2_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 95.240 114.000 95.840 ;
    END
  END clk_2_E_in
  PIN clk_2_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 104.760 114.000 105.360 ;
    END
  END clk_2_E_out
  PIN clk_2_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.770 110.000 96.050 114.000 ;
    END
  END clk_2_N_in
  PIN clk_2_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.270 110.000 107.550 114.000 ;
    END
  END clk_2_N_out
  PIN clk_2_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END clk_2_S_in
  PIN clk_2_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END clk_2_S_out
  PIN clk_2_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END clk_2_W_in
  PIN clk_2_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END clk_2_W_out
  PIN clk_3_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 96.600 114.000 97.200 ;
    END
  END clk_3_E_in
  PIN clk_3_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 106.800 114.000 107.400 ;
    END
  END clk_3_E_out
  PIN clk_3_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.610 110.000 97.890 114.000 ;
    END
  END clk_3_N_in
  PIN clk_3_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.110 110.000 109.390 114.000 ;
    END
  END clk_3_N_out
  PIN clk_3_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END clk_3_S_in
  PIN clk_3_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END clk_3_S_out
  PIN clk_3_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END clk_3_W_in
  PIN clk_3_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END clk_3_W_out
  PIN left_bottom_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END left_bottom_grid_pin_34_
  PIN left_bottom_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END left_bottom_grid_pin_35_
  PIN left_bottom_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END left_bottom_grid_pin_36_
  PIN left_bottom_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END left_bottom_grid_pin_37_
  PIN left_bottom_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END left_bottom_grid_pin_38_
  PIN left_bottom_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END left_bottom_grid_pin_39_
  PIN left_bottom_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END left_bottom_grid_pin_40_
  PIN left_bottom_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END left_bottom_grid_pin_41_
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.450 110.000 99.730 114.000 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_1_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 108.840 114.000 109.440 ;
    END
  END prog_clk_1_E_out
  PIN prog_clk_1_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.750 110.000 102.030 114.000 ;
    END
  END prog_clk_1_N_in
  PIN prog_clk_1_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END prog_clk_1_S_in
  PIN prog_clk_1_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END prog_clk_1_W_out
  PIN prog_clk_2_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 98.640 114.000 99.240 ;
    END
  END prog_clk_2_E_in
  PIN prog_clk_2_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 110.880 114.000 111.480 ;
    END
  END prog_clk_2_E_out
  PIN prog_clk_2_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.590 110.000 103.870 114.000 ;
    END
  END prog_clk_2_N_in
  PIN prog_clk_2_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 110.000 111.230 114.000 ;
    END
  END prog_clk_2_N_out
  PIN prog_clk_2_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END prog_clk_2_S_in
  PIN prog_clk_2_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END prog_clk_2_S_out
  PIN prog_clk_2_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END prog_clk_2_W_in
  PIN prog_clk_2_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END prog_clk_2_W_out
  PIN prog_clk_3_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 100.680 114.000 101.280 ;
    END
  END prog_clk_3_E_in
  PIN prog_clk_3_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 112.920 114.000 113.520 ;
    END
  END prog_clk_3_E_out
  PIN prog_clk_3_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 110.000 105.710 114.000 ;
    END
  END prog_clk_3_N_in
  PIN prog_clk_3_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.790 110.000 113.070 114.000 ;
    END
  END prog_clk_3_N_out
  PIN prog_clk_3_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END prog_clk_3_S_in
  PIN prog_clk_3_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END prog_clk_3_S_out
  PIN prog_clk_3_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END prog_clk_3_W_in
  PIN prog_clk_3_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END prog_clk_3_W_out
  PIN right_bottom_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 0.720 114.000 1.320 ;
    END
  END right_bottom_grid_pin_34_
  PIN right_bottom_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 2.080 114.000 2.680 ;
    END
  END right_bottom_grid_pin_35_
  PIN right_bottom_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 4.120 114.000 4.720 ;
    END
  END right_bottom_grid_pin_36_
  PIN right_bottom_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 6.160 114.000 6.760 ;
    END
  END right_bottom_grid_pin_37_
  PIN right_bottom_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 8.200 114.000 8.800 ;
    END
  END right_bottom_grid_pin_38_
  PIN right_bottom_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 10.240 114.000 10.840 ;
    END
  END right_bottom_grid_pin_39_
  PIN right_bottom_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 12.280 114.000 12.880 ;
    END
  END right_bottom_grid_pin_40_
  PIN right_bottom_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 14.320 114.000 14.920 ;
    END
  END right_bottom_grid_pin_41_
  PIN top_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 110.000 1.290 114.000 ;
    END
  END top_left_grid_pin_42_
  PIN top_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 110.000 3.130 114.000 ;
    END
  END top_left_grid_pin_43_
  PIN top_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 110.000 4.970 114.000 ;
    END
  END top_left_grid_pin_44_
  PIN top_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.530 110.000 6.810 114.000 ;
    END
  END top_left_grid_pin_45_
  PIN top_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.370 110.000 8.650 114.000 ;
    END
  END top_left_grid_pin_46_
  PIN top_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 110.000 10.490 114.000 ;
    END
  END top_left_grid_pin_47_
  PIN top_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 110.000 12.330 114.000 ;
    END
  END top_left_grid_pin_48_
  PIN top_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 110.000 14.170 114.000 ;
    END
  END top_left_grid_pin_49_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.880 10.640 23.480 100.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.040 10.640 40.640 100.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.100 100.725 ;
      LAYER met1 ;
        RECT 0.990 4.460 113.090 102.980 ;
      LAYER met2 ;
        RECT 1.570 109.720 2.570 113.405 ;
        RECT 3.410 109.720 4.410 113.405 ;
        RECT 5.250 109.720 6.250 113.405 ;
        RECT 7.090 109.720 8.090 113.405 ;
        RECT 8.930 109.720 9.930 113.405 ;
        RECT 10.770 109.720 11.770 113.405 ;
        RECT 12.610 109.720 13.610 113.405 ;
        RECT 14.450 109.720 15.910 113.405 ;
        RECT 16.750 109.720 17.750 113.405 ;
        RECT 18.590 109.720 19.590 113.405 ;
        RECT 20.430 109.720 21.430 113.405 ;
        RECT 22.270 109.720 23.270 113.405 ;
        RECT 24.110 109.720 25.110 113.405 ;
        RECT 25.950 109.720 26.950 113.405 ;
        RECT 27.790 109.720 29.250 113.405 ;
        RECT 30.090 109.720 31.090 113.405 ;
        RECT 31.930 109.720 32.930 113.405 ;
        RECT 33.770 109.720 34.770 113.405 ;
        RECT 35.610 109.720 36.610 113.405 ;
        RECT 37.450 109.720 38.450 113.405 ;
        RECT 39.290 109.720 40.290 113.405 ;
        RECT 41.130 109.720 42.130 113.405 ;
        RECT 42.970 109.720 44.430 113.405 ;
        RECT 45.270 109.720 46.270 113.405 ;
        RECT 47.110 109.720 48.110 113.405 ;
        RECT 48.950 109.720 49.950 113.405 ;
        RECT 50.790 109.720 51.790 113.405 ;
        RECT 52.630 109.720 53.630 113.405 ;
        RECT 54.470 109.720 55.470 113.405 ;
        RECT 56.310 109.720 57.770 113.405 ;
        RECT 58.610 109.720 59.610 113.405 ;
        RECT 60.450 109.720 61.450 113.405 ;
        RECT 62.290 109.720 63.290 113.405 ;
        RECT 64.130 109.720 65.130 113.405 ;
        RECT 65.970 109.720 66.970 113.405 ;
        RECT 67.810 109.720 68.810 113.405 ;
        RECT 69.650 109.720 70.650 113.405 ;
        RECT 71.490 109.720 72.950 113.405 ;
        RECT 73.790 109.720 74.790 113.405 ;
        RECT 75.630 109.720 76.630 113.405 ;
        RECT 77.470 109.720 78.470 113.405 ;
        RECT 79.310 109.720 80.310 113.405 ;
        RECT 81.150 109.720 82.150 113.405 ;
        RECT 82.990 109.720 83.990 113.405 ;
        RECT 84.830 109.720 86.290 113.405 ;
        RECT 87.130 109.720 88.130 113.405 ;
        RECT 88.970 109.720 89.970 113.405 ;
        RECT 90.810 109.720 91.810 113.405 ;
        RECT 92.650 109.720 93.650 113.405 ;
        RECT 94.490 109.720 95.490 113.405 ;
        RECT 96.330 109.720 97.330 113.405 ;
        RECT 98.170 109.720 99.170 113.405 ;
        RECT 100.010 109.720 101.470 113.405 ;
        RECT 102.310 109.720 103.310 113.405 ;
        RECT 104.150 109.720 105.150 113.405 ;
        RECT 105.990 109.720 106.990 113.405 ;
        RECT 107.830 109.720 108.830 113.405 ;
        RECT 109.670 109.720 110.670 113.405 ;
        RECT 111.510 109.720 112.510 113.405 ;
        RECT 1.020 4.280 113.060 109.720 ;
        RECT 1.570 0.835 2.570 4.280 ;
        RECT 3.410 0.835 4.410 4.280 ;
        RECT 5.250 0.835 6.250 4.280 ;
        RECT 7.090 0.835 8.090 4.280 ;
        RECT 8.930 0.835 9.930 4.280 ;
        RECT 10.770 0.835 11.770 4.280 ;
        RECT 12.610 0.835 13.610 4.280 ;
        RECT 14.450 0.835 15.450 4.280 ;
        RECT 16.290 0.835 17.290 4.280 ;
        RECT 18.130 0.835 19.130 4.280 ;
        RECT 19.970 0.835 20.970 4.280 ;
        RECT 21.810 0.835 22.810 4.280 ;
        RECT 23.650 0.835 24.650 4.280 ;
        RECT 25.490 0.835 26.490 4.280 ;
        RECT 27.330 0.835 28.330 4.280 ;
        RECT 29.170 0.835 30.630 4.280 ;
        RECT 31.470 0.835 32.470 4.280 ;
        RECT 33.310 0.835 34.310 4.280 ;
        RECT 35.150 0.835 36.150 4.280 ;
        RECT 36.990 0.835 37.990 4.280 ;
        RECT 38.830 0.835 39.830 4.280 ;
        RECT 40.670 0.835 41.670 4.280 ;
        RECT 42.510 0.835 43.510 4.280 ;
        RECT 44.350 0.835 45.350 4.280 ;
        RECT 46.190 0.835 47.190 4.280 ;
        RECT 48.030 0.835 49.030 4.280 ;
        RECT 49.870 0.835 50.870 4.280 ;
        RECT 51.710 0.835 52.710 4.280 ;
        RECT 53.550 0.835 54.550 4.280 ;
        RECT 55.390 0.835 56.390 4.280 ;
        RECT 57.230 0.835 58.690 4.280 ;
        RECT 59.530 0.835 60.530 4.280 ;
        RECT 61.370 0.835 62.370 4.280 ;
        RECT 63.210 0.835 64.210 4.280 ;
        RECT 65.050 0.835 66.050 4.280 ;
        RECT 66.890 0.835 67.890 4.280 ;
        RECT 68.730 0.835 69.730 4.280 ;
        RECT 70.570 0.835 71.570 4.280 ;
        RECT 72.410 0.835 73.410 4.280 ;
        RECT 74.250 0.835 75.250 4.280 ;
        RECT 76.090 0.835 77.090 4.280 ;
        RECT 77.930 0.835 78.930 4.280 ;
        RECT 79.770 0.835 80.770 4.280 ;
        RECT 81.610 0.835 82.610 4.280 ;
        RECT 83.450 0.835 84.450 4.280 ;
        RECT 85.290 0.835 86.750 4.280 ;
        RECT 87.590 0.835 88.590 4.280 ;
        RECT 89.430 0.835 90.430 4.280 ;
        RECT 91.270 0.835 92.270 4.280 ;
        RECT 93.110 0.835 94.110 4.280 ;
        RECT 94.950 0.835 95.950 4.280 ;
        RECT 96.790 0.835 97.790 4.280 ;
        RECT 98.630 0.835 99.630 4.280 ;
        RECT 100.470 0.835 101.470 4.280 ;
        RECT 102.310 0.835 103.310 4.280 ;
        RECT 104.150 0.835 105.150 4.280 ;
        RECT 105.990 0.835 106.990 4.280 ;
        RECT 107.830 0.835 108.830 4.280 ;
        RECT 109.670 0.835 110.670 4.280 ;
        RECT 111.510 0.835 112.510 4.280 ;
      LAYER met3 ;
        RECT 4.400 112.520 109.600 113.385 ;
        RECT 4.000 111.880 110.000 112.520 ;
        RECT 4.400 110.480 109.600 111.880 ;
        RECT 4.000 109.840 110.000 110.480 ;
        RECT 4.400 108.440 109.600 109.840 ;
        RECT 4.000 107.800 110.000 108.440 ;
        RECT 4.400 106.400 109.600 107.800 ;
        RECT 4.000 105.760 110.000 106.400 ;
        RECT 4.400 104.360 109.600 105.760 ;
        RECT 4.000 103.720 110.000 104.360 ;
        RECT 4.400 102.320 109.600 103.720 ;
        RECT 4.000 101.680 110.000 102.320 ;
        RECT 4.400 100.280 109.600 101.680 ;
        RECT 4.000 99.640 110.000 100.280 ;
        RECT 4.400 98.240 109.600 99.640 ;
        RECT 4.000 97.600 110.000 98.240 ;
        RECT 4.400 94.840 109.600 97.600 ;
        RECT 4.000 94.200 110.000 94.840 ;
        RECT 4.400 92.800 109.600 94.200 ;
        RECT 4.000 92.160 110.000 92.800 ;
        RECT 4.400 90.760 109.600 92.160 ;
        RECT 4.000 90.120 110.000 90.760 ;
        RECT 4.400 88.720 109.600 90.120 ;
        RECT 4.000 88.080 110.000 88.720 ;
        RECT 4.400 86.680 109.600 88.080 ;
        RECT 4.000 86.040 110.000 86.680 ;
        RECT 4.400 84.640 109.600 86.040 ;
        RECT 4.000 84.000 110.000 84.640 ;
        RECT 4.400 82.600 109.600 84.000 ;
        RECT 4.000 81.960 110.000 82.600 ;
        RECT 4.400 80.560 109.600 81.960 ;
        RECT 4.000 79.920 110.000 80.560 ;
        RECT 4.400 78.520 109.600 79.920 ;
        RECT 4.000 77.880 110.000 78.520 ;
        RECT 4.400 75.120 109.600 77.880 ;
        RECT 4.000 74.480 110.000 75.120 ;
        RECT 4.400 73.080 109.600 74.480 ;
        RECT 4.000 72.440 110.000 73.080 ;
        RECT 4.400 71.040 109.600 72.440 ;
        RECT 4.000 70.400 110.000 71.040 ;
        RECT 4.400 69.000 109.600 70.400 ;
        RECT 4.000 68.360 110.000 69.000 ;
        RECT 4.400 66.960 109.600 68.360 ;
        RECT 4.000 66.320 110.000 66.960 ;
        RECT 4.400 64.920 109.600 66.320 ;
        RECT 4.000 64.280 110.000 64.920 ;
        RECT 4.400 62.880 109.600 64.280 ;
        RECT 4.000 62.240 110.000 62.880 ;
        RECT 4.400 60.840 109.600 62.240 ;
        RECT 4.000 60.200 110.000 60.840 ;
        RECT 4.400 57.440 109.600 60.200 ;
        RECT 4.000 56.800 110.000 57.440 ;
        RECT 4.400 55.400 109.600 56.800 ;
        RECT 4.000 54.760 110.000 55.400 ;
        RECT 4.400 53.360 109.600 54.760 ;
        RECT 4.000 52.720 110.000 53.360 ;
        RECT 4.400 51.320 109.600 52.720 ;
        RECT 4.000 50.680 110.000 51.320 ;
        RECT 4.400 49.280 109.600 50.680 ;
        RECT 4.000 48.640 110.000 49.280 ;
        RECT 4.400 47.240 109.600 48.640 ;
        RECT 4.000 46.600 110.000 47.240 ;
        RECT 4.400 45.200 109.600 46.600 ;
        RECT 4.000 44.560 110.000 45.200 ;
        RECT 4.400 43.160 109.600 44.560 ;
        RECT 4.000 42.520 110.000 43.160 ;
        RECT 4.400 41.120 109.600 42.520 ;
        RECT 4.000 40.480 110.000 41.120 ;
        RECT 4.400 37.720 109.600 40.480 ;
        RECT 4.000 37.080 110.000 37.720 ;
        RECT 4.400 35.680 109.600 37.080 ;
        RECT 4.000 35.040 110.000 35.680 ;
        RECT 4.400 33.640 109.600 35.040 ;
        RECT 4.000 33.000 110.000 33.640 ;
        RECT 4.400 31.600 109.600 33.000 ;
        RECT 4.000 30.960 110.000 31.600 ;
        RECT 4.400 29.560 109.600 30.960 ;
        RECT 4.000 28.920 110.000 29.560 ;
        RECT 4.400 27.520 109.600 28.920 ;
        RECT 4.000 26.880 110.000 27.520 ;
        RECT 4.400 25.480 109.600 26.880 ;
        RECT 4.000 24.840 110.000 25.480 ;
        RECT 4.400 23.440 109.600 24.840 ;
        RECT 4.000 22.800 110.000 23.440 ;
        RECT 4.400 21.400 109.600 22.800 ;
        RECT 4.000 20.760 110.000 21.400 ;
        RECT 4.400 18.000 109.600 20.760 ;
        RECT 4.000 17.360 110.000 18.000 ;
        RECT 4.400 15.960 109.600 17.360 ;
        RECT 4.000 15.320 110.000 15.960 ;
        RECT 4.400 13.920 109.600 15.320 ;
        RECT 4.000 13.280 110.000 13.920 ;
        RECT 4.400 11.880 109.600 13.280 ;
        RECT 4.000 11.240 110.000 11.880 ;
        RECT 4.400 9.840 109.600 11.240 ;
        RECT 4.000 9.200 110.000 9.840 ;
        RECT 4.400 7.800 109.600 9.200 ;
        RECT 4.000 7.160 110.000 7.800 ;
        RECT 4.400 5.760 109.600 7.160 ;
        RECT 4.000 5.120 110.000 5.760 ;
        RECT 4.400 3.720 109.600 5.120 ;
        RECT 4.000 3.080 110.000 3.720 ;
        RECT 4.400 0.855 109.600 3.080 ;
      LAYER met4 ;
        RECT 24.215 10.240 38.640 100.880 ;
        RECT 41.040 10.240 100.905 100.880 ;
        RECT 24.215 9.695 100.905 10.240 ;
  END
END sb_1__1_
END LIBRARY

