magic
tech EFS8A
magscale 1 2
timestamp 1602269183
<< locali >>
rect 2823 24225 2858 24259
rect 8493 23137 8654 23171
rect 11563 23137 11598 23171
rect 8493 22967 8527 23137
rect 1639 18921 1777 18955
rect 10103 18377 10241 18411
rect 6319 16609 6354 16643
rect 7107 14569 7113 14603
rect 10051 14569 10057 14603
rect 7107 14501 7141 14569
rect 10051 14501 10085 14569
rect 2139 13719 2173 13787
rect 2139 13685 2145 13719
rect 4623 13481 4629 13515
rect 11707 13481 11713 13515
rect 4623 13413 4657 13481
rect 11707 13413 11741 13481
rect 6469 12767 6503 12869
rect 13179 12393 13185 12427
rect 13179 12325 13213 12393
rect 12863 11577 13001 11611
rect 1955 10455 1989 10523
rect 1955 10421 1961 10455
rect 3243 9367 3277 9435
rect 3243 9333 3249 9367
rect 16543 8585 16681 8619
rect 4353 8279 4387 8449
rect 2139 8041 2145 8075
rect 12351 8041 12357 8075
rect 2139 7973 2173 8041
rect 12351 7973 12385 8041
rect 15485 6239 15519 6409
rect 14335 5797 14473 5831
rect 8401 5015 8435 5185
rect 13461 5015 13495 5117
rect 13921 5015 13955 5321
rect 1443 4641 1478 4675
rect 6411 4233 6503 4267
rect 5549 3995 5583 4097
rect 6653 3927 6687 4233
rect 9413 3995 9447 4165
rect 11287 4029 11322 4063
rect 13363 3689 13369 3723
rect 13363 3621 13397 3689
rect 8619 3553 8654 3587
rect 14841 2975 14875 3145
rect 4399 2601 4537 2635
rect 6009 2397 6135 2431
rect 6101 2295 6135 2397
<< viali >>
rect 15485 24361 15519 24395
rect 2789 24225 2823 24259
rect 11964 24225 11998 24259
rect 12976 24225 13010 24259
rect 15301 24225 15335 24259
rect 24660 24225 24694 24259
rect 12541 24089 12575 24123
rect 2927 24021 2961 24055
rect 12035 24021 12069 24055
rect 13047 24021 13081 24055
rect 24731 24021 24765 24055
rect 2881 23817 2915 23851
rect 3157 23817 3191 23851
rect 4813 23817 4847 23851
rect 7021 23817 7055 23851
rect 9781 23817 9815 23851
rect 11989 23817 12023 23851
rect 13461 23817 13495 23851
rect 15853 23817 15887 23851
rect 17049 23817 17083 23851
rect 19533 23817 19567 23851
rect 21465 23817 21499 23851
rect 24593 23817 24627 23851
rect 25237 23817 25271 23851
rect 4399 23749 4433 23783
rect 19119 23749 19153 23783
rect 24225 23749 24259 23783
rect 9045 23681 9079 23715
rect 11621 23681 11655 23715
rect 12541 23681 12575 23715
rect 12817 23681 12851 23715
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 2973 23613 3007 23647
rect 4328 23613 4362 23647
rect 6837 23613 6871 23647
rect 7389 23613 7423 23647
rect 8652 23613 8686 23647
rect 9597 23613 9631 23647
rect 10149 23613 10183 23647
rect 16865 23613 16899 23647
rect 17417 23613 17451 23647
rect 19048 23613 19082 23647
rect 20980 23613 21014 23647
rect 23740 23613 23774 23647
rect 24752 23613 24786 23647
rect 12633 23545 12667 23579
rect 14933 23545 14967 23579
rect 15025 23545 15059 23579
rect 15577 23545 15611 23579
rect 1547 23477 1581 23511
rect 3617 23477 3651 23511
rect 8723 23477 8757 23511
rect 14749 23477 14783 23511
rect 21051 23477 21085 23511
rect 23811 23477 23845 23511
rect 24823 23477 24857 23511
rect 11667 23273 11701 23307
rect 14933 23273 14967 23307
rect 8723 23205 8757 23239
rect 12725 23205 12759 23239
rect 15485 23205 15519 23239
rect 11529 23137 11563 23171
rect 12633 23069 12667 23103
rect 13277 23069 13311 23103
rect 15393 23069 15427 23103
rect 15669 23069 15703 23103
rect 8493 22933 8527 22967
rect 1593 22729 1627 22763
rect 13461 22729 13495 22763
rect 14749 22729 14783 22763
rect 15945 22729 15979 22763
rect 12541 22593 12575 22627
rect 13829 22593 13863 22627
rect 1409 22525 1443 22559
rect 10701 22525 10735 22559
rect 11437 22525 11471 22559
rect 11897 22525 11931 22559
rect 14565 22525 14599 22559
rect 15485 22525 15519 22559
rect 11529 22457 11563 22491
rect 12173 22457 12207 22491
rect 12633 22457 12667 22491
rect 13185 22457 13219 22491
rect 2053 22389 2087 22423
rect 8585 22389 8619 22423
rect 14289 22389 14323 22423
rect 12541 22117 12575 22151
rect 12449 21981 12483 22015
rect 12725 21981 12759 22015
rect 11621 21845 11655 21879
rect 11897 21641 11931 21675
rect 12265 21505 12299 21539
rect 12449 21505 12483 21539
rect 12541 21437 12575 21471
rect 12449 20757 12483 20791
rect 1593 20553 1627 20587
rect 1409 20349 1443 20383
rect 1961 20349 1995 20383
rect 25145 19465 25179 19499
rect 1444 19261 1478 19295
rect 1869 19261 1903 19295
rect 24660 19261 24694 19295
rect 1547 19125 1581 19159
rect 24731 19125 24765 19159
rect 1777 18921 1811 18955
rect 2651 18921 2685 18955
rect 1568 18785 1602 18819
rect 2580 18785 2614 18819
rect 2053 18581 2087 18615
rect 10241 18377 10275 18411
rect 2145 18173 2179 18207
rect 2421 18173 2455 18207
rect 10032 18173 10066 18207
rect 10425 18173 10459 18207
rect 1777 18105 1811 18139
rect 1961 18037 1995 18071
rect 2973 18037 3007 18071
rect 4215 17833 4249 17867
rect 7757 17833 7791 17867
rect 9873 17765 9907 17799
rect 2145 17697 2179 17731
rect 2421 17697 2455 17731
rect 4144 17697 4178 17731
rect 7573 17697 7607 17731
rect 2329 17629 2363 17663
rect 9781 17629 9815 17663
rect 10149 17629 10183 17663
rect 1685 17493 1719 17527
rect 4629 17289 4663 17323
rect 9137 17289 9171 17323
rect 8309 17221 8343 17255
rect 8769 17153 8803 17187
rect 10149 17153 10183 17187
rect 11161 17153 11195 17187
rect 1961 17085 1995 17119
rect 2513 17085 2547 17119
rect 2789 17085 2823 17119
rect 3868 17085 3902 17119
rect 4261 17085 4295 17119
rect 7205 17085 7239 17119
rect 7665 17085 7699 17119
rect 9689 17017 9723 17051
rect 9781 17017 9815 17051
rect 2329 16949 2363 16983
rect 3249 16949 3283 16983
rect 3709 16949 3743 16983
rect 3939 16949 3973 16983
rect 7573 16949 7607 16983
rect 9505 16949 9539 16983
rect 10701 16949 10735 16983
rect 4721 16745 4755 16779
rect 6423 16745 6457 16779
rect 7481 16677 7515 16711
rect 9873 16677 9907 16711
rect 10425 16677 10459 16711
rect 11253 16677 11287 16711
rect 1869 16609 1903 16643
rect 4077 16609 4111 16643
rect 6285 16609 6319 16643
rect 11345 16609 11379 16643
rect 1777 16541 1811 16575
rect 4445 16541 4479 16575
rect 7389 16541 7423 16575
rect 9781 16541 9815 16575
rect 7941 16473 7975 16507
rect 2881 16405 2915 16439
rect 4215 16405 4249 16439
rect 4353 16405 4387 16439
rect 5089 16405 5123 16439
rect 1685 16201 1719 16235
rect 3157 16201 3191 16235
rect 5825 16201 5859 16235
rect 6653 16201 6687 16235
rect 7297 16201 7331 16235
rect 11621 16201 11655 16235
rect 3479 16133 3513 16167
rect 10977 16133 11011 16167
rect 1869 16065 1903 16099
rect 6285 16065 6319 16099
rect 7941 16065 7975 16099
rect 9137 16065 9171 16099
rect 10333 16065 10367 16099
rect 3376 15997 3410 16031
rect 5089 15997 5123 16031
rect 1961 15929 1995 15963
rect 2513 15929 2547 15963
rect 4445 15929 4479 15963
rect 7481 15929 7515 15963
rect 7573 15929 7607 15963
rect 8401 15929 8435 15963
rect 9689 15929 9723 15963
rect 9781 15929 9815 15963
rect 2881 15861 2915 15895
rect 4169 15861 4203 15895
rect 5457 15861 5491 15895
rect 9505 15861 9539 15895
rect 10701 15861 10735 15895
rect 11161 15861 11195 15895
rect 1685 15657 1719 15691
rect 8217 15657 8251 15691
rect 1961 15589 1995 15623
rect 6837 15589 6871 15623
rect 7389 15589 7423 15623
rect 8033 15589 8067 15623
rect 9689 15589 9723 15623
rect 4997 15521 5031 15555
rect 9781 15521 9815 15555
rect 11621 15521 11655 15555
rect 1869 15453 1903 15487
rect 6745 15453 6779 15487
rect 11253 15453 11287 15487
rect 2421 15385 2455 15419
rect 2881 15317 2915 15351
rect 3893 15317 3927 15351
rect 4629 15317 4663 15351
rect 7757 15317 7791 15351
rect 3157 15113 3191 15147
rect 3617 15113 3651 15147
rect 4077 15113 4111 15147
rect 5181 15113 5215 15147
rect 6193 15113 6227 15147
rect 11621 15113 11655 15147
rect 25145 15113 25179 15147
rect 2697 15045 2731 15079
rect 7113 15045 7147 15079
rect 11253 15045 11287 15079
rect 2145 14977 2179 15011
rect 4261 14977 4295 15011
rect 4721 14977 4755 15011
rect 5733 14977 5767 15011
rect 7757 14977 7791 15011
rect 8953 14977 8987 15011
rect 10149 14977 10183 15011
rect 10701 14977 10735 15011
rect 8861 14909 8895 14943
rect 9045 14909 9079 14943
rect 12449 14909 12483 14943
rect 12909 14909 12943 14943
rect 24660 14909 24694 14943
rect 2237 14841 2271 14875
rect 4353 14841 4387 14875
rect 7481 14841 7515 14875
rect 7573 14841 7607 14875
rect 10793 14841 10827 14875
rect 1869 14773 1903 14807
rect 6653 14773 6687 14807
rect 10517 14773 10551 14807
rect 12173 14773 12207 14807
rect 12541 14773 12575 14807
rect 24731 14773 24765 14807
rect 2237 14569 2271 14603
rect 7113 14569 7147 14603
rect 7665 14569 7699 14603
rect 9505 14569 9539 14603
rect 10057 14569 10091 14603
rect 10609 14569 10643 14603
rect 13093 14569 13127 14603
rect 2605 14501 2639 14535
rect 4537 14501 4571 14535
rect 11621 14501 11655 14535
rect 24225 14501 24259 14535
rect 1476 14433 1510 14467
rect 13001 14433 13035 14467
rect 13461 14433 13495 14467
rect 2513 14365 2547 14399
rect 2973 14365 3007 14399
rect 4445 14365 4479 14399
rect 4721 14365 4755 14399
rect 6745 14365 6779 14399
rect 9689 14365 9723 14399
rect 11345 14365 11379 14399
rect 11529 14365 11563 14399
rect 11805 14365 11839 14399
rect 24133 14365 24167 14399
rect 24777 14365 24811 14399
rect 1547 14229 1581 14263
rect 1961 14229 1995 14263
rect 5457 14229 5491 14263
rect 8953 14229 8987 14263
rect 12449 14229 12483 14263
rect 1593 14025 1627 14059
rect 2697 14025 2731 14059
rect 4077 14025 4111 14059
rect 4445 14025 4479 14059
rect 7757 14025 7791 14059
rect 8033 14025 8067 14059
rect 9781 14025 9815 14059
rect 11529 14025 11563 14059
rect 11805 14025 11839 14059
rect 12265 14025 12299 14059
rect 12817 14025 12851 14059
rect 14197 14025 14231 14059
rect 25145 14025 25179 14059
rect 1777 13889 1811 13923
rect 3341 13889 3375 13923
rect 3525 13889 3559 13923
rect 4629 13889 4663 13923
rect 4905 13889 4939 13923
rect 6837 13889 6871 13923
rect 8861 13889 8895 13923
rect 10609 13889 10643 13923
rect 14473 13889 14507 13923
rect 24225 13889 24259 13923
rect 13277 13821 13311 13855
rect 4721 13753 4755 13787
rect 5549 13753 5583 13787
rect 7158 13753 7192 13787
rect 9182 13753 9216 13787
rect 10930 13753 10964 13787
rect 13598 13753 13632 13787
rect 24317 13753 24351 13787
rect 24869 13753 24903 13787
rect 2145 13685 2179 13719
rect 2973 13685 3007 13719
rect 6285 13685 6319 13719
rect 6653 13685 6687 13719
rect 8677 13685 8711 13719
rect 10057 13685 10091 13719
rect 10425 13685 10459 13719
rect 13185 13685 13219 13719
rect 23489 13685 23523 13719
rect 24041 13685 24075 13719
rect 4629 13481 4663 13515
rect 5181 13481 5215 13515
rect 7849 13481 7883 13515
rect 9781 13481 9815 13515
rect 10793 13481 10827 13515
rect 11713 13481 11747 13515
rect 12265 13481 12299 13515
rect 13369 13481 13403 13515
rect 24041 13481 24075 13515
rect 2190 13413 2224 13447
rect 6193 13413 6227 13447
rect 7757 13345 7791 13379
rect 8033 13345 8067 13379
rect 9689 13345 9723 13379
rect 10149 13345 10183 13379
rect 13093 13345 13127 13379
rect 13553 13345 13587 13379
rect 23857 13345 23891 13379
rect 1869 13277 1903 13311
rect 3893 13277 3927 13311
rect 4261 13277 4295 13311
rect 5917 13277 5951 13311
rect 6101 13277 6135 13311
rect 6377 13277 6411 13311
rect 7481 13277 7515 13311
rect 8677 13277 8711 13311
rect 11345 13277 11379 13311
rect 2789 13141 2823 13175
rect 3157 13141 3191 13175
rect 7113 13141 7147 13175
rect 9413 13141 9447 13175
rect 11161 13141 11195 13175
rect 14289 13141 14323 13175
rect 24869 13141 24903 13175
rect 5365 12937 5399 12971
rect 7849 12937 7883 12971
rect 8217 12937 8251 12971
rect 6469 12869 6503 12903
rect 6561 12869 6595 12903
rect 13369 12869 13403 12903
rect 1869 12801 1903 12835
rect 3571 12801 3605 12835
rect 6285 12801 6319 12835
rect 9137 12801 9171 12835
rect 11161 12801 11195 12835
rect 12449 12801 12483 12835
rect 14289 12801 14323 12835
rect 14565 12801 14599 12835
rect 23857 12801 23891 12835
rect 2513 12733 2547 12767
rect 2881 12733 2915 12767
rect 3468 12733 3502 12767
rect 3893 12733 3927 12767
rect 4445 12733 4479 12767
rect 6469 12733 6503 12767
rect 6837 12733 6871 12767
rect 7389 12733 7423 12767
rect 8401 12733 8435 12767
rect 8953 12733 8987 12767
rect 10517 12733 10551 12767
rect 10977 12733 11011 12767
rect 13645 12733 13679 12767
rect 4353 12665 4387 12699
rect 4807 12665 4841 12699
rect 9689 12665 9723 12699
rect 10333 12665 10367 12699
rect 12770 12665 12804 12699
rect 14013 12665 14047 12699
rect 14381 12665 14415 12699
rect 1777 12597 1811 12631
rect 5733 12597 5767 12631
rect 7113 12597 7147 12631
rect 11529 12597 11563 12631
rect 12173 12597 12207 12631
rect 2605 12393 2639 12427
rect 4353 12393 4387 12427
rect 6009 12393 6043 12427
rect 10793 12393 10827 12427
rect 12541 12393 12575 12427
rect 13185 12393 13219 12427
rect 14381 12393 14415 12427
rect 6929 12325 6963 12359
rect 8769 12325 8803 12359
rect 9413 12325 9447 12359
rect 1685 12257 1719 12291
rect 4077 12257 4111 12291
rect 4905 12257 4939 12291
rect 5089 12257 5123 12291
rect 6193 12257 6227 12291
rect 7481 12257 7515 12291
rect 8033 12257 8067 12291
rect 9689 12257 9723 12291
rect 10149 12257 10183 12291
rect 11253 12257 11287 12291
rect 11713 12257 11747 12291
rect 13737 12257 13771 12291
rect 15761 12257 15795 12291
rect 6561 12189 6595 12223
rect 8401 12189 8435 12223
rect 10425 12189 10459 12223
rect 11069 12189 11103 12223
rect 11989 12189 12023 12223
rect 12817 12189 12851 12223
rect 15301 12189 15335 12223
rect 6358 12121 6392 12155
rect 7849 12121 7883 12155
rect 8171 12121 8205 12155
rect 2053 12053 2087 12087
rect 3893 12053 3927 12087
rect 6469 12053 6503 12087
rect 8309 12053 8343 12087
rect 14105 12053 14139 12087
rect 3525 11849 3559 11883
rect 6561 11849 6595 11883
rect 8585 11849 8619 11883
rect 9689 11849 9723 11883
rect 10149 11849 10183 11883
rect 11529 11849 11563 11883
rect 12173 11849 12207 11883
rect 15761 11849 15795 11883
rect 24731 11849 24765 11883
rect 2789 11781 2823 11815
rect 8217 11781 8251 11815
rect 14381 11781 14415 11815
rect 1869 11713 1903 11747
rect 3985 11713 4019 11747
rect 7665 11713 7699 11747
rect 9137 11713 9171 11747
rect 10609 11713 10643 11747
rect 13829 11713 13863 11747
rect 15301 11713 15335 11747
rect 4077 11645 4111 11679
rect 4905 11645 4939 11679
rect 5089 11645 5123 11679
rect 11897 11645 11931 11679
rect 12792 11645 12826 11679
rect 24660 11645 24694 11679
rect 1961 11577 1995 11611
rect 2513 11577 2547 11611
rect 7757 11577 7791 11611
rect 10971 11577 11005 11611
rect 13001 11577 13035 11611
rect 13645 11577 13679 11611
rect 13921 11577 13955 11611
rect 1685 11509 1719 11543
rect 3157 11509 3191 11543
rect 4169 11509 4203 11543
rect 5457 11509 5491 11543
rect 5917 11509 5951 11543
rect 6285 11509 6319 11543
rect 7113 11509 7147 11543
rect 7481 11509 7515 11543
rect 9045 11509 9079 11543
rect 10517 11509 10551 11543
rect 13185 11509 13219 11543
rect 25145 11509 25179 11543
rect 4537 11305 4571 11339
rect 7205 11305 7239 11339
rect 8585 11305 8619 11339
rect 10333 11305 10367 11339
rect 10793 11305 10827 11339
rect 12725 11305 12759 11339
rect 1961 11237 1995 11271
rect 2513 11237 2547 11271
rect 7481 11237 7515 11271
rect 8033 11237 8067 11271
rect 11758 11237 11792 11271
rect 13277 11237 13311 11271
rect 13369 11237 13403 11271
rect 4112 11169 4146 11203
rect 5641 11169 5675 11203
rect 5825 11169 5859 11203
rect 6193 11169 6227 11203
rect 9689 11169 9723 11203
rect 1869 11101 1903 11135
rect 6837 11101 6871 11135
rect 7389 11101 7423 11135
rect 9836 11101 9870 11135
rect 10057 11101 10091 11135
rect 11437 11101 11471 11135
rect 13553 11101 13587 11135
rect 2881 11033 2915 11067
rect 4215 11033 4249 11067
rect 9505 11033 9539 11067
rect 1685 10965 1719 10999
rect 3617 10965 3651 10999
rect 4997 10965 5031 10999
rect 6469 10965 6503 10999
rect 9965 10965 9999 10999
rect 11253 10965 11287 10999
rect 12357 10965 12391 10999
rect 13093 10965 13127 10999
rect 14197 10965 14231 10999
rect 2513 10761 2547 10795
rect 4537 10761 4571 10795
rect 9229 10761 9263 10795
rect 14473 10761 14507 10795
rect 8861 10693 8895 10727
rect 10149 10693 10183 10727
rect 14151 10693 14185 10727
rect 14289 10693 14323 10727
rect 3617 10625 3651 10659
rect 4261 10625 4295 10659
rect 6837 10625 6871 10659
rect 8953 10625 8987 10659
rect 9689 10625 9723 10659
rect 11253 10625 11287 10659
rect 14381 10625 14415 10659
rect 1593 10557 1627 10591
rect 3157 10557 3191 10591
rect 5733 10557 5767 10591
rect 7757 10557 7791 10591
rect 8732 10557 8766 10591
rect 10701 10557 10735 10591
rect 10977 10557 11011 10591
rect 3709 10489 3743 10523
rect 5089 10489 5123 10523
rect 7158 10489 7192 10523
rect 8585 10489 8619 10523
rect 12541 10489 12575 10523
rect 12633 10489 12667 10523
rect 13185 10489 13219 10523
rect 13553 10489 13587 10523
rect 14013 10489 14047 10523
rect 1961 10421 1995 10455
rect 2789 10421 2823 10455
rect 4997 10421 5031 10455
rect 6101 10421 6135 10455
rect 6653 10421 6687 10455
rect 8033 10421 8067 10455
rect 8493 10421 8527 10455
rect 11529 10421 11563 10455
rect 12265 10421 12299 10455
rect 13829 10421 13863 10455
rect 15577 10421 15611 10455
rect 2053 10217 2087 10251
rect 2973 10217 3007 10251
rect 3709 10217 3743 10251
rect 5733 10217 5767 10251
rect 6101 10217 6135 10251
rect 7665 10217 7699 10251
rect 8861 10217 8895 10251
rect 11345 10217 11379 10251
rect 12909 10217 12943 10251
rect 3433 10149 3467 10183
rect 4261 10149 4295 10183
rect 6469 10149 6503 10183
rect 7021 10149 7055 10183
rect 7849 10149 7883 10183
rect 11529 10149 11563 10183
rect 11621 10149 11655 10183
rect 13001 10149 13035 10183
rect 2329 10081 2363 10115
rect 2476 10081 2510 10115
rect 7389 10081 7423 10115
rect 8309 10081 8343 10115
rect 9873 10081 9907 10115
rect 10149 10081 10183 10115
rect 13093 10081 13127 10115
rect 15336 10081 15370 10115
rect 2697 10013 2731 10047
rect 4169 10013 4203 10047
rect 4813 10013 4847 10047
rect 6377 10013 6411 10047
rect 10333 10013 10367 10047
rect 11805 10013 11839 10047
rect 12541 10013 12575 10047
rect 1685 9877 1719 9911
rect 2605 9877 2639 9911
rect 5365 9877 5399 9911
rect 9413 9877 9447 9911
rect 10701 9877 10735 9911
rect 14105 9877 14139 9911
rect 15439 9877 15473 9911
rect 2697 9673 2731 9707
rect 3801 9673 3835 9707
rect 4077 9673 4111 9707
rect 4445 9673 4479 9707
rect 9781 9673 9815 9707
rect 12265 9673 12299 9707
rect 13461 9673 13495 9707
rect 15301 9673 15335 9707
rect 8861 9605 8895 9639
rect 2881 9537 2915 9571
rect 5917 9537 5951 9571
rect 6285 9537 6319 9571
rect 7205 9537 7239 9571
rect 8953 9537 8987 9571
rect 9321 9537 9355 9571
rect 10333 9537 10367 9571
rect 1685 9469 1719 9503
rect 5089 9469 5123 9503
rect 5273 9469 5307 9503
rect 8732 9469 8766 9503
rect 11253 9469 11287 9503
rect 12449 9469 12483 9503
rect 13001 9469 13035 9503
rect 13921 9469 13955 9503
rect 14105 9469 14139 9503
rect 16656 9469 16690 9503
rect 17049 9469 17083 9503
rect 1501 9401 1535 9435
rect 2053 9401 2087 9435
rect 6929 9401 6963 9435
rect 7021 9401 7055 9435
rect 8585 9401 8619 9435
rect 10654 9401 10688 9435
rect 11621 9401 11655 9435
rect 14013 9401 14047 9435
rect 2421 9333 2455 9367
rect 3249 9333 3283 9367
rect 8033 9333 8067 9367
rect 8401 9333 8435 9367
rect 10149 9333 10183 9367
rect 12541 9333 12575 9367
rect 16727 9333 16761 9367
rect 3525 9129 3559 9163
rect 4077 9129 4111 9163
rect 6469 9129 6503 9163
rect 6837 9129 6871 9163
rect 7941 9129 7975 9163
rect 8309 9129 8343 9163
rect 9045 9129 9079 9163
rect 10333 9129 10367 9163
rect 10701 9129 10735 9163
rect 12081 9129 12115 9163
rect 12725 9129 12759 9163
rect 1961 9061 1995 9095
rect 7342 9061 7376 9095
rect 11253 9061 11287 9095
rect 14933 9061 14967 9095
rect 5273 8993 5307 9027
rect 5549 8993 5583 9027
rect 5917 8993 5951 9027
rect 12909 8993 12943 9027
rect 13093 8993 13127 9027
rect 15301 8993 15335 9027
rect 1869 8925 1903 8959
rect 2513 8925 2547 8959
rect 2789 8925 2823 8959
rect 6193 8925 6227 8959
rect 7021 8925 7055 8959
rect 9873 8925 9907 8959
rect 11161 8925 11195 8959
rect 14197 8925 14231 8959
rect 15669 8925 15703 8959
rect 11713 8857 11747 8891
rect 15577 8857 15611 8891
rect 1593 8789 1627 8823
rect 3157 8789 3191 8823
rect 4905 8789 4939 8823
rect 8585 8789 8619 8823
rect 12449 8789 12483 8823
rect 15439 8789 15473 8823
rect 15761 8789 15795 8823
rect 4905 8585 4939 8619
rect 6009 8585 6043 8619
rect 8401 8585 8435 8619
rect 9321 8585 9355 8619
rect 10149 8585 10183 8619
rect 11621 8585 11655 8619
rect 11989 8585 12023 8619
rect 13001 8585 13035 8619
rect 14657 8585 14691 8619
rect 16221 8585 16255 8619
rect 16681 8585 16715 8619
rect 2513 8517 2547 8551
rect 4537 8517 4571 8551
rect 9045 8517 9079 8551
rect 9781 8517 9815 8551
rect 1777 8449 1811 8483
rect 3433 8449 3467 8483
rect 4353 8449 4387 8483
rect 9652 8449 9686 8483
rect 9873 8449 9907 8483
rect 13737 8449 13771 8483
rect 2973 8381 3007 8415
rect 3341 8381 3375 8415
rect 3525 8381 3559 8415
rect 1961 8313 1995 8347
rect 2053 8313 2087 8347
rect 5273 8381 5307 8415
rect 5549 8381 5583 8415
rect 6872 8381 6906 8415
rect 7297 8381 7331 8415
rect 8033 8381 8067 8415
rect 9505 8381 9539 8415
rect 10885 8381 10919 8415
rect 11136 8381 11170 8415
rect 14841 8381 14875 8415
rect 15393 8381 15427 8415
rect 16440 8381 16474 8415
rect 17233 8381 17267 8415
rect 6975 8313 7009 8347
rect 10517 8313 10551 8347
rect 13369 8313 13403 8347
rect 13461 8313 13495 8347
rect 4353 8245 4387 8279
rect 5089 8245 5123 8279
rect 6561 8245 6595 8279
rect 7849 8245 7883 8279
rect 11207 8245 11241 8279
rect 12725 8245 12759 8279
rect 14933 8245 14967 8279
rect 15853 8245 15887 8279
rect 16865 8245 16899 8279
rect 2145 8041 2179 8075
rect 2697 8041 2731 8075
rect 3065 8041 3099 8075
rect 7481 8041 7515 8075
rect 11161 8041 11195 8075
rect 12357 8041 12391 8075
rect 13737 8041 13771 8075
rect 15393 8041 15427 8075
rect 8033 7973 8067 8007
rect 3341 7905 3375 7939
rect 5365 7905 5399 7939
rect 5825 7905 5859 7939
rect 6561 7905 6595 7939
rect 9873 7905 9907 7939
rect 11989 7905 12023 7939
rect 15301 7905 15335 7939
rect 15853 7905 15887 7939
rect 1777 7837 1811 7871
rect 4721 7837 4755 7871
rect 7205 7837 7239 7871
rect 8401 7837 8435 7871
rect 10517 7837 10551 7871
rect 13921 7837 13955 7871
rect 8309 7769 8343 7803
rect 1685 7701 1719 7735
rect 3709 7701 3743 7735
rect 8171 7701 8205 7735
rect 8493 7701 8527 7735
rect 12909 7701 12943 7735
rect 13277 7701 13311 7735
rect 15025 7701 15059 7735
rect 4077 7497 4111 7531
rect 10609 7497 10643 7531
rect 13737 7497 13771 7531
rect 11805 7429 11839 7463
rect 12173 7429 12207 7463
rect 2697 7361 2731 7395
rect 5089 7361 5123 7395
rect 5549 7361 5583 7395
rect 10885 7361 10919 7395
rect 11529 7361 11563 7395
rect 12449 7361 12483 7395
rect 14289 7361 14323 7395
rect 14565 7361 14599 7395
rect 1444 7293 1478 7327
rect 1869 7293 1903 7327
rect 7757 7293 7791 7327
rect 9045 7293 9079 7327
rect 16037 7293 16071 7327
rect 16313 7293 16347 7327
rect 1547 7225 1581 7259
rect 3018 7225 3052 7259
rect 4537 7225 4571 7259
rect 4905 7225 4939 7259
rect 5181 7225 5215 7259
rect 8217 7225 8251 7259
rect 9407 7225 9441 7259
rect 10977 7225 11011 7259
rect 12770 7225 12804 7259
rect 14105 7225 14139 7259
rect 14381 7225 14415 7259
rect 15393 7225 15427 7259
rect 16773 7225 16807 7259
rect 2513 7157 2547 7191
rect 3617 7157 3651 7191
rect 6561 7157 6595 7191
rect 7297 7157 7331 7191
rect 8585 7157 8619 7191
rect 8861 7157 8895 7191
rect 9965 7157 9999 7191
rect 10241 7157 10275 7191
rect 13369 7157 13403 7191
rect 15853 7157 15887 7191
rect 2329 6953 2363 6987
rect 3433 6953 3467 6987
rect 5825 6953 5859 6987
rect 8125 6953 8159 6987
rect 8493 6953 8527 6987
rect 10885 6953 10919 6987
rect 11989 6953 12023 6987
rect 13093 6953 13127 6987
rect 14749 6953 14783 6987
rect 17509 6953 17543 6987
rect 24731 6953 24765 6987
rect 2605 6885 2639 6919
rect 4721 6885 4755 6919
rect 5267 6885 5301 6919
rect 6837 6885 6871 6919
rect 9873 6885 9907 6919
rect 10425 6885 10459 6919
rect 13829 6885 13863 6919
rect 14381 6885 14415 6919
rect 9137 6817 9171 6851
rect 12173 6817 12207 6851
rect 15301 6817 15335 6851
rect 15448 6817 15482 6851
rect 16865 6817 16899 6851
rect 17012 6817 17046 6851
rect 24644 6817 24678 6851
rect 1409 6749 1443 6783
rect 2513 6749 2547 6783
rect 3157 6749 3191 6783
rect 4905 6749 4939 6783
rect 6745 6749 6779 6783
rect 8585 6749 8619 6783
rect 9781 6749 9815 6783
rect 13737 6749 13771 6783
rect 15025 6749 15059 6783
rect 15669 6749 15703 6783
rect 17233 6749 17267 6783
rect 7297 6681 7331 6715
rect 1961 6613 1995 6647
rect 7757 6613 7791 6647
rect 12357 6613 12391 6647
rect 13461 6613 13495 6647
rect 15577 6613 15611 6647
rect 15945 6613 15979 6647
rect 16313 6613 16347 6647
rect 17141 6613 17175 6647
rect 2973 6409 3007 6443
rect 4629 6409 4663 6443
rect 6285 6409 6319 6443
rect 9781 6409 9815 6443
rect 11897 6409 11931 6443
rect 12265 6409 12299 6443
rect 13645 6409 13679 6443
rect 14473 6409 14507 6443
rect 15485 6409 15519 6443
rect 15577 6409 15611 6443
rect 17601 6409 17635 6443
rect 24685 6409 24719 6443
rect 4261 6341 4295 6375
rect 8033 6341 8067 6375
rect 3249 6273 3283 6307
rect 3525 6273 3559 6307
rect 4813 6273 4847 6307
rect 5457 6273 5491 6307
rect 10333 6273 10367 6307
rect 11345 6273 11379 6307
rect 13369 6273 13403 6307
rect 17233 6341 17267 6375
rect 16865 6273 16899 6307
rect 1869 6205 1903 6239
rect 2145 6205 2179 6239
rect 7021 6205 7055 6239
rect 7665 6205 7699 6239
rect 8217 6205 8251 6239
rect 14105 6205 14139 6239
rect 14289 6205 14323 6239
rect 15209 6205 15243 6239
rect 15485 6205 15519 6239
rect 15761 6205 15795 6239
rect 16313 6205 16347 6239
rect 18924 6205 18958 6239
rect 19349 6205 19383 6239
rect 3341 6137 3375 6171
rect 4905 6137 4939 6171
rect 6561 6137 6595 6171
rect 6837 6137 6871 6171
rect 8538 6137 8572 6171
rect 10057 6137 10091 6171
rect 10149 6137 10183 6171
rect 12725 6137 12759 6171
rect 12817 6137 12851 6171
rect 1685 6069 1719 6103
rect 2697 6069 2731 6103
rect 5825 6069 5859 6103
rect 7113 6069 7147 6103
rect 9137 6069 9171 6103
rect 9505 6069 9539 6103
rect 10977 6069 11011 6103
rect 15853 6069 15887 6103
rect 19027 6069 19061 6103
rect 1547 5865 1581 5899
rect 1961 5865 1995 5899
rect 3525 5865 3559 5899
rect 5273 5865 5307 5899
rect 6653 5865 6687 5899
rect 7297 5865 7331 5899
rect 9873 5865 9907 5899
rect 13737 5865 13771 5899
rect 14749 5865 14783 5899
rect 15577 5865 15611 5899
rect 16313 5865 16347 5899
rect 17325 5865 17359 5899
rect 6095 5797 6129 5831
rect 8217 5797 8251 5831
rect 8769 5797 8803 5831
rect 10057 5797 10091 5831
rect 12725 5797 12759 5831
rect 12817 5797 12851 5831
rect 14473 5797 14507 5831
rect 1444 5729 1478 5763
rect 3065 5729 3099 5763
rect 4721 5729 4755 5763
rect 4905 5729 4939 5763
rect 9045 5729 9079 5763
rect 11253 5729 11287 5763
rect 11529 5729 11563 5763
rect 14264 5729 14298 5763
rect 15669 5729 15703 5763
rect 20913 5729 20947 5763
rect 2421 5661 2455 5695
rect 5733 5661 5767 5695
rect 8125 5661 8159 5695
rect 11805 5661 11839 5695
rect 13001 5661 13035 5695
rect 16865 5661 16899 5695
rect 15117 5593 15151 5627
rect 2237 5525 2271 5559
rect 6929 5525 6963 5559
rect 10793 5525 10827 5559
rect 12449 5525 12483 5559
rect 21097 5525 21131 5559
rect 2973 5321 3007 5355
rect 8815 5321 8849 5355
rect 9321 5321 9355 5355
rect 12265 5321 12299 5355
rect 13645 5321 13679 5355
rect 13921 5321 13955 5355
rect 15393 5321 15427 5355
rect 20913 5321 20947 5355
rect 8217 5253 8251 5287
rect 8953 5253 8987 5287
rect 9689 5253 9723 5287
rect 2053 5185 2087 5219
rect 3157 5185 3191 5219
rect 6929 5185 6963 5219
rect 7297 5185 7331 5219
rect 8401 5185 8435 5219
rect 9045 5185 9079 5219
rect 11529 5185 11563 5219
rect 12449 5185 12483 5219
rect 1869 5117 1903 5151
rect 2145 5117 2179 5151
rect 3617 5117 3651 5151
rect 4169 5117 4203 5151
rect 5549 5117 5583 5151
rect 2697 5049 2731 5083
rect 5917 5049 5951 5083
rect 6561 5049 6595 5083
rect 7021 5049 7055 5083
rect 8677 5117 8711 5151
rect 10701 5117 10735 5151
rect 11069 5117 11103 5151
rect 11253 5117 11287 5151
rect 13461 5117 13495 5151
rect 12770 5049 12804 5083
rect 4629 4981 4663 5015
rect 4997 4981 5031 5015
rect 6285 4981 6319 5015
rect 8401 4981 8435 5015
rect 8493 4981 8527 5015
rect 11805 4981 11839 5015
rect 13369 4981 13403 5015
rect 13461 4981 13495 5015
rect 20085 5253 20119 5287
rect 14105 5185 14139 5219
rect 14473 5117 14507 5151
rect 14749 5117 14783 5151
rect 15853 5117 15887 5151
rect 16773 5117 16807 5151
rect 18096 5117 18130 5151
rect 18521 5117 18555 5151
rect 19901 5117 19935 5151
rect 20453 5117 20487 5151
rect 15761 5049 15795 5083
rect 13921 4981 13955 5015
rect 14289 4981 14323 5015
rect 18199 4981 18233 5015
rect 2237 4777 2271 4811
rect 3065 4777 3099 4811
rect 4997 4777 5031 4811
rect 6009 4777 6043 4811
rect 9045 4777 9079 4811
rect 9873 4777 9907 4811
rect 11345 4777 11379 4811
rect 12725 4777 12759 4811
rect 14565 4777 14599 4811
rect 15393 4777 15427 4811
rect 1961 4709 1995 4743
rect 2421 4709 2455 4743
rect 3433 4709 3467 4743
rect 6469 4709 6503 4743
rect 10517 4709 10551 4743
rect 13277 4709 13311 4743
rect 1409 4641 1443 4675
rect 1547 4641 1581 4675
rect 5181 4641 5215 4675
rect 5365 4641 5399 4675
rect 6808 4641 6842 4675
rect 8309 4641 8343 4675
rect 8493 4641 8527 4675
rect 11989 4641 12023 4675
rect 15301 4641 15335 4675
rect 15761 4641 15795 4675
rect 16865 4641 16899 4675
rect 18705 4641 18739 4675
rect 2789 4573 2823 4607
rect 8769 4573 8803 4607
rect 10425 4573 10459 4607
rect 11069 4573 11103 4607
rect 13185 4573 13219 4607
rect 13461 4573 13495 4607
rect 14289 4573 14323 4607
rect 2586 4505 2620 4539
rect 12173 4505 12207 4539
rect 17049 4505 17083 4539
rect 2697 4437 2731 4471
rect 3801 4437 3835 4471
rect 4629 4437 4663 4471
rect 6607 4437 6641 4471
rect 6745 4437 6779 4471
rect 6929 4437 6963 4471
rect 7849 4437 7883 4471
rect 16405 4437 16439 4471
rect 18889 4437 18923 4471
rect 1685 4233 1719 4267
rect 3065 4233 3099 4267
rect 4077 4233 4111 4267
rect 6377 4233 6411 4267
rect 6653 4233 6687 4267
rect 10793 4233 10827 4267
rect 18889 4233 18923 4267
rect 4445 4165 4479 4199
rect 4767 4165 4801 4199
rect 4905 4165 4939 4199
rect 5641 4165 5675 4199
rect 4997 4097 5031 4131
rect 5549 4097 5583 4131
rect 6193 4097 6227 4131
rect 1501 4029 1535 4063
rect 2973 4029 3007 4063
rect 3709 4029 3743 4063
rect 4629 3961 4663 3995
rect 5549 3961 5583 3995
rect 9413 4165 9447 4199
rect 9505 4165 9539 4199
rect 11069 4165 11103 4199
rect 11897 4165 11931 4199
rect 12265 4165 12299 4199
rect 14105 4165 14139 4199
rect 16773 4165 16807 4199
rect 6837 4097 6871 4131
rect 8125 4029 8159 4063
rect 8677 4029 8711 4063
rect 9137 4029 9171 4063
rect 9781 4097 9815 4131
rect 12817 4097 12851 4131
rect 14933 4097 14967 4131
rect 16221 4097 16255 4131
rect 18199 4097 18233 4131
rect 11253 4029 11287 4063
rect 12633 4029 12667 4063
rect 13737 4029 13771 4063
rect 18096 4029 18130 4063
rect 18521 4029 18555 4063
rect 19140 4029 19174 4063
rect 7297 3961 7331 3995
rect 8861 3961 8895 3995
rect 9413 3961 9447 3995
rect 9873 3961 9907 3995
rect 10425 3961 10459 3995
rect 13138 3961 13172 3995
rect 14657 3961 14691 3995
rect 14749 3961 14783 3995
rect 16037 3961 16071 3995
rect 16313 3961 16347 3995
rect 19533 3961 19567 3995
rect 2421 3893 2455 3927
rect 2789 3893 2823 3927
rect 5273 3893 5307 3927
rect 6653 3893 6687 3927
rect 7941 3893 7975 3927
rect 11391 3893 11425 3927
rect 14381 3893 14415 3927
rect 15669 3893 15703 3927
rect 17233 3893 17267 3927
rect 19211 3893 19245 3927
rect 1869 3689 1903 3723
rect 3525 3689 3559 3723
rect 4215 3689 4249 3723
rect 5089 3689 5123 3723
rect 6469 3689 6503 3723
rect 8033 3689 8067 3723
rect 8493 3689 8527 3723
rect 9413 3689 9447 3723
rect 10609 3689 10643 3723
rect 12817 3689 12851 3723
rect 13369 3689 13403 3723
rect 13921 3689 13955 3723
rect 3893 3621 3927 3655
rect 5594 3621 5628 3655
rect 7205 3621 7239 3655
rect 10051 3621 10085 3655
rect 11529 3621 11563 3655
rect 11621 3621 11655 3655
rect 12541 3621 12575 3655
rect 15485 3621 15519 3655
rect 18429 3621 18463 3655
rect 1444 3553 1478 3587
rect 2237 3553 2271 3587
rect 3065 3553 3099 3587
rect 4144 3553 4178 3587
rect 6193 3553 6227 3587
rect 8585 3553 8619 3587
rect 16957 3553 16991 3587
rect 19073 3553 19107 3587
rect 3157 3485 3191 3519
rect 5273 3485 5307 3519
rect 7113 3485 7147 3519
rect 7573 3485 7607 3519
rect 9689 3485 9723 3519
rect 11805 3485 11839 3519
rect 13001 3485 13035 3519
rect 15393 3485 15427 3519
rect 16865 3485 16899 3519
rect 1547 3417 1581 3451
rect 4629 3417 4663 3451
rect 11345 3417 11379 3451
rect 15945 3417 15979 3451
rect 16405 3417 16439 3451
rect 6929 3349 6963 3383
rect 8723 3349 8757 3383
rect 9045 3349 9079 3383
rect 14657 3349 14691 3383
rect 2513 3145 2547 3179
rect 2973 3145 3007 3179
rect 4905 3145 4939 3179
rect 6193 3145 6227 3179
rect 6561 3145 6595 3179
rect 7849 3145 7883 3179
rect 8861 3145 8895 3179
rect 9229 3145 9263 3179
rect 11069 3145 11103 3179
rect 12265 3145 12299 3179
rect 13093 3145 13127 3179
rect 14565 3145 14599 3179
rect 14841 3145 14875 3179
rect 15025 3145 15059 3179
rect 15669 3145 15703 3179
rect 16221 3145 16255 3179
rect 17325 3145 17359 3179
rect 19763 3145 19797 3179
rect 4537 3077 4571 3111
rect 8217 3077 8251 3111
rect 10333 3077 10367 3111
rect 1869 3009 1903 3043
rect 4169 3009 4203 3043
rect 8401 3009 8435 3043
rect 9413 3009 9447 3043
rect 15301 3077 15335 3111
rect 19073 3077 19107 3111
rect 16405 3009 16439 3043
rect 16681 3009 16715 3043
rect 18061 3009 18095 3043
rect 1501 2941 1535 2975
rect 2237 2941 2271 2975
rect 3525 2941 3559 2975
rect 3893 2941 3927 2975
rect 4997 2941 5031 2975
rect 11161 2941 11195 2975
rect 12725 2941 12759 2975
rect 13369 2941 13403 2975
rect 14841 2941 14875 2975
rect 15117 2941 15151 2975
rect 18153 2941 18187 2975
rect 19660 2941 19694 2975
rect 20085 2941 20119 2975
rect 20704 2941 20738 2975
rect 24384 2941 24418 2975
rect 3249 2873 3283 2907
rect 5318 2873 5352 2907
rect 6929 2873 6963 2907
rect 7021 2873 7055 2907
rect 7573 2873 7607 2907
rect 9734 2873 9768 2907
rect 13690 2873 13724 2907
rect 16497 2873 16531 2907
rect 17785 2873 17819 2907
rect 21189 2873 21223 2907
rect 5917 2805 5951 2839
rect 11345 2805 11379 2839
rect 11805 2805 11839 2839
rect 14289 2805 14323 2839
rect 20775 2805 20809 2839
rect 24455 2805 24489 2839
rect 24869 2805 24903 2839
rect 1547 2601 1581 2635
rect 3525 2601 3559 2635
rect 4537 2601 4571 2635
rect 6377 2601 6411 2635
rect 6653 2601 6687 2635
rect 8309 2601 8343 2635
rect 9505 2601 9539 2635
rect 9965 2601 9999 2635
rect 12357 2601 12391 2635
rect 13369 2601 13403 2635
rect 15945 2601 15979 2635
rect 18061 2601 18095 2635
rect 21327 2601 21361 2635
rect 5457 2533 5491 2567
rect 7021 2533 7055 2567
rect 7113 2533 7147 2567
rect 7941 2533 7975 2567
rect 10517 2533 10551 2567
rect 11069 2533 11103 2567
rect 11713 2533 11747 2567
rect 14013 2533 14047 2567
rect 14933 2533 14967 2567
rect 16313 2533 16347 2567
rect 18337 2533 18371 2567
rect 23489 2533 23523 2567
rect 1476 2465 1510 2499
rect 3065 2465 3099 2499
rect 3801 2465 3835 2499
rect 4328 2465 4362 2499
rect 8493 2465 8527 2499
rect 12633 2465 12667 2499
rect 14565 2465 14599 2499
rect 15301 2465 15335 2499
rect 18429 2465 18463 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 21256 2465 21290 2499
rect 23004 2465 23038 2499
rect 24660 2465 24694 2499
rect 3157 2397 3191 2431
rect 5089 2397 5123 2431
rect 5365 2397 5399 2431
rect 10425 2397 10459 2431
rect 11437 2397 11471 2431
rect 13921 2397 13955 2431
rect 16221 2397 16255 2431
rect 16681 2397 16715 2431
rect 17233 2397 17267 2431
rect 21649 2397 21683 2431
rect 2329 2329 2363 2363
rect 7573 2329 7607 2363
rect 8677 2329 8711 2363
rect 12817 2329 12851 2363
rect 24731 2329 24765 2363
rect 1961 2261 1995 2295
rect 4813 2261 4847 2295
rect 6101 2261 6135 2295
rect 9045 2261 9079 2295
rect 20085 2261 20119 2295
rect 23075 2261 23109 2295
rect 25145 2261 25179 2295
<< metal1 >>
rect 7742 27480 7748 27532
rect 7800 27520 7806 27532
rect 8846 27520 8852 27532
rect 7800 27492 8852 27520
rect 7800 27480 7806 27492
rect 8846 27480 8852 27492
rect 8904 27480 8910 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 16850 24392 16856 24404
rect 15519 24364 16856 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 16850 24352 16856 24364
rect 16908 24352 16914 24404
rect 2777 24259 2835 24265
rect 2777 24225 2789 24259
rect 2823 24256 2835 24259
rect 2866 24256 2872 24268
rect 2823 24228 2872 24256
rect 2823 24225 2835 24228
rect 2777 24219 2835 24225
rect 2866 24216 2872 24228
rect 2924 24216 2930 24268
rect 11974 24265 11980 24268
rect 11952 24259 11980 24265
rect 11952 24256 11964 24259
rect 11887 24228 11964 24256
rect 11952 24225 11964 24228
rect 12032 24256 12038 24268
rect 12526 24256 12532 24268
rect 12032 24228 12532 24256
rect 11952 24219 11980 24225
rect 11974 24216 11980 24219
rect 12032 24216 12038 24228
rect 12526 24216 12532 24228
rect 12584 24216 12590 24268
rect 12964 24259 13022 24265
rect 12964 24225 12976 24259
rect 13010 24256 13022 24259
rect 13446 24256 13452 24268
rect 13010 24228 13452 24256
rect 13010 24225 13022 24228
rect 12964 24219 13022 24225
rect 13446 24216 13452 24228
rect 13504 24216 13510 24268
rect 15289 24259 15347 24265
rect 15289 24225 15301 24259
rect 15335 24256 15347 24259
rect 15838 24256 15844 24268
rect 15335 24228 15844 24256
rect 15335 24225 15347 24228
rect 15289 24219 15347 24225
rect 15838 24216 15844 24228
rect 15896 24216 15902 24268
rect 24670 24265 24676 24268
rect 24648 24259 24676 24265
rect 24648 24256 24660 24259
rect 24583 24228 24660 24256
rect 24648 24225 24660 24228
rect 24728 24256 24734 24268
rect 26878 24256 26884 24268
rect 24728 24228 26884 24256
rect 24648 24219 24676 24225
rect 24670 24216 24676 24219
rect 24728 24216 24734 24228
rect 26878 24216 26884 24228
rect 26936 24216 26942 24268
rect 12529 24123 12587 24129
rect 12529 24089 12541 24123
rect 12575 24120 12587 24123
rect 12710 24120 12716 24132
rect 12575 24092 12716 24120
rect 12575 24089 12587 24092
rect 12529 24083 12587 24089
rect 12710 24080 12716 24092
rect 12768 24080 12774 24132
rect 2915 24055 2973 24061
rect 2915 24021 2927 24055
rect 2961 24052 2973 24055
rect 3602 24052 3608 24064
rect 2961 24024 3608 24052
rect 2961 24021 2973 24024
rect 2915 24015 2973 24021
rect 3602 24012 3608 24024
rect 3660 24012 3666 24064
rect 12023 24055 12081 24061
rect 12023 24021 12035 24055
rect 12069 24052 12081 24055
rect 12342 24052 12348 24064
rect 12069 24024 12348 24052
rect 12069 24021 12081 24024
rect 12023 24015 12081 24021
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 12618 24012 12624 24064
rect 12676 24052 12682 24064
rect 13035 24055 13093 24061
rect 13035 24052 13047 24055
rect 12676 24024 13047 24052
rect 12676 24012 12682 24024
rect 13035 24021 13047 24024
rect 13081 24021 13093 24055
rect 13035 24015 13093 24021
rect 20622 24012 20628 24064
rect 20680 24052 20686 24064
rect 24719 24055 24777 24061
rect 24719 24052 24731 24055
rect 20680 24024 24731 24052
rect 20680 24012 20686 24024
rect 24719 24021 24731 24024
rect 24765 24021 24777 24055
rect 24719 24015 24777 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2866 23848 2872 23860
rect 2827 23820 2872 23848
rect 2866 23808 2872 23820
rect 2924 23808 2930 23860
rect 3142 23848 3148 23860
rect 3103 23820 3148 23848
rect 3142 23808 3148 23820
rect 3200 23808 3206 23860
rect 4798 23848 4804 23860
rect 4759 23820 4804 23848
rect 4798 23808 4804 23820
rect 4856 23808 4862 23860
rect 7006 23848 7012 23860
rect 6967 23820 7012 23848
rect 7006 23808 7012 23820
rect 7064 23808 7070 23860
rect 9769 23851 9827 23857
rect 9769 23817 9781 23851
rect 9815 23848 9827 23851
rect 10870 23848 10876 23860
rect 9815 23820 10876 23848
rect 9815 23817 9827 23820
rect 9769 23811 9827 23817
rect 10870 23808 10876 23820
rect 10928 23808 10934 23860
rect 11974 23848 11980 23860
rect 11935 23820 11980 23848
rect 11974 23808 11980 23820
rect 12032 23808 12038 23860
rect 13446 23848 13452 23860
rect 13407 23820 13452 23848
rect 13446 23808 13452 23820
rect 13504 23848 13510 23860
rect 14826 23848 14832 23860
rect 13504 23820 14832 23848
rect 13504 23808 13510 23820
rect 14826 23808 14832 23820
rect 14884 23808 14890 23860
rect 15838 23848 15844 23860
rect 15799 23820 15844 23848
rect 15838 23808 15844 23820
rect 15896 23848 15902 23860
rect 16482 23848 16488 23860
rect 15896 23820 16488 23848
rect 15896 23808 15902 23820
rect 16482 23808 16488 23820
rect 16540 23808 16546 23860
rect 17037 23851 17095 23857
rect 17037 23817 17049 23851
rect 17083 23848 17095 23851
rect 18874 23848 18880 23860
rect 17083 23820 18880 23848
rect 17083 23817 17095 23820
rect 17037 23811 17095 23817
rect 18874 23808 18880 23820
rect 18932 23808 18938 23860
rect 19521 23851 19579 23857
rect 19521 23817 19533 23851
rect 19567 23848 19579 23851
rect 20898 23848 20904 23860
rect 19567 23820 20904 23848
rect 19567 23817 19579 23820
rect 19521 23811 19579 23817
rect 3418 23740 3424 23792
rect 3476 23780 3482 23792
rect 4387 23783 4445 23789
rect 4387 23780 4399 23783
rect 3476 23752 4399 23780
rect 3476 23740 3482 23752
rect 4387 23749 4399 23752
rect 4433 23749 4445 23783
rect 19107 23783 19165 23789
rect 19107 23780 19119 23783
rect 4387 23743 4445 23749
rect 12544 23752 19119 23780
rect 8294 23672 8300 23724
rect 8352 23712 8358 23724
rect 12544 23721 12572 23752
rect 19107 23749 19119 23752
rect 19153 23749 19165 23783
rect 19107 23743 19165 23749
rect 9033 23715 9091 23721
rect 9033 23712 9045 23715
rect 8352 23684 9045 23712
rect 8352 23672 8358 23684
rect 934 23604 940 23656
rect 992 23644 998 23656
rect 1432 23647 1490 23653
rect 1432 23644 1444 23647
rect 992 23616 1444 23644
rect 992 23604 998 23616
rect 1432 23613 1444 23616
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1432 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 2961 23647 3019 23653
rect 2961 23613 2973 23647
rect 3007 23644 3019 23647
rect 4316 23647 4374 23653
rect 3007 23616 3648 23644
rect 3007 23613 3019 23616
rect 2961 23607 3019 23613
rect 1302 23468 1308 23520
rect 1360 23508 1366 23520
rect 3620 23517 3648 23616
rect 4316 23613 4328 23647
rect 4362 23644 4374 23647
rect 4798 23644 4804 23656
rect 4362 23616 4804 23644
rect 4362 23613 4374 23616
rect 4316 23607 4374 23613
rect 4798 23604 4804 23616
rect 4856 23604 4862 23656
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 7377 23647 7435 23653
rect 7377 23644 7389 23647
rect 6871 23616 7389 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 7377 23613 7389 23616
rect 7423 23644 7435 23647
rect 7466 23644 7472 23656
rect 7423 23616 7472 23644
rect 7423 23613 7435 23616
rect 7377 23607 7435 23613
rect 7466 23604 7472 23616
rect 7524 23604 7530 23656
rect 8655 23653 8683 23684
rect 9033 23681 9045 23684
rect 9079 23681 9091 23715
rect 9033 23675 9091 23681
rect 11609 23715 11667 23721
rect 11609 23681 11621 23715
rect 11655 23712 11667 23715
rect 12529 23715 12587 23721
rect 12529 23712 12541 23715
rect 11655 23684 12541 23712
rect 11655 23681 11667 23684
rect 11609 23675 11667 23681
rect 12529 23681 12541 23684
rect 12575 23681 12587 23715
rect 12802 23712 12808 23724
rect 12763 23684 12808 23712
rect 12529 23675 12587 23681
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 8640 23647 8698 23653
rect 8640 23613 8652 23647
rect 8686 23613 8698 23647
rect 8640 23607 8698 23613
rect 9585 23647 9643 23653
rect 9585 23613 9597 23647
rect 9631 23644 9643 23647
rect 10134 23644 10140 23656
rect 9631 23616 10140 23644
rect 9631 23613 9643 23616
rect 9585 23607 9643 23613
rect 10134 23604 10140 23616
rect 10192 23604 10198 23656
rect 16850 23644 16856 23656
rect 16763 23616 16856 23644
rect 16850 23604 16856 23616
rect 16908 23644 16914 23656
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 16908 23616 17417 23644
rect 16908 23604 16914 23616
rect 17405 23613 17417 23616
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 19036 23647 19094 23653
rect 19036 23613 19048 23647
rect 19082 23644 19094 23647
rect 19536 23644 19564 23811
rect 20898 23808 20904 23820
rect 20956 23808 20962 23860
rect 21453 23851 21511 23857
rect 21453 23817 21465 23851
rect 21499 23848 21511 23851
rect 22830 23848 22836 23860
rect 21499 23820 22836 23848
rect 21499 23817 21511 23820
rect 21453 23811 21511 23817
rect 19082 23616 19564 23644
rect 20968 23647 21026 23653
rect 19082 23613 19094 23616
rect 19036 23607 19094 23613
rect 20968 23613 20980 23647
rect 21014 23644 21026 23647
rect 21468 23644 21496 23811
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 24581 23851 24639 23857
rect 24581 23817 24593 23851
rect 24627 23848 24639 23851
rect 24670 23848 24676 23860
rect 24627 23820 24676 23848
rect 24627 23817 24639 23820
rect 24581 23811 24639 23817
rect 24670 23808 24676 23820
rect 24728 23808 24734 23860
rect 25222 23848 25228 23860
rect 25183 23820 25228 23848
rect 25222 23808 25228 23820
rect 25280 23808 25286 23860
rect 24213 23783 24271 23789
rect 24213 23749 24225 23783
rect 24259 23780 24271 23783
rect 24854 23780 24860 23792
rect 24259 23752 24860 23780
rect 24259 23749 24271 23752
rect 24213 23743 24271 23749
rect 21014 23616 21496 23644
rect 23728 23647 23786 23653
rect 21014 23613 21026 23616
rect 20968 23607 21026 23613
rect 23728 23613 23740 23647
rect 23774 23644 23786 23647
rect 24228 23644 24256 23743
rect 24854 23740 24860 23752
rect 24912 23740 24918 23792
rect 23774 23616 24256 23644
rect 24740 23647 24798 23653
rect 23774 23613 23786 23616
rect 23728 23607 23786 23613
rect 24740 23613 24752 23647
rect 24786 23644 24798 23647
rect 25222 23644 25228 23656
rect 24786 23616 25228 23644
rect 24786 23613 24798 23616
rect 24740 23607 24798 23613
rect 25222 23604 25228 23616
rect 25280 23604 25286 23656
rect 12621 23579 12679 23585
rect 12621 23545 12633 23579
rect 12667 23576 12679 23579
rect 12710 23576 12716 23588
rect 12667 23548 12716 23576
rect 12667 23545 12679 23548
rect 12621 23539 12679 23545
rect 1535 23511 1593 23517
rect 1535 23508 1547 23511
rect 1360 23480 1547 23508
rect 1360 23468 1366 23480
rect 1535 23477 1547 23480
rect 1581 23477 1593 23511
rect 1535 23471 1593 23477
rect 3605 23511 3663 23517
rect 3605 23477 3617 23511
rect 3651 23508 3663 23511
rect 4062 23508 4068 23520
rect 3651 23480 4068 23508
rect 3651 23477 3663 23480
rect 3605 23471 3663 23477
rect 4062 23468 4068 23480
rect 4120 23468 4126 23520
rect 8711 23511 8769 23517
rect 8711 23477 8723 23511
rect 8757 23508 8769 23511
rect 8846 23508 8852 23520
rect 8757 23480 8852 23508
rect 8757 23477 8769 23480
rect 8711 23471 8769 23477
rect 8846 23468 8852 23480
rect 8904 23468 8910 23520
rect 12434 23468 12440 23520
rect 12492 23508 12498 23520
rect 12636 23508 12664 23539
rect 12710 23536 12716 23548
rect 12768 23536 12774 23588
rect 14918 23576 14924 23588
rect 14879 23548 14924 23576
rect 14918 23536 14924 23548
rect 14976 23536 14982 23588
rect 15013 23579 15071 23585
rect 15013 23545 15025 23579
rect 15059 23545 15071 23579
rect 15562 23576 15568 23588
rect 15523 23548 15568 23576
rect 15013 23539 15071 23545
rect 14734 23508 14740 23520
rect 12492 23480 12664 23508
rect 14647 23480 14740 23508
rect 12492 23468 12498 23480
rect 14734 23468 14740 23480
rect 14792 23508 14798 23520
rect 15028 23508 15056 23539
rect 15562 23536 15568 23548
rect 15620 23536 15626 23588
rect 14792 23480 15056 23508
rect 14792 23468 14798 23480
rect 20070 23468 20076 23520
rect 20128 23508 20134 23520
rect 21039 23511 21097 23517
rect 21039 23508 21051 23511
rect 20128 23480 21051 23508
rect 20128 23468 20134 23480
rect 21039 23477 21051 23480
rect 21085 23477 21097 23511
rect 21039 23471 21097 23477
rect 22738 23468 22744 23520
rect 22796 23508 22802 23520
rect 23799 23511 23857 23517
rect 23799 23508 23811 23511
rect 22796 23480 23811 23508
rect 22796 23468 22802 23480
rect 23799 23477 23811 23480
rect 23845 23477 23857 23511
rect 23799 23471 23857 23477
rect 24578 23468 24584 23520
rect 24636 23508 24642 23520
rect 24811 23511 24869 23517
rect 24811 23508 24823 23511
rect 24636 23480 24823 23508
rect 24636 23468 24642 23480
rect 24811 23477 24823 23480
rect 24857 23477 24869 23511
rect 24811 23471 24869 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 7466 23264 7472 23316
rect 7524 23304 7530 23316
rect 11655 23307 11713 23313
rect 11655 23304 11667 23307
rect 7524 23276 11667 23304
rect 7524 23264 7530 23276
rect 11655 23273 11667 23276
rect 11701 23273 11713 23307
rect 11655 23267 11713 23273
rect 12250 23264 12256 23316
rect 12308 23304 12314 23316
rect 14918 23304 14924 23316
rect 12308 23276 12756 23304
rect 14879 23276 14924 23304
rect 12308 23264 12314 23276
rect 8711 23239 8769 23245
rect 8711 23205 8723 23239
rect 8757 23236 8769 23239
rect 12618 23236 12624 23248
rect 8757 23208 12624 23236
rect 8757 23205 8769 23208
rect 8711 23199 8769 23205
rect 12618 23196 12624 23208
rect 12676 23196 12682 23248
rect 12728 23245 12756 23276
rect 14918 23264 14924 23276
rect 14976 23264 14982 23316
rect 12713 23239 12771 23245
rect 12713 23205 12725 23239
rect 12759 23205 12771 23239
rect 15470 23236 15476 23248
rect 15431 23208 15476 23236
rect 12713 23199 12771 23205
rect 15470 23196 15476 23208
rect 15528 23196 15534 23248
rect 11517 23171 11575 23177
rect 11517 23137 11529 23171
rect 11563 23168 11575 23171
rect 11606 23168 11612 23180
rect 11563 23140 11612 23168
rect 11563 23137 11575 23140
rect 11517 23131 11575 23137
rect 11606 23128 11612 23140
rect 11664 23128 11670 23180
rect 12621 23103 12679 23109
rect 12621 23069 12633 23103
rect 12667 23100 12679 23103
rect 13078 23100 13084 23112
rect 12667 23072 13084 23100
rect 12667 23069 12679 23072
rect 12621 23063 12679 23069
rect 13078 23060 13084 23072
rect 13136 23060 13142 23112
rect 13262 23100 13268 23112
rect 13223 23072 13268 23100
rect 13262 23060 13268 23072
rect 13320 23060 13326 23112
rect 15378 23100 15384 23112
rect 15339 23072 15384 23100
rect 15378 23060 15384 23072
rect 15436 23060 15442 23112
rect 15562 23060 15568 23112
rect 15620 23100 15626 23112
rect 15657 23103 15715 23109
rect 15657 23100 15669 23103
rect 15620 23072 15669 23100
rect 15620 23060 15626 23072
rect 15657 23069 15669 23072
rect 15703 23069 15715 23103
rect 15657 23063 15715 23069
rect 8478 22964 8484 22976
rect 8439 22936 8484 22964
rect 8478 22924 8484 22936
rect 8536 22924 8542 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 13078 22720 13084 22772
rect 13136 22760 13142 22772
rect 13449 22763 13507 22769
rect 13449 22760 13461 22763
rect 13136 22732 13461 22760
rect 13136 22720 13142 22732
rect 13449 22729 13461 22732
rect 13495 22729 13507 22763
rect 14734 22760 14740 22772
rect 14695 22732 14740 22760
rect 13449 22723 13507 22729
rect 14734 22720 14740 22732
rect 14792 22720 14798 22772
rect 15378 22720 15384 22772
rect 15436 22760 15442 22772
rect 15933 22763 15991 22769
rect 15933 22760 15945 22763
rect 15436 22732 15945 22760
rect 15436 22720 15442 22732
rect 15933 22729 15945 22732
rect 15979 22760 15991 22763
rect 20070 22760 20076 22772
rect 15979 22732 20076 22760
rect 15979 22729 15991 22732
rect 15933 22723 15991 22729
rect 20070 22720 20076 22732
rect 20128 22720 20134 22772
rect 12342 22584 12348 22636
rect 12400 22624 12406 22636
rect 12529 22627 12587 22633
rect 12529 22624 12541 22627
rect 12400 22596 12541 22624
rect 12400 22584 12406 22596
rect 12529 22593 12541 22596
rect 12575 22624 12587 22627
rect 13817 22627 13875 22633
rect 13817 22624 13829 22627
rect 12575 22596 13829 22624
rect 12575 22593 12587 22596
rect 12529 22587 12587 22593
rect 13817 22593 13829 22596
rect 13863 22593 13875 22627
rect 13817 22587 13875 22593
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 10689 22559 10747 22565
rect 1443 22528 2084 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 2056 22432 2084 22528
rect 10689 22525 10701 22559
rect 10735 22556 10747 22559
rect 11425 22559 11483 22565
rect 11425 22556 11437 22559
rect 10735 22528 11437 22556
rect 10735 22525 10747 22528
rect 10689 22519 10747 22525
rect 11425 22525 11437 22528
rect 11471 22556 11483 22559
rect 11885 22559 11943 22565
rect 11885 22556 11897 22559
rect 11471 22528 11897 22556
rect 11471 22525 11483 22528
rect 11425 22519 11483 22525
rect 11885 22525 11897 22528
rect 11931 22556 11943 22559
rect 12250 22556 12256 22568
rect 11931 22528 12256 22556
rect 11931 22525 11943 22528
rect 11885 22519 11943 22525
rect 12250 22516 12256 22528
rect 12308 22516 12314 22568
rect 14553 22559 14611 22565
rect 14553 22556 14565 22559
rect 14292 22528 14565 22556
rect 11517 22491 11575 22497
rect 11517 22457 11529 22491
rect 11563 22488 11575 22491
rect 12161 22491 12219 22497
rect 12161 22488 12173 22491
rect 11563 22460 12173 22488
rect 11563 22457 11575 22460
rect 11517 22451 11575 22457
rect 12161 22457 12173 22460
rect 12207 22457 12219 22491
rect 12161 22451 12219 22457
rect 12621 22491 12679 22497
rect 12621 22457 12633 22491
rect 12667 22457 12679 22491
rect 12621 22451 12679 22457
rect 13173 22491 13231 22497
rect 13173 22457 13185 22491
rect 13219 22488 13231 22491
rect 13262 22488 13268 22500
rect 13219 22460 13268 22488
rect 13219 22457 13231 22460
rect 13173 22451 13231 22457
rect 2038 22420 2044 22432
rect 1999 22392 2044 22420
rect 2038 22380 2044 22392
rect 2096 22380 2102 22432
rect 7834 22380 7840 22432
rect 7892 22420 7898 22432
rect 8478 22420 8484 22432
rect 7892 22392 8484 22420
rect 7892 22380 7898 22392
rect 8478 22380 8484 22392
rect 8536 22420 8542 22432
rect 8573 22423 8631 22429
rect 8573 22420 8585 22423
rect 8536 22392 8585 22420
rect 8536 22380 8542 22392
rect 8573 22389 8585 22392
rect 8619 22389 8631 22423
rect 12176 22420 12204 22451
rect 12636 22420 12664 22451
rect 13262 22448 13268 22460
rect 13320 22448 13326 22500
rect 12176 22392 12664 22420
rect 8573 22383 8631 22389
rect 14182 22380 14188 22432
rect 14240 22420 14246 22432
rect 14292 22429 14320 22528
rect 14553 22525 14565 22528
rect 14599 22556 14611 22559
rect 15470 22556 15476 22568
rect 14599 22528 15476 22556
rect 14599 22525 14611 22528
rect 14553 22519 14611 22525
rect 15470 22516 15476 22528
rect 15528 22516 15534 22568
rect 14277 22423 14335 22429
rect 14277 22420 14289 22423
rect 14240 22392 14289 22420
rect 14240 22380 14246 22392
rect 14277 22389 14289 22392
rect 14323 22389 14335 22423
rect 14277 22383 14335 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 12434 22108 12440 22160
rect 12492 22148 12498 22160
rect 12529 22151 12587 22157
rect 12529 22148 12541 22151
rect 12492 22120 12541 22148
rect 12492 22108 12498 22120
rect 12529 22117 12541 22120
rect 12575 22117 12587 22151
rect 12529 22111 12587 22117
rect 12437 22015 12495 22021
rect 12437 21981 12449 22015
rect 12483 22012 12495 22015
rect 12526 22012 12532 22024
rect 12483 21984 12532 22012
rect 12483 21981 12495 21984
rect 12437 21975 12495 21981
rect 12526 21972 12532 21984
rect 12584 21972 12590 22024
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 22012 12771 22015
rect 12802 22012 12808 22024
rect 12759 21984 12808 22012
rect 12759 21981 12771 21984
rect 12713 21975 12771 21981
rect 11422 21904 11428 21956
rect 11480 21944 11486 21956
rect 12728 21944 12756 21975
rect 12802 21972 12808 21984
rect 12860 21972 12866 22024
rect 11480 21916 12756 21944
rect 11480 21904 11486 21916
rect 11606 21876 11612 21888
rect 11519 21848 11612 21876
rect 11606 21836 11612 21848
rect 11664 21876 11670 21888
rect 12066 21876 12072 21888
rect 11664 21848 12072 21876
rect 11664 21836 11670 21848
rect 12066 21836 12072 21848
rect 12124 21836 12130 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 11885 21675 11943 21681
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 12526 21672 12532 21684
rect 11931 21644 12532 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 12253 21539 12311 21545
rect 12253 21505 12265 21539
rect 12299 21536 12311 21539
rect 12434 21536 12440 21548
rect 12299 21508 12440 21536
rect 12299 21505 12311 21508
rect 12253 21499 12311 21505
rect 12434 21496 12440 21508
rect 12492 21496 12498 21548
rect 12342 21428 12348 21480
rect 12400 21468 12406 21480
rect 12526 21468 12532 21480
rect 12400 21440 12532 21468
rect 12400 21428 12406 21440
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 11882 20748 11888 20800
rect 11940 20788 11946 20800
rect 12437 20791 12495 20797
rect 12437 20788 12449 20791
rect 11940 20760 12449 20788
rect 11940 20748 11946 20760
rect 12437 20757 12449 20760
rect 12483 20788 12495 20791
rect 12526 20788 12532 20800
rect 12483 20760 12532 20788
rect 12483 20757 12495 20760
rect 12437 20751 12495 20757
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 1762 20380 1768 20392
rect 1443 20352 1768 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1762 20340 1768 20352
rect 1820 20380 1826 20392
rect 1949 20383 2007 20389
rect 1949 20380 1961 20383
rect 1820 20352 1961 20380
rect 1820 20340 1826 20352
rect 1949 20349 1961 20352
rect 1995 20349 2007 20383
rect 1949 20343 2007 20349
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 15562 20040 15568 20052
rect 14332 20012 15568 20040
rect 14332 20000 14338 20012
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 25130 19496 25136 19508
rect 25091 19468 25136 19496
rect 25130 19456 25136 19468
rect 25188 19456 25194 19508
rect 1210 19252 1216 19304
rect 1268 19292 1274 19304
rect 1432 19295 1490 19301
rect 1432 19292 1444 19295
rect 1268 19264 1444 19292
rect 1268 19252 1274 19264
rect 1432 19261 1444 19264
rect 1478 19292 1490 19295
rect 1857 19295 1915 19301
rect 1857 19292 1869 19295
rect 1478 19264 1869 19292
rect 1478 19261 1490 19264
rect 1432 19255 1490 19261
rect 1857 19261 1869 19264
rect 1903 19261 1915 19295
rect 1857 19255 1915 19261
rect 24648 19295 24706 19301
rect 24648 19261 24660 19295
rect 24694 19292 24706 19295
rect 25130 19292 25136 19304
rect 24694 19264 25136 19292
rect 24694 19261 24706 19264
rect 24648 19255 24706 19261
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 1394 19116 1400 19168
rect 1452 19156 1458 19168
rect 1535 19159 1593 19165
rect 1535 19156 1547 19159
rect 1452 19128 1547 19156
rect 1452 19116 1458 19128
rect 1535 19125 1547 19128
rect 1581 19125 1593 19159
rect 1535 19119 1593 19125
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 24719 19159 24777 19165
rect 24719 19156 24731 19159
rect 22152 19128 24731 19156
rect 22152 19116 22158 19128
rect 24719 19125 24731 19128
rect 24765 19125 24777 19159
rect 24719 19119 24777 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1762 18952 1768 18964
rect 1723 18924 1768 18952
rect 1762 18912 1768 18924
rect 1820 18912 1826 18964
rect 2038 18912 2044 18964
rect 2096 18952 2102 18964
rect 2639 18955 2697 18961
rect 2639 18952 2651 18955
rect 2096 18924 2651 18952
rect 2096 18912 2102 18924
rect 2639 18921 2651 18924
rect 2685 18921 2697 18955
rect 2639 18915 2697 18921
rect 1556 18819 1614 18825
rect 1556 18785 1568 18819
rect 1602 18816 1614 18819
rect 1670 18816 1676 18828
rect 1602 18788 1676 18816
rect 1602 18785 1614 18788
rect 1556 18779 1614 18785
rect 1670 18776 1676 18788
rect 1728 18776 1734 18828
rect 2568 18819 2626 18825
rect 2568 18785 2580 18819
rect 2614 18816 2626 18819
rect 2958 18816 2964 18828
rect 2614 18788 2964 18816
rect 2614 18785 2626 18788
rect 2568 18779 2626 18785
rect 2958 18776 2964 18788
rect 3016 18776 3022 18828
rect 2041 18615 2099 18621
rect 2041 18581 2053 18615
rect 2087 18612 2099 18615
rect 2406 18612 2412 18624
rect 2087 18584 2412 18612
rect 2087 18581 2099 18584
rect 2041 18575 2099 18581
rect 2406 18572 2412 18584
rect 2464 18572 2470 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 10134 18368 10140 18420
rect 10192 18408 10198 18420
rect 10229 18411 10287 18417
rect 10229 18408 10241 18411
rect 10192 18380 10241 18408
rect 10192 18368 10198 18380
rect 10229 18377 10241 18380
rect 10275 18377 10287 18411
rect 10229 18371 10287 18377
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18173 2191 18207
rect 2406 18204 2412 18216
rect 2367 18176 2412 18204
rect 2133 18167 2191 18173
rect 1765 18139 1823 18145
rect 1765 18105 1777 18139
rect 1811 18136 1823 18139
rect 2148 18136 2176 18167
rect 2406 18164 2412 18176
rect 2464 18164 2470 18216
rect 10020 18207 10078 18213
rect 10020 18173 10032 18207
rect 10066 18204 10078 18207
rect 10134 18204 10140 18216
rect 10066 18176 10140 18204
rect 10066 18173 10078 18176
rect 10020 18167 10078 18173
rect 10134 18164 10140 18176
rect 10192 18204 10198 18216
rect 10413 18207 10471 18213
rect 10413 18204 10425 18207
rect 10192 18176 10425 18204
rect 10192 18164 10198 18176
rect 10413 18173 10425 18176
rect 10459 18173 10471 18207
rect 10413 18167 10471 18173
rect 3786 18136 3792 18148
rect 1811 18108 3792 18136
rect 1811 18105 1823 18108
rect 1765 18099 1823 18105
rect 3786 18096 3792 18108
rect 3844 18096 3850 18148
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2958 18068 2964 18080
rect 2919 18040 2964 18068
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4203 17867 4261 17873
rect 4203 17864 4215 17867
rect 4120 17836 4215 17864
rect 4120 17824 4126 17836
rect 4203 17833 4215 17836
rect 4249 17833 4261 17867
rect 7742 17864 7748 17876
rect 7703 17836 7748 17864
rect 4203 17827 4261 17833
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 9582 17756 9588 17808
rect 9640 17796 9646 17808
rect 9861 17799 9919 17805
rect 9861 17796 9873 17799
rect 9640 17768 9873 17796
rect 9640 17756 9646 17768
rect 9861 17765 9873 17768
rect 9907 17765 9919 17799
rect 9861 17759 9919 17765
rect 2130 17728 2136 17740
rect 2091 17700 2136 17728
rect 2130 17688 2136 17700
rect 2188 17688 2194 17740
rect 2406 17728 2412 17740
rect 2319 17700 2412 17728
rect 2406 17688 2412 17700
rect 2464 17728 2470 17740
rect 3694 17728 3700 17740
rect 2464 17700 3700 17728
rect 2464 17688 2470 17700
rect 3694 17688 3700 17700
rect 3752 17688 3758 17740
rect 4132 17731 4190 17737
rect 4132 17697 4144 17731
rect 4178 17728 4190 17731
rect 4614 17728 4620 17740
rect 4178 17700 4620 17728
rect 4178 17697 4190 17700
rect 4132 17691 4190 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 7374 17688 7380 17740
rect 7432 17728 7438 17740
rect 7561 17731 7619 17737
rect 7561 17728 7573 17731
rect 7432 17700 7573 17728
rect 7432 17688 7438 17700
rect 7561 17697 7573 17700
rect 7607 17697 7619 17731
rect 7561 17691 7619 17697
rect 2314 17660 2320 17672
rect 2275 17632 2320 17660
rect 2314 17620 2320 17632
rect 2372 17620 2378 17672
rect 9769 17663 9827 17669
rect 9769 17629 9781 17663
rect 9815 17629 9827 17663
rect 10134 17660 10140 17672
rect 10095 17632 10140 17660
rect 9769 17623 9827 17629
rect 9122 17552 9128 17604
rect 9180 17592 9186 17604
rect 9784 17592 9812 17623
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 11146 17592 11152 17604
rect 9180 17564 11152 17592
rect 9180 17552 9186 17564
rect 11146 17552 11152 17564
rect 11204 17552 11210 17604
rect 1670 17524 1676 17536
rect 1583 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17524 1734 17536
rect 2682 17524 2688 17536
rect 1728 17496 2688 17524
rect 1728 17484 1734 17496
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 4614 17320 4620 17332
rect 4575 17292 4620 17320
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 9122 17320 9128 17332
rect 9083 17292 9128 17320
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 7374 17212 7380 17264
rect 7432 17252 7438 17264
rect 8297 17255 8355 17261
rect 8297 17252 8309 17255
rect 7432 17224 8309 17252
rect 7432 17212 7438 17224
rect 8297 17221 8309 17224
rect 8343 17221 8355 17255
rect 8297 17215 8355 17221
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 9766 17184 9772 17196
rect 8803 17156 9772 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10134 17184 10140 17196
rect 10095 17156 10140 17184
rect 10134 17144 10140 17156
rect 10192 17144 10198 17196
rect 11146 17184 11152 17196
rect 11107 17156 11152 17184
rect 11146 17144 11152 17156
rect 11204 17144 11210 17196
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17116 2007 17119
rect 2130 17116 2136 17128
rect 1995 17088 2136 17116
rect 1995 17085 2007 17088
rect 1949 17079 2007 17085
rect 2130 17076 2136 17088
rect 2188 17116 2194 17128
rect 2501 17119 2559 17125
rect 2501 17116 2513 17119
rect 2188 17088 2513 17116
rect 2188 17076 2194 17088
rect 2501 17085 2513 17088
rect 2547 17085 2559 17119
rect 2501 17079 2559 17085
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17116 2835 17119
rect 2866 17116 2872 17128
rect 2823 17088 2872 17116
rect 2823 17085 2835 17088
rect 2777 17079 2835 17085
rect 1486 17008 1492 17060
rect 1544 17048 1550 17060
rect 2516 17048 2544 17079
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 3856 17119 3914 17125
rect 3856 17085 3868 17119
rect 3902 17116 3914 17119
rect 3970 17116 3976 17128
rect 3902 17088 3976 17116
rect 3902 17085 3914 17088
rect 3856 17079 3914 17085
rect 3970 17076 3976 17088
rect 4028 17116 4034 17128
rect 4249 17119 4307 17125
rect 4249 17116 4261 17119
rect 4028 17088 4261 17116
rect 4028 17076 4034 17088
rect 4249 17085 4261 17088
rect 4295 17085 4307 17119
rect 4249 17079 4307 17085
rect 7193 17119 7251 17125
rect 7193 17085 7205 17119
rect 7239 17116 7251 17119
rect 7650 17116 7656 17128
rect 7239 17088 7656 17116
rect 7239 17085 7251 17088
rect 7193 17079 7251 17085
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 6178 17048 6184 17060
rect 1544 17020 2176 17048
rect 2516 17020 3280 17048
rect 1544 17008 1550 17020
rect 2148 16980 2176 17020
rect 3252 16992 3280 17020
rect 4126 17020 6184 17048
rect 2317 16983 2375 16989
rect 2317 16980 2329 16983
rect 2148 16952 2329 16980
rect 2317 16949 2329 16952
rect 2363 16949 2375 16983
rect 3234 16980 3240 16992
rect 3195 16952 3240 16980
rect 2317 16943 2375 16949
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 3694 16980 3700 16992
rect 3655 16952 3700 16980
rect 3694 16940 3700 16952
rect 3752 16940 3758 16992
rect 3927 16983 3985 16989
rect 3927 16949 3939 16983
rect 3973 16980 3985 16983
rect 4126 16980 4154 17020
rect 6178 17008 6184 17020
rect 6236 17008 6242 17060
rect 9677 17051 9735 17057
rect 9677 17017 9689 17051
rect 9723 17017 9735 17051
rect 9677 17011 9735 17017
rect 7558 16980 7564 16992
rect 3973 16952 4154 16980
rect 7519 16952 7564 16980
rect 3973 16949 3985 16952
rect 3927 16943 3985 16949
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 9493 16983 9551 16989
rect 9493 16949 9505 16983
rect 9539 16980 9551 16983
rect 9582 16980 9588 16992
rect 9539 16952 9588 16980
rect 9539 16949 9551 16952
rect 9493 16943 9551 16949
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 9692 16980 9720 17011
rect 9766 17008 9772 17060
rect 9824 17048 9830 17060
rect 11330 17048 11336 17060
rect 9824 17020 11336 17048
rect 9824 17008 9830 17020
rect 11330 17008 11336 17020
rect 11388 17008 11394 17060
rect 10686 16980 10692 16992
rect 9692 16952 10692 16980
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 3694 16736 3700 16788
rect 3752 16776 3758 16788
rect 4709 16779 4767 16785
rect 4709 16776 4721 16779
rect 3752 16748 4721 16776
rect 3752 16736 3758 16748
rect 4709 16745 4721 16748
rect 4755 16745 4767 16779
rect 4709 16739 4767 16745
rect 6411 16779 6469 16785
rect 6411 16745 6423 16779
rect 6457 16776 6469 16779
rect 7374 16776 7380 16788
rect 6457 16748 7380 16776
rect 6457 16745 6469 16748
rect 6411 16739 6469 16745
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 9582 16736 9588 16788
rect 9640 16776 9646 16788
rect 9640 16748 10824 16776
rect 9640 16736 9646 16748
rect 7469 16711 7527 16717
rect 7469 16677 7481 16711
rect 7515 16708 7527 16711
rect 7558 16708 7564 16720
rect 7515 16680 7564 16708
rect 7515 16677 7527 16680
rect 7469 16671 7527 16677
rect 7558 16668 7564 16680
rect 7616 16668 7622 16720
rect 9490 16668 9496 16720
rect 9548 16708 9554 16720
rect 9861 16711 9919 16717
rect 9861 16708 9873 16711
rect 9548 16680 9873 16708
rect 9548 16668 9554 16680
rect 9861 16677 9873 16680
rect 9907 16677 9919 16711
rect 9861 16671 9919 16677
rect 10413 16711 10471 16717
rect 10413 16677 10425 16711
rect 10459 16708 10471 16711
rect 10686 16708 10692 16720
rect 10459 16680 10692 16708
rect 10459 16677 10471 16680
rect 10413 16671 10471 16677
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 10796 16708 10824 16748
rect 11241 16711 11299 16717
rect 11241 16708 11253 16711
rect 10796 16680 11253 16708
rect 11241 16677 11253 16680
rect 11287 16677 11299 16711
rect 11241 16671 11299 16677
rect 1670 16600 1676 16652
rect 1728 16640 1734 16652
rect 1857 16643 1915 16649
rect 1857 16640 1869 16643
rect 1728 16612 1869 16640
rect 1728 16600 1734 16612
rect 1857 16609 1869 16612
rect 1903 16609 1915 16643
rect 1857 16603 1915 16609
rect 3970 16600 3976 16652
rect 4028 16640 4034 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 4028 16612 4077 16640
rect 4028 16600 4034 16612
rect 4065 16609 4077 16612
rect 4111 16640 4123 16643
rect 4982 16640 4988 16652
rect 4111 16612 4988 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4982 16600 4988 16612
rect 5040 16600 5046 16652
rect 6270 16640 6276 16652
rect 6231 16612 6276 16640
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 11330 16640 11336 16652
rect 11291 16612 11336 16640
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 1762 16572 1768 16584
rect 1723 16544 1768 16572
rect 1762 16532 1768 16544
rect 1820 16532 1826 16584
rect 4433 16575 4491 16581
rect 4433 16541 4445 16575
rect 4479 16572 4491 16575
rect 5442 16572 5448 16584
rect 4479 16544 5448 16572
rect 4479 16541 4491 16544
rect 4433 16535 4491 16541
rect 5442 16532 5448 16544
rect 5500 16532 5506 16584
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 7377 16575 7435 16581
rect 7377 16572 7389 16575
rect 6696 16544 7389 16572
rect 6696 16532 6702 16544
rect 7377 16541 7389 16544
rect 7423 16572 7435 16575
rect 8202 16572 8208 16584
rect 7423 16544 8208 16572
rect 7423 16541 7435 16544
rect 7377 16535 7435 16541
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 9030 16532 9036 16584
rect 9088 16572 9094 16584
rect 9769 16575 9827 16581
rect 9769 16572 9781 16575
rect 9088 16544 9781 16572
rect 9088 16532 9094 16544
rect 9769 16541 9781 16544
rect 9815 16541 9827 16575
rect 9769 16535 9827 16541
rect 7926 16504 7932 16516
rect 7887 16476 7932 16504
rect 7926 16464 7932 16476
rect 7984 16464 7990 16516
rect 2866 16436 2872 16448
rect 2827 16408 2872 16436
rect 2866 16396 2872 16408
rect 2924 16396 2930 16448
rect 3878 16396 3884 16448
rect 3936 16436 3942 16448
rect 4203 16439 4261 16445
rect 4203 16436 4215 16439
rect 3936 16408 4215 16436
rect 3936 16396 3942 16408
rect 4203 16405 4215 16408
rect 4249 16405 4261 16439
rect 4338 16436 4344 16448
rect 4299 16408 4344 16436
rect 4203 16399 4261 16405
rect 4338 16396 4344 16408
rect 4396 16396 4402 16448
rect 5074 16436 5080 16448
rect 5035 16408 5080 16436
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1673 16235 1731 16241
rect 1673 16201 1685 16235
rect 1719 16232 1731 16235
rect 1762 16232 1768 16244
rect 1719 16204 1768 16232
rect 1719 16201 1731 16204
rect 1673 16195 1731 16201
rect 1762 16192 1768 16204
rect 1820 16192 1826 16244
rect 3142 16232 3148 16244
rect 3103 16204 3148 16232
rect 3142 16192 3148 16204
rect 3200 16192 3206 16244
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5813 16235 5871 16241
rect 5813 16232 5825 16235
rect 5040 16204 5825 16232
rect 5040 16192 5046 16204
rect 5813 16201 5825 16204
rect 5859 16201 5871 16235
rect 6638 16232 6644 16244
rect 6599 16204 6644 16232
rect 5813 16195 5871 16201
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 7285 16235 7343 16241
rect 7285 16201 7297 16235
rect 7331 16232 7343 16235
rect 7558 16232 7564 16244
rect 7331 16204 7564 16232
rect 7331 16201 7343 16204
rect 7285 16195 7343 16201
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 11609 16235 11667 16241
rect 11609 16232 11621 16235
rect 11388 16204 11621 16232
rect 11388 16192 11394 16204
rect 11609 16201 11621 16204
rect 11655 16201 11667 16235
rect 11609 16195 11667 16201
rect 3467 16167 3525 16173
rect 3467 16133 3479 16167
rect 3513 16164 3525 16167
rect 9030 16164 9036 16176
rect 3513 16136 9036 16164
rect 3513 16133 3525 16136
rect 3467 16127 3525 16133
rect 9030 16124 9036 16136
rect 9088 16164 9094 16176
rect 10965 16167 11023 16173
rect 10965 16164 10977 16167
rect 9088 16136 10977 16164
rect 9088 16124 9094 16136
rect 10965 16133 10977 16136
rect 11011 16133 11023 16167
rect 10965 16127 11023 16133
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 6270 16096 6276 16108
rect 1903 16068 2912 16096
rect 6183 16068 6276 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 1949 15963 2007 15969
rect 1949 15929 1961 15963
rect 1995 15929 2007 15963
rect 1949 15923 2007 15929
rect 2501 15963 2559 15969
rect 2501 15929 2513 15963
rect 2547 15960 2559 15963
rect 2682 15960 2688 15972
rect 2547 15932 2688 15960
rect 2547 15929 2559 15932
rect 2501 15923 2559 15929
rect 1762 15852 1768 15904
rect 1820 15892 1826 15904
rect 1964 15892 1992 15923
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 2884 15901 2912 16068
rect 6270 16056 6276 16068
rect 6328 16096 6334 16108
rect 7926 16096 7932 16108
rect 6328 16068 7932 16096
rect 6328 16056 6334 16068
rect 7926 16056 7932 16068
rect 7984 16056 7990 16108
rect 9125 16099 9183 16105
rect 9125 16065 9137 16099
rect 9171 16096 9183 16099
rect 9766 16096 9772 16108
rect 9171 16068 9772 16096
rect 9171 16065 9183 16068
rect 9125 16059 9183 16065
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16096 10379 16099
rect 10686 16096 10692 16108
rect 10367 16068 10692 16096
rect 10367 16065 10379 16068
rect 10321 16059 10379 16065
rect 10686 16056 10692 16068
rect 10744 16056 10750 16108
rect 3142 15988 3148 16040
rect 3200 16028 3206 16040
rect 3364 16031 3422 16037
rect 3364 16028 3376 16031
rect 3200 16000 3376 16028
rect 3200 15988 3206 16000
rect 3364 15997 3376 16000
rect 3410 15997 3422 16031
rect 5074 16028 5080 16040
rect 5035 16000 5080 16028
rect 3364 15991 3422 15997
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 4430 15960 4436 15972
rect 4391 15932 4436 15960
rect 4430 15920 4436 15932
rect 4488 15920 4494 15972
rect 7466 15960 7472 15972
rect 7427 15932 7472 15960
rect 7466 15920 7472 15932
rect 7524 15920 7530 15972
rect 7561 15963 7619 15969
rect 7561 15929 7573 15963
rect 7607 15960 7619 15963
rect 7650 15960 7656 15972
rect 7607 15932 7656 15960
rect 7607 15929 7619 15932
rect 7561 15923 7619 15929
rect 7650 15920 7656 15932
rect 7708 15960 7714 15972
rect 8389 15963 8447 15969
rect 8389 15960 8401 15963
rect 7708 15932 8401 15960
rect 7708 15920 7714 15932
rect 8389 15929 8401 15932
rect 8435 15929 8447 15963
rect 8389 15923 8447 15929
rect 9677 15963 9735 15969
rect 9677 15929 9689 15963
rect 9723 15929 9735 15963
rect 9677 15923 9735 15929
rect 1820 15864 1992 15892
rect 2869 15895 2927 15901
rect 1820 15852 1826 15864
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 3050 15892 3056 15904
rect 2915 15864 3056 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 4157 15895 4215 15901
rect 4157 15861 4169 15895
rect 4203 15892 4215 15895
rect 4338 15892 4344 15904
rect 4203 15864 4344 15892
rect 4203 15861 4215 15864
rect 4157 15855 4215 15861
rect 4338 15852 4344 15864
rect 4396 15892 4402 15904
rect 5258 15892 5264 15904
rect 4396 15864 5264 15892
rect 4396 15852 4402 15864
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 5442 15892 5448 15904
rect 5403 15864 5448 15892
rect 5442 15852 5448 15864
rect 5500 15852 5506 15904
rect 9490 15892 9496 15904
rect 9451 15864 9496 15892
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 9692 15892 9720 15923
rect 9766 15920 9772 15972
rect 9824 15960 9830 15972
rect 9824 15932 9869 15960
rect 9824 15920 9830 15932
rect 10686 15892 10692 15904
rect 9692 15864 10692 15892
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 11146 15892 11152 15904
rect 11107 15864 11152 15892
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 8202 15688 8208 15700
rect 8163 15660 8208 15688
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 1854 15580 1860 15632
rect 1912 15620 1918 15632
rect 1949 15623 2007 15629
rect 1949 15620 1961 15623
rect 1912 15592 1961 15620
rect 1912 15580 1918 15592
rect 1949 15589 1961 15592
rect 1995 15589 2007 15623
rect 6822 15620 6828 15632
rect 6783 15592 6828 15620
rect 1949 15583 2007 15589
rect 6822 15580 6828 15592
rect 6880 15580 6886 15632
rect 7377 15623 7435 15629
rect 7377 15589 7389 15623
rect 7423 15620 7435 15623
rect 7466 15620 7472 15632
rect 7423 15592 7472 15620
rect 7423 15589 7435 15592
rect 7377 15583 7435 15589
rect 7466 15580 7472 15592
rect 7524 15620 7530 15632
rect 8021 15623 8079 15629
rect 8021 15620 8033 15623
rect 7524 15592 8033 15620
rect 7524 15580 7530 15592
rect 8021 15589 8033 15592
rect 8067 15589 8079 15623
rect 8021 15583 8079 15589
rect 9490 15580 9496 15632
rect 9548 15620 9554 15632
rect 9677 15623 9735 15629
rect 9677 15620 9689 15623
rect 9548 15592 9689 15620
rect 9548 15580 9554 15592
rect 9677 15589 9689 15592
rect 9723 15589 9735 15623
rect 9677 15583 9735 15589
rect 4982 15552 4988 15564
rect 4943 15524 4988 15552
rect 4982 15512 4988 15524
rect 5040 15512 5046 15564
rect 9766 15552 9772 15564
rect 9727 15524 9772 15552
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 11606 15552 11612 15564
rect 11567 15524 11612 15552
rect 11606 15512 11612 15524
rect 11664 15512 11670 15564
rect 1302 15444 1308 15496
rect 1360 15484 1366 15496
rect 1857 15487 1915 15493
rect 1857 15484 1869 15487
rect 1360 15456 1869 15484
rect 1360 15444 1366 15456
rect 1857 15453 1869 15456
rect 1903 15484 1915 15487
rect 3142 15484 3148 15496
rect 1903 15456 3148 15484
rect 1903 15453 1915 15456
rect 1857 15447 1915 15453
rect 3142 15444 3148 15456
rect 3200 15444 3206 15496
rect 6178 15444 6184 15496
rect 6236 15484 6242 15496
rect 6733 15487 6791 15493
rect 6733 15484 6745 15487
rect 6236 15456 6745 15484
rect 6236 15444 6242 15456
rect 6733 15453 6745 15456
rect 6779 15453 6791 15487
rect 6733 15447 6791 15453
rect 10778 15444 10784 15496
rect 10836 15484 10842 15496
rect 11241 15487 11299 15493
rect 11241 15484 11253 15487
rect 10836 15456 11253 15484
rect 10836 15444 10842 15456
rect 11241 15453 11253 15456
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 2409 15419 2467 15425
rect 2409 15385 2421 15419
rect 2455 15385 2467 15419
rect 2409 15379 2467 15385
rect 2424 15348 2452 15379
rect 2869 15351 2927 15357
rect 2869 15348 2881 15351
rect 2424 15320 2881 15348
rect 2869 15317 2881 15320
rect 2915 15348 2927 15351
rect 2958 15348 2964 15360
rect 2915 15320 2964 15348
rect 2915 15317 2927 15320
rect 2869 15311 2927 15317
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 3878 15348 3884 15360
rect 3839 15320 3884 15348
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 4614 15348 4620 15360
rect 4575 15320 4620 15348
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 7742 15348 7748 15360
rect 7703 15320 7748 15348
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 3142 15144 3148 15156
rect 3103 15116 3148 15144
rect 3142 15104 3148 15116
rect 3200 15104 3206 15156
rect 3602 15144 3608 15156
rect 3563 15116 3608 15144
rect 3602 15104 3608 15116
rect 3660 15104 3666 15156
rect 4065 15147 4123 15153
rect 4065 15113 4077 15147
rect 4111 15144 4123 15147
rect 4430 15144 4436 15156
rect 4111 15116 4436 15144
rect 4111 15113 4123 15116
rect 4065 15107 4123 15113
rect 4430 15104 4436 15116
rect 4488 15104 4494 15156
rect 4982 15104 4988 15156
rect 5040 15144 5046 15156
rect 5169 15147 5227 15153
rect 5169 15144 5181 15147
rect 5040 15116 5181 15144
rect 5040 15104 5046 15116
rect 5169 15113 5181 15116
rect 5215 15113 5227 15147
rect 6178 15144 6184 15156
rect 6139 15116 6184 15144
rect 5169 15107 5227 15113
rect 6178 15104 6184 15116
rect 6236 15104 6242 15156
rect 11606 15144 11612 15156
rect 11567 15116 11612 15144
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 25130 15144 25136 15156
rect 25091 15116 25136 15144
rect 25130 15104 25136 15116
rect 25188 15104 25194 15156
rect 2682 15076 2688 15088
rect 2643 15048 2688 15076
rect 2682 15036 2688 15048
rect 2740 15036 2746 15088
rect 3050 15036 3056 15088
rect 3108 15076 3114 15088
rect 3108 15048 5764 15076
rect 3108 15036 3114 15048
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 15008 2191 15011
rect 2958 15008 2964 15020
rect 2179 14980 2964 15008
rect 2179 14977 2191 14980
rect 2133 14971 2191 14977
rect 2958 14968 2964 14980
rect 3016 14968 3022 15020
rect 3602 14968 3608 15020
rect 3660 15008 3666 15020
rect 4249 15011 4307 15017
rect 4249 15008 4261 15011
rect 3660 14980 4261 15008
rect 3660 14968 3666 14980
rect 4249 14977 4261 14980
rect 4295 14977 4307 15011
rect 4706 15008 4712 15020
rect 4667 14980 4712 15008
rect 4249 14971 4307 14977
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 5736 15017 5764 15048
rect 6822 15036 6828 15088
rect 6880 15076 6886 15088
rect 7101 15079 7159 15085
rect 7101 15076 7113 15079
rect 6880 15048 7113 15076
rect 6880 15036 6886 15048
rect 7101 15045 7113 15048
rect 7147 15076 7159 15079
rect 11238 15076 11244 15088
rect 7147 15048 8892 15076
rect 11199 15048 11244 15076
rect 7147 15045 7159 15048
rect 7101 15039 7159 15045
rect 5721 15011 5779 15017
rect 5721 14977 5733 15011
rect 5767 14977 5779 15011
rect 5721 14971 5779 14977
rect 7466 14968 7472 15020
rect 7524 15008 7530 15020
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 7524 14980 7757 15008
rect 7524 14968 7530 14980
rect 7745 14977 7757 14980
rect 7791 14977 7803 15011
rect 8864 15008 8892 15048
rect 11238 15036 11244 15048
rect 11296 15036 11302 15088
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8864 14980 8953 15008
rect 7745 14971 7803 14977
rect 8941 14977 8953 14980
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 15008 10195 15011
rect 10689 15011 10747 15017
rect 10689 15008 10701 15011
rect 10183 14980 10701 15008
rect 10183 14977 10195 14980
rect 10137 14971 10195 14977
rect 10689 14977 10701 14980
rect 10735 15008 10747 15011
rect 11146 15008 11152 15020
rect 10735 14980 11152 15008
rect 10735 14977 10747 14980
rect 10689 14971 10747 14977
rect 11146 14968 11152 14980
rect 11204 14968 11210 15020
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14940 8907 14943
rect 9033 14943 9091 14949
rect 9033 14940 9045 14943
rect 8895 14912 9045 14940
rect 8895 14909 8907 14912
rect 8849 14903 8907 14909
rect 9033 14909 9045 14912
rect 9079 14909 9091 14943
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 9033 14903 9091 14909
rect 12176 14912 12449 14940
rect 1670 14832 1676 14884
rect 1728 14872 1734 14884
rect 2222 14872 2228 14884
rect 1728 14844 2228 14872
rect 1728 14832 1734 14844
rect 2222 14832 2228 14844
rect 2280 14832 2286 14884
rect 4341 14875 4399 14881
rect 4341 14841 4353 14875
rect 4387 14872 4399 14875
rect 4430 14872 4436 14884
rect 4387 14844 4436 14872
rect 4387 14841 4399 14844
rect 4341 14835 4399 14841
rect 4430 14832 4436 14844
rect 4488 14832 4494 14884
rect 7469 14875 7527 14881
rect 7469 14841 7481 14875
rect 7515 14841 7527 14875
rect 7469 14835 7527 14841
rect 7561 14875 7619 14881
rect 7561 14841 7573 14875
rect 7607 14872 7619 14875
rect 7742 14872 7748 14884
rect 7607 14844 7748 14872
rect 7607 14841 7619 14844
rect 7561 14835 7619 14841
rect 1854 14804 1860 14816
rect 1815 14776 1860 14804
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 6641 14807 6699 14813
rect 6641 14773 6653 14807
rect 6687 14804 6699 14807
rect 7484 14804 7512 14835
rect 7742 14832 7748 14844
rect 7800 14872 7806 14884
rect 8864 14872 8892 14903
rect 7800 14844 8892 14872
rect 7800 14832 7806 14844
rect 10778 14832 10784 14884
rect 10836 14872 10842 14884
rect 10836 14844 10881 14872
rect 10836 14832 10842 14844
rect 8202 14804 8208 14816
rect 6687 14776 8208 14804
rect 6687 14773 6699 14776
rect 6641 14767 6699 14773
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 10505 14807 10563 14813
rect 10505 14773 10517 14807
rect 10551 14804 10563 14807
rect 10796 14804 10824 14832
rect 12176 14816 12204 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 24648 14943 24706 14949
rect 24648 14909 24660 14943
rect 24694 14940 24706 14943
rect 25130 14940 25136 14952
rect 24694 14912 25136 14940
rect 24694 14909 24706 14912
rect 24648 14903 24706 14909
rect 12250 14832 12256 14884
rect 12308 14872 12314 14884
rect 12912 14872 12940 14903
rect 25130 14900 25136 14912
rect 25188 14900 25194 14952
rect 12308 14844 12940 14872
rect 12308 14832 12314 14844
rect 12158 14804 12164 14816
rect 10551 14776 10824 14804
rect 12119 14776 12164 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 12158 14764 12164 14776
rect 12216 14764 12222 14816
rect 12526 14804 12532 14816
rect 12487 14776 12532 14804
rect 12526 14764 12532 14776
rect 12584 14764 12590 14816
rect 24719 14807 24777 14813
rect 24719 14773 24731 14807
rect 24765 14804 24777 14807
rect 25130 14804 25136 14816
rect 24765 14776 25136 14804
rect 24765 14773 24777 14776
rect 24719 14767 24777 14773
rect 25130 14764 25136 14776
rect 25188 14764 25194 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 7101 14603 7159 14609
rect 7101 14600 7113 14603
rect 7064 14572 7113 14600
rect 7064 14560 7070 14572
rect 7101 14569 7113 14572
rect 7147 14569 7159 14603
rect 7650 14600 7656 14612
rect 7611 14572 7656 14600
rect 7101 14563 7159 14569
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 9493 14603 9551 14609
rect 9493 14569 9505 14603
rect 9539 14600 9551 14603
rect 9766 14600 9772 14612
rect 9539 14572 9772 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10045 14603 10103 14609
rect 10045 14600 10057 14603
rect 9916 14572 10057 14600
rect 9916 14560 9922 14572
rect 10045 14569 10057 14572
rect 10091 14569 10103 14603
rect 10045 14563 10103 14569
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 11330 14600 11336 14612
rect 10643 14572 11336 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 13078 14600 13084 14612
rect 13039 14572 13084 14600
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 2593 14535 2651 14541
rect 2593 14501 2605 14535
rect 2639 14532 2651 14535
rect 2774 14532 2780 14544
rect 2639 14504 2780 14532
rect 2639 14501 2651 14504
rect 2593 14495 2651 14501
rect 2774 14492 2780 14504
rect 2832 14492 2838 14544
rect 4525 14535 4583 14541
rect 4525 14501 4537 14535
rect 4571 14532 4583 14535
rect 4614 14532 4620 14544
rect 4571 14504 4620 14532
rect 4571 14501 4583 14504
rect 4525 14495 4583 14501
rect 4614 14492 4620 14504
rect 4672 14492 4678 14544
rect 11606 14532 11612 14544
rect 11567 14504 11612 14532
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 23842 14492 23848 14544
rect 23900 14532 23906 14544
rect 24213 14535 24271 14541
rect 24213 14532 24225 14535
rect 23900 14504 24225 14532
rect 23900 14492 23906 14504
rect 24213 14501 24225 14504
rect 24259 14501 24271 14535
rect 24213 14495 24271 14501
rect 1464 14467 1522 14473
rect 1464 14433 1476 14467
rect 1510 14464 1522 14467
rect 1578 14464 1584 14476
rect 1510 14436 1584 14464
rect 1510 14433 1522 14436
rect 1464 14427 1522 14433
rect 1578 14424 1584 14436
rect 1636 14424 1642 14476
rect 12986 14464 12992 14476
rect 12947 14436 12992 14464
rect 12986 14424 12992 14436
rect 13044 14424 13050 14476
rect 13449 14467 13507 14473
rect 13449 14433 13461 14467
rect 13495 14464 13507 14467
rect 14458 14464 14464 14476
rect 13495 14436 14464 14464
rect 13495 14433 13507 14436
rect 13449 14427 13507 14433
rect 2498 14396 2504 14408
rect 2459 14368 2504 14396
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 2958 14396 2964 14408
rect 2919 14368 2964 14396
rect 2958 14356 2964 14368
rect 3016 14356 3022 14408
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 4433 14399 4491 14405
rect 4433 14396 4445 14399
rect 4120 14368 4445 14396
rect 4120 14356 4126 14368
rect 4433 14365 4445 14368
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 4522 14356 4528 14408
rect 4580 14396 4586 14408
rect 4709 14399 4767 14405
rect 4709 14396 4721 14399
rect 4580 14368 4721 14396
rect 4580 14356 4586 14368
rect 4709 14365 4721 14368
rect 4755 14365 4767 14399
rect 4709 14359 4767 14365
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14396 6791 14399
rect 8018 14396 8024 14408
rect 6779 14368 8024 14396
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 9490 14356 9496 14408
rect 9548 14396 9554 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 9548 14368 9689 14396
rect 9548 14356 9554 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14396 11391 14399
rect 11514 14396 11520 14408
rect 11379 14368 11520 14396
rect 11379 14365 11391 14368
rect 11333 14359 11391 14365
rect 11514 14356 11520 14368
rect 11572 14356 11578 14408
rect 11793 14399 11851 14405
rect 11793 14365 11805 14399
rect 11839 14365 11851 14399
rect 13464 14396 13492 14427
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 11793 14359 11851 14365
rect 12452 14368 13492 14396
rect 24121 14399 24179 14405
rect 11238 14288 11244 14340
rect 11296 14328 11302 14340
rect 11808 14328 11836 14359
rect 11296 14300 11836 14328
rect 11296 14288 11302 14300
rect 1535 14263 1593 14269
rect 1535 14229 1547 14263
rect 1581 14260 1593 14263
rect 1762 14260 1768 14272
rect 1581 14232 1768 14260
rect 1581 14229 1593 14232
rect 1535 14223 1593 14229
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 1949 14263 2007 14269
rect 1949 14229 1961 14263
rect 1995 14260 2007 14263
rect 2038 14260 2044 14272
rect 1995 14232 2044 14260
rect 1995 14229 2007 14232
rect 1949 14223 2007 14229
rect 2038 14220 2044 14232
rect 2096 14220 2102 14272
rect 4706 14220 4712 14272
rect 4764 14260 4770 14272
rect 5445 14263 5503 14269
rect 5445 14260 5457 14263
rect 4764 14232 5457 14260
rect 4764 14220 4770 14232
rect 5445 14229 5457 14232
rect 5491 14260 5503 14263
rect 6362 14260 6368 14272
rect 5491 14232 6368 14260
rect 5491 14229 5503 14232
rect 5445 14223 5503 14229
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 8938 14260 8944 14272
rect 8899 14232 8944 14260
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 12250 14220 12256 14272
rect 12308 14260 12314 14272
rect 12452 14269 12480 14368
rect 24121 14365 24133 14399
rect 24167 14365 24179 14399
rect 24121 14359 24179 14365
rect 24765 14399 24823 14405
rect 24765 14365 24777 14399
rect 24811 14396 24823 14399
rect 24854 14396 24860 14408
rect 24811 14368 24860 14396
rect 24811 14365 24823 14368
rect 24765 14359 24823 14365
rect 24136 14328 24164 14359
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 25130 14328 25136 14340
rect 24136 14300 25136 14328
rect 25130 14288 25136 14300
rect 25188 14288 25194 14340
rect 12437 14263 12495 14269
rect 12437 14260 12449 14263
rect 12308 14232 12449 14260
rect 12308 14220 12314 14232
rect 12437 14229 12449 14232
rect 12483 14229 12495 14263
rect 12437 14223 12495 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 2222 14016 2228 14068
rect 2280 14056 2286 14068
rect 2685 14059 2743 14065
rect 2685 14056 2697 14059
rect 2280 14028 2697 14056
rect 2280 14016 2286 14028
rect 2685 14025 2697 14028
rect 2731 14025 2743 14059
rect 4062 14056 4068 14068
rect 2685 14019 2743 14025
rect 3528 14028 4068 14056
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 2314 13920 2320 13932
rect 1811 13892 2320 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 2314 13880 2320 13892
rect 2372 13920 2378 13932
rect 3528 13929 3556 14028
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 4433 14059 4491 14065
rect 4433 14025 4445 14059
rect 4479 14056 4491 14059
rect 4614 14056 4620 14068
rect 4479 14028 4620 14056
rect 4479 14025 4491 14028
rect 4433 14019 4491 14025
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 7742 14056 7748 14068
rect 7703 14028 7748 14056
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8018 14056 8024 14068
rect 7979 14028 8024 14056
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 9766 14056 9772 14068
rect 9727 14028 9772 14056
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 11606 14056 11612 14068
rect 11563 14028 11612 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 11606 14016 11612 14028
rect 11664 14056 11670 14068
rect 11793 14059 11851 14065
rect 11793 14056 11805 14059
rect 11664 14028 11805 14056
rect 11664 14016 11670 14028
rect 11793 14025 11805 14028
rect 11839 14025 11851 14059
rect 12250 14056 12256 14068
rect 12211 14028 12256 14056
rect 11793 14019 11851 14025
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 12805 14059 12863 14065
rect 12805 14025 12817 14059
rect 12851 14056 12863 14059
rect 12986 14056 12992 14068
rect 12851 14028 12992 14056
rect 12851 14025 12863 14028
rect 12805 14019 12863 14025
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 14182 14056 14188 14068
rect 14143 14028 14188 14056
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 25130 14056 25136 14068
rect 25091 14028 25136 14056
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 4522 13948 4528 14000
rect 4580 13988 4586 14000
rect 4580 13960 4936 13988
rect 4580 13948 4586 13960
rect 3329 13923 3387 13929
rect 3329 13920 3341 13923
rect 2372 13892 3341 13920
rect 2372 13880 2378 13892
rect 3329 13889 3341 13892
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13920 4675 13923
rect 4706 13920 4712 13932
rect 4663 13892 4712 13920
rect 4663 13889 4675 13892
rect 4617 13883 4675 13889
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 4908 13929 4936 13960
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13920 6883 13923
rect 7098 13920 7104 13932
rect 6871 13892 7104 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 8849 13923 8907 13929
rect 8849 13889 8861 13923
rect 8895 13920 8907 13923
rect 8938 13920 8944 13932
rect 8895 13892 8944 13920
rect 8895 13889 8907 13892
rect 8849 13883 8907 13889
rect 8938 13880 8944 13892
rect 8996 13920 9002 13932
rect 10597 13923 10655 13929
rect 8996 13892 9628 13920
rect 8996 13880 9002 13892
rect 4709 13787 4767 13793
rect 4709 13753 4721 13787
rect 4755 13784 4767 13787
rect 4890 13784 4896 13796
rect 4755 13756 4896 13784
rect 4755 13753 4767 13756
rect 4709 13747 4767 13753
rect 4890 13744 4896 13756
rect 4948 13784 4954 13796
rect 5537 13787 5595 13793
rect 5537 13784 5549 13787
rect 4948 13756 5549 13784
rect 4948 13744 4954 13756
rect 5537 13753 5549 13756
rect 5583 13753 5595 13787
rect 5537 13747 5595 13753
rect 7146 13787 7204 13793
rect 7146 13753 7158 13787
rect 7192 13753 7204 13787
rect 7146 13747 7204 13753
rect 9170 13787 9228 13793
rect 9170 13753 9182 13787
rect 9216 13753 9228 13787
rect 9600 13784 9628 13892
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 10778 13920 10784 13932
rect 10643 13892 10784 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 10778 13880 10784 13892
rect 10836 13920 10842 13932
rect 13078 13920 13084 13932
rect 10836 13892 13084 13920
rect 10836 13880 10842 13892
rect 13078 13880 13084 13892
rect 13136 13880 13142 13932
rect 14461 13923 14519 13929
rect 14461 13920 14473 13923
rect 13786 13892 14473 13920
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13852 13323 13855
rect 13354 13852 13360 13864
rect 13311 13824 13360 13852
rect 13311 13821 13323 13824
rect 13265 13815 13323 13821
rect 13354 13812 13360 13824
rect 13412 13852 13418 13864
rect 13786 13852 13814 13892
rect 14461 13889 14473 13892
rect 14507 13889 14519 13923
rect 14461 13883 14519 13889
rect 24213 13923 24271 13929
rect 24213 13889 24225 13923
rect 24259 13920 24271 13923
rect 24670 13920 24676 13932
rect 24259 13892 24676 13920
rect 24259 13889 24271 13892
rect 24213 13883 24271 13889
rect 24670 13880 24676 13892
rect 24728 13880 24734 13932
rect 13412 13824 13814 13852
rect 13412 13812 13418 13824
rect 9766 13784 9772 13796
rect 9600 13756 9772 13784
rect 9170 13747 9228 13753
rect 2038 13676 2044 13728
rect 2096 13716 2102 13728
rect 2133 13719 2191 13725
rect 2133 13716 2145 13719
rect 2096 13688 2145 13716
rect 2096 13676 2102 13688
rect 2133 13685 2145 13688
rect 2179 13685 2191 13719
rect 2133 13679 2191 13685
rect 2774 13676 2780 13728
rect 2832 13716 2838 13728
rect 2961 13719 3019 13725
rect 2961 13716 2973 13719
rect 2832 13688 2973 13716
rect 2832 13676 2838 13688
rect 2961 13685 2973 13688
rect 3007 13685 3019 13719
rect 2961 13679 3019 13685
rect 6273 13719 6331 13725
rect 6273 13685 6285 13719
rect 6319 13716 6331 13719
rect 6638 13716 6644 13728
rect 6319 13688 6644 13716
rect 6319 13685 6331 13688
rect 6273 13679 6331 13685
rect 6638 13676 6644 13688
rect 6696 13716 6702 13728
rect 7006 13716 7012 13728
rect 6696 13688 7012 13716
rect 6696 13676 6702 13688
rect 7006 13676 7012 13688
rect 7064 13716 7070 13728
rect 7161 13716 7189 13747
rect 8665 13719 8723 13725
rect 8665 13716 8677 13719
rect 7064 13688 8677 13716
rect 7064 13676 7070 13688
rect 8665 13685 8677 13688
rect 8711 13716 8723 13719
rect 9185 13716 9213 13747
rect 9766 13744 9772 13756
rect 9824 13744 9830 13796
rect 10918 13787 10976 13793
rect 10918 13784 10930 13787
rect 10428 13756 10930 13784
rect 9858 13716 9864 13728
rect 8711 13688 9864 13716
rect 8711 13685 8723 13688
rect 8665 13679 8723 13685
rect 9858 13676 9864 13688
rect 9916 13716 9922 13728
rect 10428 13725 10456 13756
rect 10918 13753 10930 13756
rect 10964 13753 10976 13787
rect 13586 13787 13644 13793
rect 13586 13784 13598 13787
rect 10918 13747 10976 13753
rect 13188 13756 13598 13784
rect 13188 13728 13216 13756
rect 13586 13753 13598 13756
rect 13632 13753 13644 13787
rect 13586 13747 13644 13753
rect 24305 13787 24363 13793
rect 24305 13753 24317 13787
rect 24351 13753 24363 13787
rect 24854 13784 24860 13796
rect 24815 13756 24860 13784
rect 24305 13747 24363 13753
rect 10045 13719 10103 13725
rect 10045 13716 10057 13719
rect 9916 13688 10057 13716
rect 9916 13676 9922 13688
rect 10045 13685 10057 13688
rect 10091 13716 10103 13719
rect 10413 13719 10471 13725
rect 10413 13716 10425 13719
rect 10091 13688 10425 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 10413 13685 10425 13688
rect 10459 13685 10471 13719
rect 13170 13716 13176 13728
rect 13131 13688 13176 13716
rect 10413 13679 10471 13685
rect 13170 13676 13176 13688
rect 13228 13676 13234 13728
rect 23477 13719 23535 13725
rect 23477 13685 23489 13719
rect 23523 13716 23535 13719
rect 23842 13716 23848 13728
rect 23523 13688 23848 13716
rect 23523 13685 23535 13688
rect 23477 13679 23535 13685
rect 23842 13676 23848 13688
rect 23900 13676 23906 13728
rect 24026 13716 24032 13728
rect 23987 13688 24032 13716
rect 24026 13676 24032 13688
rect 24084 13716 24090 13728
rect 24320 13716 24348 13747
rect 24854 13744 24860 13756
rect 24912 13744 24918 13796
rect 24084 13688 24348 13716
rect 24084 13676 24090 13688
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 4614 13512 4620 13524
rect 4575 13484 4620 13512
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 4890 13472 4896 13524
rect 4948 13512 4954 13524
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 4948 13484 5181 13512
rect 4948 13472 4954 13484
rect 5169 13481 5181 13484
rect 5215 13481 5227 13515
rect 5169 13475 5227 13481
rect 7837 13515 7895 13521
rect 7837 13481 7849 13515
rect 7883 13512 7895 13515
rect 8018 13512 8024 13524
rect 7883 13484 8024 13512
rect 7883 13481 7895 13484
rect 7837 13475 7895 13481
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 9766 13512 9772 13524
rect 9727 13484 9772 13512
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 10778 13512 10784 13524
rect 10739 13484 10784 13512
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12250 13512 12256 13524
rect 12211 13484 12256 13512
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 13354 13512 13360 13524
rect 13315 13484 13360 13512
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 24026 13512 24032 13524
rect 23987 13484 24032 13512
rect 24026 13472 24032 13484
rect 24084 13472 24090 13524
rect 2038 13404 2044 13456
rect 2096 13444 2102 13456
rect 2178 13447 2236 13453
rect 2178 13444 2190 13447
rect 2096 13416 2190 13444
rect 2096 13404 2102 13416
rect 2178 13413 2190 13416
rect 2224 13413 2236 13447
rect 2178 13407 2236 13413
rect 5074 13404 5080 13456
rect 5132 13444 5138 13456
rect 6181 13447 6239 13453
rect 6181 13444 6193 13447
rect 5132 13416 6193 13444
rect 5132 13404 5138 13416
rect 6181 13413 6193 13416
rect 6227 13413 6239 13447
rect 6181 13407 6239 13413
rect 7742 13376 7748 13388
rect 7703 13348 7748 13376
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 8021 13379 8079 13385
rect 8021 13345 8033 13379
rect 8067 13345 8079 13379
rect 9674 13376 9680 13388
rect 9635 13348 9680 13376
rect 8021 13339 8079 13345
rect 1857 13311 1915 13317
rect 1857 13277 1869 13311
rect 1903 13308 1915 13311
rect 1946 13308 1952 13320
rect 1903 13280 1952 13308
rect 1903 13277 1915 13280
rect 1857 13271 1915 13277
rect 1946 13268 1952 13280
rect 2004 13308 2010 13320
rect 2590 13308 2596 13320
rect 2004 13280 2596 13308
rect 2004 13268 2010 13280
rect 2590 13268 2596 13280
rect 2648 13268 2654 13320
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13308 3939 13311
rect 4249 13311 4307 13317
rect 4249 13308 4261 13311
rect 3927 13280 4261 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 4249 13277 4261 13280
rect 4295 13308 4307 13311
rect 4338 13308 4344 13320
rect 4295 13280 4344 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13308 5963 13311
rect 6089 13311 6147 13317
rect 6089 13308 6101 13311
rect 5951 13280 6101 13308
rect 5951 13277 5963 13280
rect 5905 13271 5963 13277
rect 6089 13277 6101 13280
rect 6135 13308 6147 13311
rect 6178 13308 6184 13320
rect 6135 13280 6184 13308
rect 6135 13277 6147 13280
rect 6089 13271 6147 13277
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 6362 13308 6368 13320
rect 6323 13280 6368 13308
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 7432 13280 7481 13308
rect 7432 13268 7438 13280
rect 7469 13277 7481 13280
rect 7515 13308 7527 13311
rect 8036 13308 8064 13339
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 9876 13348 10149 13376
rect 7515 13280 8064 13308
rect 8665 13311 8723 13317
rect 7515 13277 7527 13280
rect 7469 13271 7527 13277
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 8938 13308 8944 13320
rect 8711 13280 8944 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 8938 13268 8944 13280
rect 8996 13308 9002 13320
rect 9876 13308 9904 13348
rect 10137 13345 10149 13348
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 12216 13348 13093 13376
rect 12216 13336 12222 13348
rect 13081 13345 13093 13348
rect 13127 13345 13139 13379
rect 13538 13376 13544 13388
rect 13499 13348 13544 13376
rect 13081 13339 13139 13345
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 23842 13376 23848 13388
rect 23803 13348 23848 13376
rect 23842 13336 23848 13348
rect 23900 13336 23906 13388
rect 8996 13280 9904 13308
rect 11333 13311 11391 13317
rect 8996 13268 9002 13280
rect 11333 13277 11345 13311
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 2498 13200 2504 13252
rect 2556 13240 2562 13252
rect 2556 13212 3188 13240
rect 2556 13200 2562 13212
rect 2774 13172 2780 13184
rect 2735 13144 2780 13172
rect 2774 13132 2780 13144
rect 2832 13132 2838 13184
rect 3160 13181 3188 13212
rect 3145 13175 3203 13181
rect 3145 13141 3157 13175
rect 3191 13172 3203 13175
rect 3510 13172 3516 13184
rect 3191 13144 3516 13172
rect 3191 13141 3203 13144
rect 3145 13135 3203 13141
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 7098 13172 7104 13184
rect 7059 13144 7104 13172
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 9122 13132 9128 13184
rect 9180 13172 9186 13184
rect 9401 13175 9459 13181
rect 9401 13172 9413 13175
rect 9180 13144 9413 13172
rect 9180 13132 9186 13144
rect 9401 13141 9413 13144
rect 9447 13172 9459 13175
rect 9490 13172 9496 13184
rect 9447 13144 9496 13172
rect 9447 13141 9459 13144
rect 9401 13135 9459 13141
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 11146 13172 11152 13184
rect 11107 13144 11152 13172
rect 11146 13132 11152 13144
rect 11204 13172 11210 13184
rect 11348 13172 11376 13271
rect 11204 13144 11376 13172
rect 14277 13175 14335 13181
rect 11204 13132 11210 13144
rect 14277 13141 14289 13175
rect 14323 13172 14335 13175
rect 14366 13172 14372 13184
rect 14323 13144 14372 13172
rect 14323 13141 14335 13144
rect 14277 13135 14335 13141
rect 14366 13132 14372 13144
rect 14424 13132 14430 13184
rect 24854 13172 24860 13184
rect 24815 13144 24860 13172
rect 24854 13132 24860 13144
rect 24912 13132 24918 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 5353 12971 5411 12977
rect 5353 12968 5365 12971
rect 5224 12940 5365 12968
rect 5224 12928 5230 12940
rect 5353 12937 5365 12940
rect 5399 12937 5411 12971
rect 5353 12931 5411 12937
rect 6270 12928 6276 12980
rect 6328 12968 6334 12980
rect 7742 12968 7748 12980
rect 6328 12940 7748 12968
rect 6328 12928 6334 12940
rect 7742 12928 7748 12940
rect 7800 12968 7806 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7800 12940 7849 12968
rect 7800 12928 7806 12940
rect 7837 12937 7849 12940
rect 7883 12968 7895 12971
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 7883 12940 8217 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 8205 12931 8263 12937
rect 3786 12860 3792 12912
rect 3844 12900 3850 12912
rect 6457 12903 6515 12909
rect 6457 12900 6469 12903
rect 3844 12872 6469 12900
rect 3844 12860 3850 12872
rect 6457 12869 6469 12872
rect 6503 12900 6515 12903
rect 6549 12903 6607 12909
rect 6549 12900 6561 12903
rect 6503 12872 6561 12900
rect 6503 12869 6515 12872
rect 6457 12863 6515 12869
rect 6549 12869 6561 12872
rect 6595 12869 6607 12903
rect 6549 12863 6607 12869
rect 1854 12832 1860 12844
rect 1815 12804 1860 12832
rect 1854 12792 1860 12804
rect 1912 12792 1918 12844
rect 3559 12835 3617 12841
rect 3559 12801 3571 12835
rect 3605 12832 3617 12835
rect 5994 12832 6000 12844
rect 3605 12804 6000 12832
rect 3605 12801 3617 12804
rect 3559 12795 3617 12801
rect 5994 12792 6000 12804
rect 6052 12792 6058 12844
rect 6273 12835 6331 12841
rect 6273 12801 6285 12835
rect 6319 12832 6331 12835
rect 6319 12804 7420 12832
rect 6319 12801 6331 12804
rect 6273 12795 6331 12801
rect 7392 12776 7420 12804
rect 2501 12767 2559 12773
rect 2501 12733 2513 12767
rect 2547 12764 2559 12767
rect 2774 12764 2780 12776
rect 2547 12736 2780 12764
rect 2547 12733 2559 12736
rect 2501 12727 2559 12733
rect 2774 12724 2780 12736
rect 2832 12764 2838 12776
rect 2869 12767 2927 12773
rect 2869 12764 2881 12767
rect 2832 12736 2881 12764
rect 2832 12724 2838 12736
rect 2869 12733 2881 12736
rect 2915 12733 2927 12767
rect 2869 12727 2927 12733
rect 3050 12724 3056 12776
rect 3108 12764 3114 12776
rect 3456 12767 3514 12773
rect 3456 12764 3468 12767
rect 3108 12736 3468 12764
rect 3108 12724 3114 12736
rect 3456 12733 3468 12736
rect 3502 12764 3514 12767
rect 3881 12767 3939 12773
rect 3881 12764 3893 12767
rect 3502 12736 3893 12764
rect 3502 12733 3514 12736
rect 3456 12727 3514 12733
rect 3881 12733 3893 12736
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 4212 12736 4445 12764
rect 4212 12724 4218 12736
rect 4433 12733 4445 12736
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 6457 12767 6515 12773
rect 6457 12733 6469 12767
rect 6503 12764 6515 12767
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6503 12736 6837 12764
rect 6503 12733 6515 12736
rect 6457 12727 6515 12733
rect 6825 12733 6837 12736
rect 6871 12733 6883 12767
rect 7374 12764 7380 12776
rect 7335 12736 7380 12764
rect 6825 12727 6883 12733
rect 4341 12699 4399 12705
rect 4341 12696 4353 12699
rect 4126 12668 4353 12696
rect 1765 12631 1823 12637
rect 1765 12597 1777 12631
rect 1811 12628 1823 12631
rect 1946 12628 1952 12640
rect 1811 12600 1952 12628
rect 1811 12597 1823 12600
rect 1765 12591 1823 12597
rect 1946 12588 1952 12600
rect 2004 12628 2010 12640
rect 4126 12628 4154 12668
rect 4341 12665 4353 12668
rect 4387 12696 4399 12699
rect 4614 12696 4620 12708
rect 4387 12668 4620 12696
rect 4387 12665 4399 12668
rect 4341 12659 4399 12665
rect 4614 12656 4620 12668
rect 4672 12696 4678 12708
rect 4795 12699 4853 12705
rect 4795 12696 4807 12699
rect 4672 12668 4807 12696
rect 4672 12656 4678 12668
rect 4795 12665 4807 12668
rect 4841 12696 4853 12699
rect 6840 12696 6868 12727
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 8220 12764 8248 12931
rect 13357 12903 13415 12909
rect 13357 12869 13369 12903
rect 13403 12900 13415 12903
rect 18598 12900 18604 12912
rect 13403 12872 18604 12900
rect 13403 12869 13415 12872
rect 13357 12863 13415 12869
rect 18598 12860 18604 12872
rect 18656 12860 18662 12912
rect 9122 12832 9128 12844
rect 9083 12804 9128 12832
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 11146 12832 11152 12844
rect 11107 12804 11152 12832
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12832 12495 12835
rect 12526 12832 12532 12844
rect 12483 12804 12532 12832
rect 12483 12801 12495 12804
rect 12437 12795 12495 12801
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 14274 12832 14280 12844
rect 14235 12804 14280 12832
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 14550 12832 14556 12844
rect 14511 12804 14556 12832
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 23842 12832 23848 12844
rect 23803 12804 23848 12832
rect 23842 12792 23848 12804
rect 23900 12792 23906 12844
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 8220 12736 8401 12764
rect 8389 12733 8401 12736
rect 8435 12733 8447 12767
rect 8938 12764 8944 12776
rect 8899 12736 8944 12764
rect 8389 12727 8447 12733
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 10505 12767 10563 12773
rect 10505 12733 10517 12767
rect 10551 12733 10563 12767
rect 10962 12764 10968 12776
rect 10923 12736 10968 12764
rect 10505 12727 10563 12733
rect 9674 12696 9680 12708
rect 4841 12668 5764 12696
rect 6840 12668 9680 12696
rect 4841 12665 4853 12668
rect 4795 12659 4853 12665
rect 5736 12637 5764 12668
rect 9674 12656 9680 12668
rect 9732 12696 9738 12708
rect 10321 12699 10379 12705
rect 10321 12696 10333 12699
rect 9732 12668 10333 12696
rect 9732 12656 9738 12668
rect 10321 12665 10333 12668
rect 10367 12696 10379 12699
rect 10520 12696 10548 12727
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 12216 12736 13645 12764
rect 12216 12724 12222 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 12176 12696 12204 12724
rect 10367 12668 12204 12696
rect 12758 12699 12816 12705
rect 10367 12665 10379 12668
rect 10321 12659 10379 12665
rect 12758 12665 12770 12699
rect 12804 12665 12816 12699
rect 12758 12659 12816 12665
rect 2004 12600 4154 12628
rect 5721 12631 5779 12637
rect 2004 12588 2010 12600
rect 5721 12597 5733 12631
rect 5767 12628 5779 12631
rect 6638 12628 6644 12640
rect 5767 12600 6644 12628
rect 5767 12597 5779 12600
rect 5721 12591 5779 12597
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 7098 12628 7104 12640
rect 7059 12600 7104 12628
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 11514 12628 11520 12640
rect 11475 12600 11520 12628
rect 11514 12588 11520 12600
rect 11572 12628 11578 12640
rect 11698 12628 11704 12640
rect 11572 12600 11704 12628
rect 11572 12588 11578 12600
rect 11698 12588 11704 12600
rect 11756 12628 11762 12640
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 11756 12600 12173 12628
rect 11756 12588 11762 12600
rect 12161 12597 12173 12600
rect 12207 12628 12219 12631
rect 12773 12628 12801 12659
rect 12894 12656 12900 12708
rect 12952 12696 12958 12708
rect 13538 12696 13544 12708
rect 12952 12668 13544 12696
rect 12952 12656 12958 12668
rect 13538 12656 13544 12668
rect 13596 12696 13602 12708
rect 14001 12699 14059 12705
rect 14001 12696 14013 12699
rect 13596 12668 14013 12696
rect 13596 12656 13602 12668
rect 14001 12665 14013 12668
rect 14047 12665 14059 12699
rect 14366 12696 14372 12708
rect 14279 12668 14372 12696
rect 14001 12659 14059 12665
rect 14366 12656 14372 12668
rect 14424 12696 14430 12708
rect 15746 12696 15752 12708
rect 14424 12668 15752 12696
rect 14424 12656 14430 12668
rect 15746 12656 15752 12668
rect 15804 12656 15810 12708
rect 12207 12600 12801 12628
rect 12207 12597 12219 12600
rect 12161 12591 12219 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2590 12424 2596 12436
rect 2551 12396 2596 12424
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 4338 12424 4344 12436
rect 4299 12396 4344 12424
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 5166 12384 5172 12436
rect 5224 12424 5230 12436
rect 5997 12427 6055 12433
rect 5997 12424 6009 12427
rect 5224 12396 6009 12424
rect 5224 12384 5230 12396
rect 5997 12393 6009 12396
rect 6043 12393 6055 12427
rect 5997 12387 6055 12393
rect 10781 12427 10839 12433
rect 10781 12393 10793 12427
rect 10827 12424 10839 12427
rect 10962 12424 10968 12436
rect 10827 12396 10968 12424
rect 10827 12393 10839 12396
rect 10781 12387 10839 12393
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 12526 12424 12532 12436
rect 12487 12396 12532 12424
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 13170 12424 13176 12436
rect 13131 12396 13176 12424
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 14274 12384 14280 12436
rect 14332 12424 14338 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 14332 12396 14381 12424
rect 14332 12384 14338 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 6917 12359 6975 12365
rect 4126 12328 6868 12356
rect 4126 12300 4154 12328
rect 1670 12288 1676 12300
rect 1631 12260 1676 12288
rect 1670 12248 1676 12260
rect 1728 12248 1734 12300
rect 4062 12288 4068 12300
rect 4023 12260 4068 12288
rect 4062 12248 4068 12260
rect 4120 12260 4154 12300
rect 4893 12291 4951 12297
rect 4120 12248 4126 12260
rect 4893 12257 4905 12291
rect 4939 12257 4951 12291
rect 5074 12288 5080 12300
rect 5035 12260 5080 12288
rect 4893 12251 4951 12257
rect 3234 12180 3240 12232
rect 3292 12220 3298 12232
rect 4908 12220 4936 12251
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 6086 12248 6092 12300
rect 6144 12288 6150 12300
rect 6181 12291 6239 12297
rect 6181 12288 6193 12291
rect 6144 12260 6193 12288
rect 6144 12248 6150 12260
rect 6181 12257 6193 12260
rect 6227 12257 6239 12291
rect 6840 12288 6868 12328
rect 6917 12325 6929 12359
rect 6963 12356 6975 12359
rect 7374 12356 7380 12368
rect 6963 12328 7380 12356
rect 6963 12325 6975 12328
rect 6917 12319 6975 12325
rect 7374 12316 7380 12328
rect 7432 12316 7438 12368
rect 8757 12359 8815 12365
rect 8757 12325 8769 12359
rect 8803 12356 8815 12359
rect 8938 12356 8944 12368
rect 8803 12328 8944 12356
rect 8803 12325 8815 12328
rect 8757 12319 8815 12325
rect 8938 12316 8944 12328
rect 8996 12356 9002 12368
rect 9401 12359 9459 12365
rect 9401 12356 9413 12359
rect 8996 12328 9413 12356
rect 8996 12316 9002 12328
rect 9401 12325 9413 12328
rect 9447 12325 9459 12359
rect 9401 12319 9459 12325
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 6840 12260 7481 12288
rect 6181 12251 6239 12257
rect 7469 12257 7481 12260
rect 7515 12288 7527 12291
rect 8021 12291 8079 12297
rect 8021 12288 8033 12291
rect 7515 12260 8033 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 8021 12257 8033 12260
rect 8067 12288 8079 12291
rect 8662 12288 8668 12300
rect 8067 12260 8668 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 8662 12248 8668 12260
rect 8720 12248 8726 12300
rect 9674 12288 9680 12300
rect 9635 12260 9680 12288
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12257 11299 12291
rect 11241 12251 11299 12257
rect 3292 12192 5304 12220
rect 3292 12180 3298 12192
rect 5276 12152 5304 12192
rect 5442 12180 5448 12232
rect 5500 12220 5506 12232
rect 6546 12220 6552 12232
rect 5500 12192 6552 12220
rect 5500 12180 5506 12192
rect 6546 12180 6552 12192
rect 6604 12220 6610 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 6604 12192 8401 12220
rect 6604 12180 6610 12192
rect 8389 12189 8401 12192
rect 8435 12220 8447 12223
rect 8570 12220 8576 12232
rect 8435 12192 8576 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12220 10471 12223
rect 10594 12220 10600 12232
rect 10459 12192 10600 12220
rect 10459 12189 10471 12192
rect 10413 12183 10471 12189
rect 10594 12180 10600 12192
rect 10652 12220 10658 12232
rect 11057 12223 11115 12229
rect 11057 12220 11069 12223
rect 10652 12192 11069 12220
rect 10652 12180 10658 12192
rect 11057 12189 11069 12192
rect 11103 12189 11115 12223
rect 11256 12220 11284 12251
rect 11330 12248 11336 12300
rect 11388 12288 11394 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 11388 12260 11713 12288
rect 11388 12248 11394 12260
rect 11701 12257 11713 12260
rect 11747 12288 11759 12291
rect 12894 12288 12900 12300
rect 11747 12260 12900 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 12894 12248 12900 12260
rect 12952 12248 12958 12300
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 14366 12288 14372 12300
rect 13771 12260 14372 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 14366 12248 14372 12260
rect 14424 12248 14430 12300
rect 15746 12288 15752 12300
rect 15707 12260 15752 12288
rect 15746 12248 15752 12260
rect 15804 12248 15810 12300
rect 11790 12220 11796 12232
rect 11256 12192 11796 12220
rect 11057 12183 11115 12189
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12220 12035 12223
rect 12158 12220 12164 12232
rect 12023 12192 12164 12220
rect 12023 12189 12035 12192
rect 11977 12183 12035 12189
rect 12158 12180 12164 12192
rect 12216 12220 12222 12232
rect 12805 12223 12863 12229
rect 12805 12220 12817 12223
rect 12216 12192 12817 12220
rect 12216 12180 12222 12192
rect 12805 12189 12817 12192
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 13964 12192 15301 12220
rect 13964 12180 13970 12192
rect 15289 12189 15301 12192
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 6178 12152 6184 12164
rect 5276 12124 6184 12152
rect 6178 12112 6184 12124
rect 6236 12112 6242 12164
rect 6346 12155 6404 12161
rect 6346 12121 6358 12155
rect 6392 12152 6404 12155
rect 7282 12152 7288 12164
rect 6392 12124 7288 12152
rect 6392 12121 6404 12124
rect 6346 12115 6404 12121
rect 7282 12112 7288 12124
rect 7340 12152 7346 12164
rect 7837 12155 7895 12161
rect 7837 12152 7849 12155
rect 7340 12124 7849 12152
rect 7340 12112 7346 12124
rect 7837 12121 7849 12124
rect 7883 12152 7895 12155
rect 8159 12155 8217 12161
rect 8159 12152 8171 12155
rect 7883 12124 8171 12152
rect 7883 12121 7895 12124
rect 7837 12115 7895 12121
rect 8159 12121 8171 12124
rect 8205 12121 8217 12155
rect 11808 12152 11836 12180
rect 12986 12152 12992 12164
rect 11808 12124 12992 12152
rect 8159 12115 8217 12121
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 2038 12084 2044 12096
rect 1999 12056 2044 12084
rect 2038 12044 2044 12056
rect 2096 12044 2102 12096
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4154 12084 4160 12096
rect 3927 12056 4160 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4154 12044 4160 12056
rect 4212 12044 4218 12096
rect 5258 12044 5264 12096
rect 5316 12084 5322 12096
rect 6454 12084 6460 12096
rect 5316 12056 6460 12084
rect 5316 12044 5322 12056
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 8294 12084 8300 12096
rect 8255 12056 8300 12084
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 14090 12084 14096 12096
rect 14051 12056 14096 12084
rect 14090 12044 14096 12056
rect 14148 12044 14154 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 3513 11883 3571 11889
rect 3513 11880 3525 11883
rect 3292 11852 3525 11880
rect 3292 11840 3298 11852
rect 3513 11849 3525 11852
rect 3559 11849 3571 11883
rect 6546 11880 6552 11892
rect 6507 11852 6552 11880
rect 3513 11843 3571 11849
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 8570 11880 8576 11892
rect 8531 11852 8576 11880
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 9674 11880 9680 11892
rect 9635 11852 9680 11880
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 10134 11880 10140 11892
rect 10095 11852 10140 11880
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11882 11880 11888 11892
rect 11563 11852 11888 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 15746 11880 15752 11892
rect 15707 11852 15752 11880
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 24210 11840 24216 11892
rect 24268 11880 24274 11892
rect 24719 11883 24777 11889
rect 24719 11880 24731 11883
rect 24268 11852 24731 11880
rect 24268 11840 24274 11852
rect 24719 11849 24731 11852
rect 24765 11849 24777 11883
rect 24719 11843 24777 11849
rect 1762 11772 1768 11824
rect 1820 11812 1826 11824
rect 2777 11815 2835 11821
rect 2777 11812 2789 11815
rect 1820 11784 2789 11812
rect 1820 11772 1826 11784
rect 1872 11753 1900 11784
rect 2777 11781 2789 11784
rect 2823 11781 2835 11815
rect 2777 11775 2835 11781
rect 7834 11772 7840 11824
rect 7892 11812 7898 11824
rect 8018 11812 8024 11824
rect 7892 11784 8024 11812
rect 7892 11772 7898 11784
rect 8018 11772 8024 11784
rect 8076 11812 8082 11824
rect 8205 11815 8263 11821
rect 8205 11812 8217 11815
rect 8076 11784 8217 11812
rect 8076 11772 8082 11784
rect 8205 11781 8217 11784
rect 8251 11781 8263 11815
rect 8205 11775 8263 11781
rect 12802 11772 12808 11824
rect 12860 11812 12866 11824
rect 14369 11815 14427 11821
rect 14369 11812 14381 11815
rect 12860 11784 14381 11812
rect 12860 11772 12866 11784
rect 14369 11781 14381 11784
rect 14415 11812 14427 11815
rect 14550 11812 14556 11824
rect 14415 11784 14556 11812
rect 14415 11781 14427 11784
rect 14369 11775 14427 11781
rect 14550 11772 14556 11784
rect 14608 11772 14614 11824
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11713 1915 11747
rect 1857 11707 1915 11713
rect 3786 11704 3792 11756
rect 3844 11744 3850 11756
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3844 11716 3985 11744
rect 3844 11704 3850 11716
rect 3973 11713 3985 11716
rect 4019 11744 4031 11747
rect 4019 11716 4936 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 4908 11688 4936 11716
rect 7190 11704 7196 11756
rect 7248 11744 7254 11756
rect 7653 11747 7711 11753
rect 7653 11744 7665 11747
rect 7248 11716 7665 11744
rect 7248 11704 7254 11716
rect 7653 11713 7665 11716
rect 7699 11744 7711 11747
rect 9125 11747 9183 11753
rect 9125 11744 9137 11747
rect 7699 11716 9137 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 9125 11713 9137 11716
rect 9171 11713 9183 11747
rect 10594 11744 10600 11756
rect 10555 11716 10600 11744
rect 9125 11707 9183 11713
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 12820 11744 12848 11772
rect 12795 11716 12848 11744
rect 13817 11747 13875 11753
rect 4062 11676 4068 11688
rect 4023 11648 4068 11676
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4890 11676 4896 11688
rect 4803 11648 4896 11676
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5074 11676 5080 11688
rect 4987 11648 5080 11676
rect 5074 11636 5080 11648
rect 5132 11676 5138 11688
rect 11882 11676 11888 11688
rect 5132 11648 5396 11676
rect 11843 11648 11888 11676
rect 5132 11636 5138 11648
rect 1949 11611 2007 11617
rect 1949 11577 1961 11611
rect 1995 11577 2007 11611
rect 2498 11608 2504 11620
rect 2459 11580 2504 11608
rect 1949 11571 2007 11577
rect 1670 11540 1676 11552
rect 1631 11512 1676 11540
rect 1670 11500 1676 11512
rect 1728 11540 1734 11552
rect 1964 11540 1992 11571
rect 2498 11568 2504 11580
rect 2556 11568 2562 11620
rect 5368 11552 5396 11648
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 12795 11685 12823 11716
rect 13817 11713 13829 11747
rect 13863 11744 13875 11747
rect 14090 11744 14096 11756
rect 13863 11716 14096 11744
rect 13863 11713 13875 11716
rect 13817 11707 13875 11713
rect 14090 11704 14096 11716
rect 14148 11744 14154 11756
rect 15289 11747 15347 11753
rect 15289 11744 15301 11747
rect 14148 11716 15301 11744
rect 14148 11704 14154 11716
rect 15289 11713 15301 11716
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 12780 11679 12838 11685
rect 12780 11645 12792 11679
rect 12826 11645 12838 11679
rect 12780 11639 12838 11645
rect 24648 11679 24706 11685
rect 24648 11645 24660 11679
rect 24694 11676 24706 11679
rect 24694 11648 25176 11676
rect 24694 11645 24706 11648
rect 24648 11639 24706 11645
rect 7745 11611 7803 11617
rect 7745 11577 7757 11611
rect 7791 11608 7803 11611
rect 7834 11608 7840 11620
rect 7791 11580 7840 11608
rect 7791 11577 7803 11580
rect 7745 11571 7803 11577
rect 1728 11512 1992 11540
rect 1728 11500 1734 11512
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 3142 11540 3148 11552
rect 2372 11512 3148 11540
rect 2372 11500 2378 11512
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 4212 11512 4257 11540
rect 4212 11500 4218 11512
rect 5350 11500 5356 11552
rect 5408 11540 5414 11552
rect 5445 11543 5503 11549
rect 5445 11540 5457 11543
rect 5408 11512 5457 11540
rect 5408 11500 5414 11512
rect 5445 11509 5457 11512
rect 5491 11509 5503 11543
rect 5902 11540 5908 11552
rect 5863 11512 5908 11540
rect 5445 11503 5503 11509
rect 5902 11500 5908 11512
rect 5960 11540 5966 11552
rect 6086 11540 6092 11552
rect 5960 11512 6092 11540
rect 5960 11500 5966 11512
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 6270 11540 6276 11552
rect 6231 11512 6276 11540
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 7101 11543 7159 11549
rect 7101 11509 7113 11543
rect 7147 11540 7159 11543
rect 7282 11540 7288 11552
rect 7147 11512 7288 11540
rect 7147 11509 7159 11512
rect 7101 11503 7159 11509
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 7469 11543 7527 11549
rect 7469 11509 7481 11543
rect 7515 11540 7527 11543
rect 7760 11540 7788 11571
rect 7834 11568 7840 11580
rect 7892 11568 7898 11620
rect 10959 11611 11017 11617
rect 10959 11577 10971 11611
rect 11005 11608 11017 11611
rect 11514 11608 11520 11620
rect 11005 11580 11520 11608
rect 11005 11577 11017 11580
rect 10959 11571 11017 11577
rect 7515 11512 7788 11540
rect 7515 11509 7527 11512
rect 7469 11503 7527 11509
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8352 11512 9045 11540
rect 8352 11500 8358 11512
rect 9033 11509 9045 11512
rect 9079 11540 9091 11543
rect 9766 11540 9772 11552
rect 9079 11512 9772 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11540 10563 11543
rect 10974 11540 11002 11571
rect 11514 11568 11520 11580
rect 11572 11608 11578 11620
rect 12989 11611 13047 11617
rect 11572 11580 11928 11608
rect 11572 11568 11578 11580
rect 11146 11540 11152 11552
rect 10551 11512 11152 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 11900 11540 11928 11580
rect 12989 11577 13001 11611
rect 13035 11608 13047 11611
rect 13538 11608 13544 11620
rect 13035 11580 13544 11608
rect 13035 11577 13047 11580
rect 12989 11571 13047 11577
rect 13538 11568 13544 11580
rect 13596 11568 13602 11620
rect 13633 11611 13691 11617
rect 13633 11577 13645 11611
rect 13679 11608 13691 11611
rect 13906 11608 13912 11620
rect 13679 11580 13912 11608
rect 13679 11577 13691 11580
rect 13633 11571 13691 11577
rect 13906 11568 13912 11580
rect 13964 11568 13970 11620
rect 13170 11540 13176 11552
rect 11900 11512 13176 11540
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 25148 11549 25176 11648
rect 25133 11543 25191 11549
rect 25133 11509 25145 11543
rect 25179 11540 25191 11543
rect 27614 11540 27620 11552
rect 25179 11512 27620 11540
rect 25179 11509 25191 11512
rect 25133 11503 25191 11509
rect 27614 11500 27620 11512
rect 27672 11500 27678 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 4062 11336 4068 11348
rect 3200 11308 4068 11336
rect 3200 11296 3206 11308
rect 4062 11296 4068 11308
rect 4120 11336 4126 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4120 11308 4537 11336
rect 4120 11296 4126 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 7190 11336 7196 11348
rect 7151 11308 7196 11336
rect 4525 11299 4583 11305
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 10321 11339 10379 11345
rect 10321 11305 10333 11339
rect 10367 11336 10379 11339
rect 10781 11339 10839 11345
rect 10781 11336 10793 11339
rect 10367 11308 10793 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 10781 11305 10793 11308
rect 10827 11336 10839 11339
rect 10962 11336 10968 11348
rect 10827 11308 10968 11336
rect 10827 11305 10839 11308
rect 10781 11299 10839 11305
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 12713 11339 12771 11345
rect 12713 11305 12725 11339
rect 12759 11336 12771 11339
rect 12802 11336 12808 11348
rect 12759 11308 12808 11336
rect 12759 11305 12771 11308
rect 12713 11299 12771 11305
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13078 11296 13084 11348
rect 13136 11336 13142 11348
rect 13136 11308 13400 11336
rect 13136 11296 13142 11308
rect 1949 11271 2007 11277
rect 1949 11237 1961 11271
rect 1995 11268 2007 11271
rect 2038 11268 2044 11280
rect 1995 11240 2044 11268
rect 1995 11237 2007 11240
rect 1949 11231 2007 11237
rect 2038 11228 2044 11240
rect 2096 11228 2102 11280
rect 2498 11268 2504 11280
rect 2459 11240 2504 11268
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 5902 11268 5908 11280
rect 5644 11240 5908 11268
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4100 11203 4158 11209
rect 4100 11200 4112 11203
rect 4028 11172 4112 11200
rect 4028 11160 4034 11172
rect 4100 11169 4112 11172
rect 4146 11169 4158 11203
rect 4100 11163 4158 11169
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5644 11209 5672 11240
rect 5902 11228 5908 11240
rect 5960 11268 5966 11280
rect 7466 11268 7472 11280
rect 5960 11240 6776 11268
rect 7427 11240 7472 11268
rect 5960 11228 5966 11240
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 5316 11172 5641 11200
rect 5316 11160 5322 11172
rect 5629 11169 5641 11172
rect 5675 11169 5687 11203
rect 5629 11163 5687 11169
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 6178 11200 6184 11212
rect 6139 11172 6184 11200
rect 5813 11163 5871 11169
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 5828 11132 5856 11163
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 1903 11104 2912 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 2884 11073 2912 11104
rect 5368 11104 5856 11132
rect 2869 11067 2927 11073
rect 2869 11033 2881 11067
rect 2915 11064 2927 11067
rect 4203 11067 4261 11073
rect 4203 11064 4215 11067
rect 2915 11036 4215 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 4203 11033 4215 11036
rect 4249 11033 4261 11067
rect 4203 11027 4261 11033
rect 5368 11008 5396 11104
rect 6748 11064 6776 11240
rect 7466 11228 7472 11240
rect 7524 11228 7530 11280
rect 8018 11268 8024 11280
rect 7979 11240 8024 11268
rect 8018 11228 8024 11240
rect 8076 11228 8082 11280
rect 11146 11228 11152 11280
rect 11204 11268 11210 11280
rect 11746 11271 11804 11277
rect 11746 11268 11758 11271
rect 11204 11240 11758 11268
rect 11204 11228 11210 11240
rect 11746 11237 11758 11240
rect 11792 11237 11804 11271
rect 13262 11268 13268 11280
rect 13223 11240 13268 11268
rect 11746 11231 11804 11237
rect 13262 11228 13268 11240
rect 13320 11228 13326 11280
rect 13372 11277 13400 11308
rect 13357 11271 13415 11277
rect 13357 11237 13369 11271
rect 13403 11237 13415 11271
rect 13357 11231 13415 11237
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 9723 11172 10180 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11132 6883 11135
rect 7006 11132 7012 11144
rect 6871 11104 7012 11132
rect 6871 11101 6883 11104
rect 6825 11095 6883 11101
rect 7006 11092 7012 11104
rect 7064 11132 7070 11144
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7064 11104 7389 11132
rect 7064 11092 7070 11104
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 9824 11135 9882 11141
rect 9824 11132 9836 11135
rect 9456 11104 9836 11132
rect 9456 11092 9462 11104
rect 9824 11101 9836 11104
rect 9870 11101 9882 11135
rect 10042 11132 10048 11144
rect 10003 11104 10048 11132
rect 9824 11095 9882 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 9030 11064 9036 11076
rect 6748 11036 9036 11064
rect 9030 11024 9036 11036
rect 9088 11064 9094 11076
rect 9493 11067 9551 11073
rect 9493 11064 9505 11067
rect 9088 11036 9505 11064
rect 9088 11024 9094 11036
rect 9493 11033 9505 11036
rect 9539 11064 9551 11067
rect 10152 11064 10180 11172
rect 11422 11132 11428 11144
rect 11383 11104 11428 11132
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 12710 11064 12716 11076
rect 9539 11036 12716 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 13170 11024 13176 11076
rect 13228 11064 13234 11076
rect 13556 11064 13584 11095
rect 13228 11036 13584 11064
rect 13228 11024 13234 11036
rect 1670 10996 1676 11008
rect 1631 10968 1676 10996
rect 1670 10956 1676 10968
rect 1728 10956 1734 11008
rect 3605 10999 3663 11005
rect 3605 10965 3617 10999
rect 3651 10996 3663 10999
rect 3694 10996 3700 11008
rect 3651 10968 3700 10996
rect 3651 10965 3663 10968
rect 3605 10959 3663 10965
rect 3694 10956 3700 10968
rect 3752 10956 3758 11008
rect 4985 10999 5043 11005
rect 4985 10965 4997 10999
rect 5031 10996 5043 10999
rect 5350 10996 5356 11008
rect 5031 10968 5356 10996
rect 5031 10965 5043 10968
rect 4985 10959 5043 10965
rect 5350 10956 5356 10968
rect 5408 10956 5414 11008
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 6512 10968 6557 10996
rect 6512 10956 6518 10968
rect 9766 10956 9772 11008
rect 9824 10996 9830 11008
rect 9953 10999 10011 11005
rect 9953 10996 9965 10999
rect 9824 10968 9965 10996
rect 9824 10956 9830 10968
rect 9953 10965 9965 10968
rect 9999 10965 10011 10999
rect 11238 10996 11244 11008
rect 11199 10968 11244 10996
rect 9953 10959 10011 10965
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 12345 10999 12403 11005
rect 12345 10965 12357 10999
rect 12391 10996 12403 10999
rect 13078 10996 13084 11008
rect 12391 10968 13084 10996
rect 12391 10965 12403 10968
rect 12345 10959 12403 10965
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14185 10999 14243 11005
rect 14185 10996 14197 10999
rect 13872 10968 14197 10996
rect 13872 10956 13878 10968
rect 14185 10965 14197 10968
rect 14231 10965 14243 10999
rect 14185 10959 14243 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 1728 10764 2513 10792
rect 1728 10752 1734 10764
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 2501 10755 2559 10761
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4028 10764 4537 10792
rect 4028 10752 4034 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4525 10755 4583 10761
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 11238 10792 11244 10804
rect 9263 10764 11244 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 14458 10792 14464 10804
rect 13464 10764 14320 10792
rect 14419 10764 14464 10792
rect 6270 10684 6276 10736
rect 6328 10724 6334 10736
rect 8846 10724 8852 10736
rect 6328 10696 8852 10724
rect 6328 10684 6334 10696
rect 8846 10684 8852 10696
rect 8904 10684 8910 10736
rect 9766 10684 9772 10736
rect 9824 10724 9830 10736
rect 10137 10727 10195 10733
rect 10137 10724 10149 10727
rect 9824 10696 10149 10724
rect 9824 10684 9830 10696
rect 10137 10693 10149 10696
rect 10183 10724 10195 10727
rect 13464 10724 13492 10764
rect 14292 10736 14320 10764
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 10183 10696 13492 10724
rect 10183 10693 10195 10696
rect 10137 10687 10195 10693
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 14139 10727 14197 10733
rect 14139 10724 14151 10727
rect 13872 10696 14151 10724
rect 13872 10684 13878 10696
rect 14139 10693 14151 10696
rect 14185 10693 14197 10727
rect 14274 10724 14280 10736
rect 14235 10696 14280 10724
rect 14139 10687 14197 10693
rect 14274 10684 14280 10696
rect 14332 10684 14338 10736
rect 2498 10616 2504 10668
rect 2556 10656 2562 10668
rect 3602 10656 3608 10668
rect 2556 10628 3608 10656
rect 2556 10616 2562 10628
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 4798 10656 4804 10668
rect 4295 10628 4804 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 6454 10616 6460 10668
rect 6512 10656 6518 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6512 10628 6837 10656
rect 6512 10616 6518 10628
rect 6825 10625 6837 10628
rect 6871 10656 6883 10659
rect 7650 10656 7656 10668
rect 6871 10628 7656 10656
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8628 10628 8953 10656
rect 8628 10616 8634 10628
rect 8941 10625 8953 10628
rect 8987 10656 8999 10659
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 8987 10628 9689 10656
rect 8987 10625 8999 10628
rect 8941 10619 8999 10625
rect 9677 10625 9689 10628
rect 9723 10656 9735 10659
rect 10042 10656 10048 10668
rect 9723 10628 10048 10656
rect 9723 10625 9735 10628
rect 9677 10619 9735 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 11241 10659 11299 10665
rect 11241 10625 11253 10659
rect 11287 10656 11299 10659
rect 11422 10656 11428 10668
rect 11287 10628 11428 10656
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 14366 10616 14372 10668
rect 14424 10656 14430 10668
rect 14424 10628 14469 10656
rect 14424 10616 14430 10628
rect 1581 10591 1639 10597
rect 1581 10557 1593 10591
rect 1627 10588 1639 10591
rect 1762 10588 1768 10600
rect 1627 10560 1768 10588
rect 1627 10557 1639 10560
rect 1581 10551 1639 10557
rect 1762 10548 1768 10560
rect 1820 10588 1826 10600
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 1820 10560 3157 10588
rect 1820 10548 1826 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 5718 10588 5724 10600
rect 3145 10551 3203 10557
rect 4356 10560 5724 10588
rect 3694 10480 3700 10532
rect 3752 10520 3758 10532
rect 3752 10492 4154 10520
rect 3752 10480 3758 10492
rect 1946 10452 1952 10464
rect 1907 10424 1952 10452
rect 1946 10412 1952 10424
rect 2004 10412 2010 10464
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 2777 10455 2835 10461
rect 2777 10452 2789 10455
rect 2188 10424 2789 10452
rect 2188 10412 2194 10424
rect 2777 10421 2789 10424
rect 2823 10421 2835 10455
rect 4126 10452 4154 10492
rect 4356 10452 4384 10560
rect 5718 10548 5724 10560
rect 5776 10548 5782 10600
rect 7466 10548 7472 10600
rect 7524 10588 7530 10600
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7524 10560 7757 10588
rect 7524 10548 7530 10560
rect 7745 10557 7757 10560
rect 7791 10588 7803 10591
rect 8294 10588 8300 10600
rect 7791 10560 8300 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 8720 10591 8778 10597
rect 8720 10588 8732 10591
rect 8404 10560 8732 10588
rect 5074 10520 5080 10532
rect 5035 10492 5080 10520
rect 5074 10480 5080 10492
rect 5132 10480 5138 10532
rect 7146 10523 7204 10529
rect 7146 10520 7158 10523
rect 6656 10492 7158 10520
rect 6656 10464 6684 10492
rect 7146 10489 7158 10492
rect 7192 10489 7204 10523
rect 7146 10483 7204 10489
rect 7282 10480 7288 10532
rect 7340 10520 7346 10532
rect 8404 10520 8432 10560
rect 8720 10557 8732 10560
rect 8766 10557 8778 10591
rect 10686 10588 10692 10600
rect 10647 10560 10692 10588
rect 8720 10551 8778 10557
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 10962 10588 10968 10600
rect 10923 10560 10968 10588
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 8570 10520 8576 10532
rect 7340 10492 8432 10520
rect 8531 10492 8576 10520
rect 7340 10480 7346 10492
rect 8036 10464 8064 10492
rect 8570 10480 8576 10492
rect 8628 10480 8634 10532
rect 12526 10520 12532 10532
rect 12487 10492 12532 10520
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 13170 10520 13176 10532
rect 12676 10492 12721 10520
rect 13131 10492 13176 10520
rect 12676 10480 12682 10492
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 13541 10523 13599 10529
rect 13541 10489 13553 10523
rect 13587 10520 13599 10523
rect 13722 10520 13728 10532
rect 13587 10492 13728 10520
rect 13587 10489 13599 10492
rect 13541 10483 13599 10489
rect 4126 10424 4384 10452
rect 4985 10455 5043 10461
rect 2777 10415 2835 10421
rect 4985 10421 4997 10455
rect 5031 10452 5043 10455
rect 5258 10452 5264 10464
rect 5031 10424 5264 10452
rect 5031 10421 5043 10424
rect 4985 10415 5043 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 6089 10455 6147 10461
rect 6089 10452 6101 10455
rect 5500 10424 6101 10452
rect 5500 10412 5506 10424
rect 6089 10421 6101 10424
rect 6135 10452 6147 10455
rect 6178 10452 6184 10464
rect 6135 10424 6184 10452
rect 6135 10421 6147 10424
rect 6089 10415 6147 10421
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6638 10452 6644 10464
rect 6599 10424 6644 10452
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 8018 10452 8024 10464
rect 7979 10424 8024 10452
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 8481 10455 8539 10461
rect 8481 10421 8493 10455
rect 8527 10452 8539 10455
rect 8846 10452 8852 10464
rect 8527 10424 8852 10452
rect 8527 10421 8539 10424
rect 8481 10415 8539 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 11204 10424 11529 10452
rect 11204 10412 11210 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 11517 10415 11575 10421
rect 12253 10455 12311 10461
rect 12253 10421 12265 10455
rect 12299 10452 12311 10455
rect 12636 10452 12664 10480
rect 12299 10424 12664 10452
rect 12299 10421 12311 10424
rect 12253 10415 12311 10421
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 13556 10452 13584 10483
rect 13722 10480 13728 10492
rect 13780 10480 13786 10532
rect 13998 10520 14004 10532
rect 13959 10492 14004 10520
rect 13998 10480 14004 10492
rect 14056 10480 14062 10532
rect 12768 10424 13584 10452
rect 12768 10412 12774 10424
rect 13630 10412 13636 10464
rect 13688 10452 13694 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13688 10424 13829 10452
rect 13688 10412 13694 10424
rect 13817 10421 13829 10424
rect 13863 10452 13875 10455
rect 14366 10452 14372 10464
rect 13863 10424 14372 10452
rect 13863 10421 13875 10424
rect 13817 10415 13875 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2038 10248 2044 10260
rect 1999 10220 2044 10248
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 2961 10251 3019 10257
rect 2961 10248 2973 10251
rect 2924 10220 2973 10248
rect 2924 10208 2930 10220
rect 2961 10217 2973 10220
rect 3007 10217 3019 10251
rect 2961 10211 3019 10217
rect 3602 10208 3608 10260
rect 3660 10248 3666 10260
rect 3697 10251 3755 10257
rect 3697 10248 3709 10251
rect 3660 10220 3709 10248
rect 3660 10208 3666 10220
rect 3697 10217 3709 10220
rect 3743 10217 3755 10251
rect 5718 10248 5724 10260
rect 5679 10220 5724 10248
rect 3697 10211 3755 10217
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6089 10251 6147 10257
rect 6089 10248 6101 10251
rect 6052 10220 6101 10248
rect 6052 10208 6058 10220
rect 6089 10217 6101 10220
rect 6135 10217 6147 10251
rect 7650 10248 7656 10260
rect 7611 10220 7656 10248
rect 6089 10211 6147 10217
rect 3421 10183 3479 10189
rect 3421 10149 3433 10183
rect 3467 10180 3479 10183
rect 3878 10180 3884 10192
rect 3467 10152 3884 10180
rect 3467 10149 3479 10152
rect 3421 10143 3479 10149
rect 2130 10072 2136 10124
rect 2188 10112 2194 10124
rect 2317 10115 2375 10121
rect 2317 10112 2329 10115
rect 2188 10084 2329 10112
rect 2188 10072 2194 10084
rect 2317 10081 2329 10084
rect 2363 10081 2375 10115
rect 2317 10075 2375 10081
rect 2464 10115 2522 10121
rect 2464 10081 2476 10115
rect 2510 10112 2522 10115
rect 3436 10112 3464 10143
rect 3878 10140 3884 10152
rect 3936 10140 3942 10192
rect 4246 10180 4252 10192
rect 4159 10152 4252 10180
rect 4246 10140 4252 10152
rect 4304 10180 4310 10192
rect 5074 10180 5080 10192
rect 4304 10152 5080 10180
rect 4304 10140 4310 10152
rect 5074 10140 5080 10152
rect 5132 10140 5138 10192
rect 2510 10084 3464 10112
rect 2510 10081 2522 10084
rect 2464 10075 2522 10081
rect 2682 10044 2688 10056
rect 2643 10016 2688 10044
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4430 10044 4436 10056
rect 4203 10016 4436 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4430 10004 4436 10016
rect 4488 10004 4494 10056
rect 4798 10044 4804 10056
rect 4759 10016 4804 10044
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 6104 10044 6132 10211
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 8662 10208 8668 10260
rect 8720 10248 8726 10260
rect 8849 10251 8907 10257
rect 8849 10248 8861 10251
rect 8720 10220 8861 10248
rect 8720 10208 8726 10220
rect 8849 10217 8861 10220
rect 8895 10217 8907 10251
rect 8849 10211 8907 10217
rect 11333 10251 11391 10257
rect 11333 10217 11345 10251
rect 11379 10248 11391 10251
rect 11422 10248 11428 10260
rect 11379 10220 11428 10248
rect 11379 10217 11391 10220
rect 11333 10211 11391 10217
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 12897 10251 12955 10257
rect 12897 10217 12909 10251
rect 12943 10248 12955 10251
rect 13262 10248 13268 10260
rect 12943 10220 13268 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13722 10208 13728 10260
rect 13780 10248 13786 10260
rect 13998 10248 14004 10260
rect 13780 10220 14004 10248
rect 13780 10208 13786 10220
rect 13998 10208 14004 10220
rect 14056 10248 14062 10260
rect 15378 10248 15384 10260
rect 14056 10220 15384 10248
rect 14056 10208 14062 10220
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 6454 10180 6460 10192
rect 6415 10152 6460 10180
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 7006 10180 7012 10192
rect 6967 10152 7012 10180
rect 7006 10140 7012 10152
rect 7064 10140 7070 10192
rect 7834 10180 7840 10192
rect 7795 10152 7840 10180
rect 7834 10140 7840 10152
rect 7892 10140 7898 10192
rect 11514 10180 11520 10192
rect 11475 10152 11520 10180
rect 11514 10140 11520 10152
rect 11572 10140 11578 10192
rect 11606 10140 11612 10192
rect 11664 10180 11670 10192
rect 11664 10152 11709 10180
rect 11664 10140 11670 10152
rect 12618 10140 12624 10192
rect 12676 10180 12682 10192
rect 12989 10183 13047 10189
rect 12989 10180 13001 10183
rect 12676 10152 13001 10180
rect 12676 10140 12682 10152
rect 12989 10149 13001 10152
rect 13035 10149 13047 10183
rect 12989 10143 13047 10149
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 8294 10112 8300 10124
rect 7423 10084 8300 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 9858 10112 9864 10124
rect 9819 10084 9864 10112
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 10134 10112 10140 10124
rect 10095 10084 10140 10112
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 13078 10112 13084 10124
rect 13039 10084 13084 10112
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 13170 10072 13176 10124
rect 13228 10112 13234 10124
rect 15286 10112 15292 10124
rect 15344 10121 15350 10124
rect 15344 10115 15382 10121
rect 13228 10084 15292 10112
rect 13228 10072 13234 10084
rect 15286 10072 15292 10084
rect 15370 10081 15382 10115
rect 15344 10075 15382 10081
rect 15344 10072 15350 10075
rect 6365 10047 6423 10053
rect 6365 10044 6377 10047
rect 6104 10016 6377 10044
rect 6365 10013 6377 10016
rect 6411 10013 6423 10047
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 6365 10007 6423 10013
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 11790 10044 11796 10056
rect 11751 10016 11796 10044
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12526 10044 12532 10056
rect 12439 10016 12532 10044
rect 12526 10004 12532 10016
rect 12584 10044 12590 10056
rect 15562 10044 15568 10056
rect 12584 10016 15568 10044
rect 12584 10004 12590 10016
rect 15562 10004 15568 10016
rect 15620 10004 15626 10056
rect 6270 9976 6276 9988
rect 2608 9948 6276 9976
rect 2608 9920 2636 9948
rect 6270 9936 6276 9948
rect 6328 9936 6334 9988
rect 1673 9911 1731 9917
rect 1673 9877 1685 9911
rect 1719 9908 1731 9911
rect 2038 9908 2044 9920
rect 1719 9880 2044 9908
rect 1719 9877 1731 9880
rect 1673 9871 1731 9877
rect 2038 9868 2044 9880
rect 2096 9868 2102 9920
rect 2590 9908 2596 9920
rect 2551 9880 2596 9908
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 5350 9908 5356 9920
rect 5311 9880 5356 9908
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 9398 9908 9404 9920
rect 9359 9880 9404 9908
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 10686 9908 10692 9920
rect 10647 9880 10692 9908
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 14090 9908 14096 9920
rect 14051 9880 14096 9908
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14458 9868 14464 9920
rect 14516 9908 14522 9920
rect 15427 9911 15485 9917
rect 15427 9908 15439 9911
rect 14516 9880 15439 9908
rect 14516 9868 14522 9880
rect 15427 9877 15439 9880
rect 15473 9877 15485 9911
rect 15427 9871 15485 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 2685 9707 2743 9713
rect 2685 9704 2697 9707
rect 2648 9676 2697 9704
rect 2648 9664 2654 9676
rect 2685 9673 2697 9676
rect 2731 9673 2743 9707
rect 2685 9667 2743 9673
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 3789 9707 3847 9713
rect 3789 9704 3801 9707
rect 3752 9676 3801 9704
rect 3752 9664 3758 9676
rect 3789 9673 3801 9676
rect 3835 9673 3847 9707
rect 3789 9667 3847 9673
rect 4065 9707 4123 9713
rect 4065 9673 4077 9707
rect 4111 9704 4123 9707
rect 4246 9704 4252 9716
rect 4111 9676 4252 9704
rect 4111 9673 4123 9676
rect 4065 9667 4123 9673
rect 4246 9664 4252 9676
rect 4304 9664 4310 9716
rect 4430 9704 4436 9716
rect 4391 9676 4436 9704
rect 4430 9664 4436 9676
rect 4488 9664 4494 9716
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 9858 9704 9864 9716
rect 9815 9676 9864 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 9858 9664 9864 9676
rect 9916 9704 9922 9716
rect 10686 9704 10692 9716
rect 9916 9676 10692 9704
rect 9916 9664 9922 9676
rect 10686 9664 10692 9676
rect 10744 9704 10750 9716
rect 11882 9704 11888 9716
rect 10744 9676 11888 9704
rect 10744 9664 10750 9676
rect 11882 9664 11888 9676
rect 11940 9664 11946 9716
rect 12250 9704 12256 9716
rect 12211 9676 12256 9704
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 13136 9676 13461 9704
rect 13136 9664 13142 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 15286 9704 15292 9716
rect 15247 9676 15292 9704
rect 13449 9667 13507 9673
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 8386 9596 8392 9648
rect 8444 9636 8450 9648
rect 8846 9636 8852 9648
rect 8444 9608 8852 9636
rect 8444 9596 8450 9608
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 10962 9596 10968 9648
rect 11020 9636 11026 9648
rect 13814 9636 13820 9648
rect 11020 9608 13820 9636
rect 11020 9596 11026 9608
rect 13814 9596 13820 9608
rect 13872 9636 13878 9648
rect 14826 9636 14832 9648
rect 13872 9608 14832 9636
rect 13872 9596 13878 9608
rect 14826 9596 14832 9608
rect 14884 9596 14890 9648
rect 1486 9528 1492 9580
rect 1544 9568 1550 9580
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 1544 9540 2881 9568
rect 1544 9528 1550 9540
rect 2869 9537 2881 9540
rect 2915 9568 2927 9571
rect 3510 9568 3516 9580
rect 2915 9540 3516 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 6273 9571 6331 9577
rect 6273 9568 6285 9571
rect 5951 9540 6285 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 6273 9537 6285 9540
rect 6319 9568 6331 9571
rect 6454 9568 6460 9580
rect 6319 9540 6460 9568
rect 6319 9537 6331 9540
rect 6273 9531 6331 9537
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 7064 9540 7205 9568
rect 7064 9528 7070 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 8570 9528 8576 9580
rect 8628 9568 8634 9580
rect 8941 9571 8999 9577
rect 8941 9568 8953 9571
rect 8628 9540 8953 9568
rect 8628 9528 8634 9540
rect 8941 9537 8953 9540
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9568 9367 9571
rect 10134 9568 10140 9580
rect 9355 9540 10140 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10318 9568 10324 9580
rect 10279 9540 10324 9568
rect 10318 9528 10324 9540
rect 10376 9568 10382 9580
rect 10686 9568 10692 9580
rect 10376 9540 10692 9568
rect 10376 9528 10382 9540
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 14642 9568 14648 9580
rect 12452 9540 14648 9568
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 5077 9503 5135 9509
rect 1719 9472 2452 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 1489 9435 1547 9441
rect 1489 9401 1501 9435
rect 1535 9432 1547 9435
rect 1578 9432 1584 9444
rect 1535 9404 1584 9432
rect 1535 9401 1547 9404
rect 1489 9395 1547 9401
rect 1578 9392 1584 9404
rect 1636 9392 1642 9444
rect 2041 9435 2099 9441
rect 2041 9401 2053 9435
rect 2087 9432 2099 9435
rect 2314 9432 2320 9444
rect 2087 9404 2320 9432
rect 2087 9401 2099 9404
rect 2041 9395 2099 9401
rect 2314 9392 2320 9404
rect 2372 9392 2378 9444
rect 2424 9376 2452 9472
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 5123 9472 5273 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5261 9469 5273 9472
rect 5307 9469 5319 9503
rect 8720 9503 8778 9509
rect 8720 9500 8732 9503
rect 5261 9463 5319 9469
rect 8036 9472 8732 9500
rect 2406 9364 2412 9376
rect 2367 9336 2412 9364
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 3234 9364 3240 9376
rect 3195 9336 3240 9364
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 5276 9364 5304 9463
rect 6454 9392 6460 9444
rect 6512 9432 6518 9444
rect 6917 9435 6975 9441
rect 6917 9432 6929 9435
rect 6512 9404 6929 9432
rect 6512 9392 6518 9404
rect 6917 9401 6929 9404
rect 6963 9401 6975 9435
rect 6917 9395 6975 9401
rect 7009 9435 7067 9441
rect 7009 9401 7021 9435
rect 7055 9401 7067 9435
rect 7009 9395 7067 9401
rect 6822 9364 6828 9376
rect 5276 9336 6828 9364
rect 6822 9324 6828 9336
rect 6880 9364 6886 9376
rect 7024 9364 7052 9395
rect 8036 9376 8064 9472
rect 8720 9469 8732 9472
rect 8766 9500 8778 9503
rect 9398 9500 9404 9512
rect 8766 9472 9404 9500
rect 8766 9469 8778 9472
rect 8720 9463 8778 9469
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 11241 9503 11299 9509
rect 11241 9469 11253 9503
rect 11287 9469 11299 9503
rect 11241 9463 11299 9469
rect 8573 9435 8631 9441
rect 8573 9401 8585 9435
rect 8619 9432 8631 9435
rect 9030 9432 9036 9444
rect 8619 9404 9036 9432
rect 8619 9401 8631 9404
rect 8573 9395 8631 9401
rect 9030 9392 9036 9404
rect 9088 9392 9094 9444
rect 10642 9435 10700 9441
rect 10642 9432 10654 9435
rect 10152 9404 10654 9432
rect 8018 9364 8024 9376
rect 6880 9336 7052 9364
rect 7979 9336 8024 9364
rect 6880 9324 6886 9336
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 8386 9364 8392 9376
rect 8347 9336 8392 9364
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 10152 9373 10180 9404
rect 10642 9401 10654 9404
rect 10688 9432 10700 9435
rect 11146 9432 11152 9444
rect 10688 9404 11152 9432
rect 10688 9401 10700 9404
rect 10642 9395 10700 9401
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 11256 9432 11284 9463
rect 12250 9460 12256 9512
rect 12308 9500 12314 9512
rect 12452 9509 12480 9540
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12308 9472 12449 9500
rect 12308 9460 12314 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12986 9500 12992 9512
rect 12947 9472 12992 9500
rect 12437 9463 12495 9469
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13786 9472 13921 9500
rect 11606 9432 11612 9444
rect 11256 9404 11612 9432
rect 11606 9392 11612 9404
rect 11664 9432 11670 9444
rect 13786 9432 13814 9472
rect 13909 9469 13921 9472
rect 13955 9500 13967 9503
rect 14093 9503 14151 9509
rect 14093 9500 14105 9503
rect 13955 9472 14105 9500
rect 13955 9469 13967 9472
rect 13909 9463 13967 9469
rect 14093 9469 14105 9472
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 16644 9503 16702 9509
rect 16644 9469 16656 9503
rect 16690 9500 16702 9503
rect 17034 9500 17040 9512
rect 16690 9472 17040 9500
rect 16690 9469 16702 9472
rect 16644 9463 16702 9469
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 13998 9432 14004 9444
rect 11664 9404 13814 9432
rect 13959 9404 14004 9432
rect 11664 9392 11670 9404
rect 13998 9392 14004 9404
rect 14056 9392 14062 9444
rect 10137 9367 10195 9373
rect 10137 9364 10149 9367
rect 10100 9336 10149 9364
rect 10100 9324 10106 9336
rect 10137 9333 10149 9336
rect 10183 9333 10195 9367
rect 12526 9364 12532 9376
rect 12487 9336 12532 9364
rect 10137 9327 10195 9333
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 16715 9367 16773 9373
rect 16715 9333 16727 9367
rect 16761 9364 16773 9367
rect 18046 9364 18052 9376
rect 16761 9336 18052 9364
rect 16761 9333 16773 9336
rect 16715 9327 16773 9333
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 3510 9160 3516 9172
rect 3471 9132 3516 9160
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 4065 9163 4123 9169
rect 4065 9129 4077 9163
rect 4111 9160 4123 9163
rect 4430 9160 4436 9172
rect 4111 9132 4436 9160
rect 4111 9129 4123 9132
rect 4065 9123 4123 9129
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 4522 9120 4528 9172
rect 4580 9160 4586 9172
rect 6454 9160 6460 9172
rect 4580 9132 6460 9160
rect 4580 9120 4586 9132
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 6822 9160 6828 9172
rect 6783 9132 6828 9160
rect 6822 9120 6828 9132
rect 6880 9160 6886 9172
rect 7929 9163 7987 9169
rect 7929 9160 7941 9163
rect 6880 9132 7941 9160
rect 6880 9120 6886 9132
rect 7929 9129 7941 9132
rect 7975 9129 7987 9163
rect 8294 9160 8300 9172
rect 8255 9132 8300 9160
rect 7929 9123 7987 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 9030 9160 9036 9172
rect 8991 9132 9036 9160
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10321 9163 10379 9169
rect 10321 9160 10333 9163
rect 10192 9132 10333 9160
rect 10192 9120 10198 9132
rect 10321 9129 10333 9132
rect 10367 9129 10379 9163
rect 10686 9160 10692 9172
rect 10647 9132 10692 9160
rect 10321 9123 10379 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11514 9120 11520 9172
rect 11572 9160 11578 9172
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 11572 9132 12081 9160
rect 11572 9120 11578 9132
rect 12069 9129 12081 9132
rect 12115 9129 12127 9163
rect 12710 9160 12716 9172
rect 12671 9132 12716 9160
rect 12069 9123 12127 9129
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 1946 9092 1952 9104
rect 1907 9064 1952 9092
rect 1946 9052 1952 9064
rect 2004 9052 2010 9104
rect 4890 9052 4896 9104
rect 4948 9092 4954 9104
rect 4948 9064 5948 9092
rect 4948 9052 4954 9064
rect 5258 9024 5264 9036
rect 4126 8996 5264 9024
rect 1854 8956 1860 8968
rect 1815 8928 1860 8956
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 2498 8956 2504 8968
rect 2459 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2774 8956 2780 8968
rect 2735 8928 2780 8956
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 2130 8848 2136 8900
rect 2188 8888 2194 8900
rect 4126 8888 4154 8996
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 5920 9033 5948 9064
rect 6178 9052 6184 9104
rect 6236 9092 6242 9104
rect 6638 9092 6644 9104
rect 6236 9064 6644 9092
rect 6236 9052 6242 9064
rect 6638 9052 6644 9064
rect 6696 9092 6702 9104
rect 7330 9095 7388 9101
rect 7330 9092 7342 9095
rect 6696 9064 7342 9092
rect 6696 9052 6702 9064
rect 7330 9061 7342 9064
rect 7376 9061 7388 9095
rect 11238 9092 11244 9104
rect 11199 9064 11244 9092
rect 7330 9055 7388 9061
rect 11238 9052 11244 9064
rect 11296 9052 11302 9104
rect 14921 9095 14979 9101
rect 14921 9061 14933 9095
rect 14967 9092 14979 9095
rect 15470 9092 15476 9104
rect 14967 9064 15476 9092
rect 14967 9061 14979 9064
rect 14921 9055 14979 9061
rect 15470 9052 15476 9064
rect 15528 9052 15534 9104
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 8993 5595 9027
rect 5537 8987 5595 8993
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 5350 8956 5356 8968
rect 2188 8860 4154 8888
rect 4908 8928 5356 8956
rect 2188 8848 2194 8860
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 2038 8780 2044 8832
rect 2096 8820 2102 8832
rect 3145 8823 3203 8829
rect 3145 8820 3157 8823
rect 2096 8792 3157 8820
rect 2096 8780 2102 8792
rect 3145 8789 3157 8792
rect 3191 8820 3203 8823
rect 3234 8820 3240 8832
rect 3191 8792 3240 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 4908 8829 4936 8928
rect 5350 8916 5356 8928
rect 5408 8956 5414 8968
rect 5552 8956 5580 8987
rect 11882 8984 11888 9036
rect 11940 9024 11946 9036
rect 12894 9024 12900 9036
rect 11940 8996 12900 9024
rect 11940 8984 11946 8996
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 12986 8984 12992 9036
rect 13044 9024 13050 9036
rect 13081 9027 13139 9033
rect 13081 9024 13093 9027
rect 13044 8996 13093 9024
rect 13044 8984 13050 8996
rect 13081 8993 13093 8996
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 13170 8984 13176 9036
rect 13228 9024 13234 9036
rect 13630 9024 13636 9036
rect 13228 8996 13636 9024
rect 13228 8984 13234 8996
rect 13630 8984 13636 8996
rect 13688 9024 13694 9036
rect 15289 9027 15347 9033
rect 13688 8996 15240 9024
rect 13688 8984 13694 8996
rect 5408 8928 5580 8956
rect 6181 8959 6239 8965
rect 5408 8916 5414 8928
rect 6181 8925 6193 8959
rect 6227 8956 6239 8959
rect 7009 8959 7067 8965
rect 7009 8956 7021 8959
rect 6227 8928 7021 8956
rect 6227 8925 6239 8928
rect 6181 8919 6239 8925
rect 7009 8925 7021 8928
rect 7055 8956 7067 8959
rect 7466 8956 7472 8968
rect 7055 8928 7472 8956
rect 7055 8925 7067 8928
rect 7009 8919 7067 8925
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8956 9919 8959
rect 10870 8956 10876 8968
rect 9907 8928 10876 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11974 8956 11980 8968
rect 11195 8928 11980 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 11974 8916 11980 8928
rect 12032 8956 12038 8968
rect 14185 8959 14243 8965
rect 14185 8956 14197 8959
rect 12032 8928 14197 8956
rect 12032 8916 12038 8928
rect 14185 8925 14197 8928
rect 14231 8925 14243 8959
rect 15212 8956 15240 8996
rect 15289 8993 15301 9027
rect 15335 9024 15347 9027
rect 15378 9024 15384 9036
rect 15335 8996 15384 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 15378 8984 15384 8996
rect 15436 9024 15442 9036
rect 16850 9024 16856 9036
rect 15436 8996 16856 9024
rect 15436 8984 15442 8996
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 15657 8959 15715 8965
rect 15657 8956 15669 8959
rect 15212 8928 15669 8956
rect 14185 8919 14243 8925
rect 15657 8925 15669 8928
rect 15703 8956 15715 8959
rect 16206 8956 16212 8968
rect 15703 8928 16212 8956
rect 15703 8925 15715 8928
rect 15657 8919 15715 8925
rect 16206 8916 16212 8928
rect 16264 8916 16270 8968
rect 11701 8891 11759 8897
rect 11701 8857 11713 8891
rect 11747 8888 11759 8891
rect 11790 8888 11796 8900
rect 11747 8860 11796 8888
rect 11747 8857 11759 8860
rect 11701 8851 11759 8857
rect 11790 8848 11796 8860
rect 11848 8848 11854 8900
rect 15565 8891 15623 8897
rect 15565 8857 15577 8891
rect 15611 8888 15623 8891
rect 15838 8888 15844 8900
rect 15611 8860 15844 8888
rect 15611 8857 15623 8860
rect 15565 8851 15623 8857
rect 15838 8848 15844 8860
rect 15896 8848 15902 8900
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4488 8792 4905 8820
rect 4488 8780 4494 8792
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 8570 8820 8576 8832
rect 8531 8792 8576 8820
rect 4893 8783 4951 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 10134 8780 10140 8832
rect 10192 8820 10198 8832
rect 12437 8823 12495 8829
rect 12437 8820 12449 8823
rect 10192 8792 12449 8820
rect 10192 8780 10198 8792
rect 12437 8789 12449 8792
rect 12483 8820 12495 8823
rect 12986 8820 12992 8832
rect 12483 8792 12992 8820
rect 12483 8789 12495 8792
rect 12437 8783 12495 8789
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 14826 8780 14832 8832
rect 14884 8820 14890 8832
rect 15427 8823 15485 8829
rect 15427 8820 15439 8823
rect 14884 8792 15439 8820
rect 14884 8780 14890 8792
rect 15427 8789 15439 8792
rect 15473 8789 15485 8823
rect 15746 8820 15752 8832
rect 15707 8792 15752 8820
rect 15427 8783 15485 8789
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2222 8576 2228 8628
rect 2280 8616 2286 8628
rect 4890 8616 4896 8628
rect 2280 8588 4896 8616
rect 2280 8576 2286 8588
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5316 8588 6009 8616
rect 5316 8576 5322 8588
rect 5997 8585 6009 8588
rect 6043 8585 6055 8619
rect 5997 8579 6055 8585
rect 8389 8619 8447 8625
rect 8389 8585 8401 8619
rect 8435 8616 8447 8619
rect 8478 8616 8484 8628
rect 8435 8588 8484 8616
rect 8435 8585 8447 8588
rect 8389 8579 8447 8585
rect 8478 8576 8484 8588
rect 8536 8616 8542 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 8536 8588 9321 8616
rect 8536 8576 8542 8588
rect 9309 8585 9321 8588
rect 9355 8616 9367 8619
rect 10134 8616 10140 8628
rect 9355 8588 9904 8616
rect 10095 8588 10140 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 2498 8548 2504 8560
rect 2459 8520 2504 8548
rect 2498 8508 2504 8520
rect 2556 8508 2562 8560
rect 4525 8551 4583 8557
rect 4525 8517 4537 8551
rect 4571 8548 4583 8551
rect 5442 8548 5448 8560
rect 4571 8520 5448 8548
rect 4571 8517 4583 8520
rect 4525 8511 4583 8517
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 9033 8551 9091 8557
rect 9033 8548 9045 8551
rect 8352 8520 9045 8548
rect 8352 8508 8358 8520
rect 9033 8517 9045 8520
rect 9079 8548 9091 8551
rect 9766 8548 9772 8560
rect 9079 8520 9772 8548
rect 9079 8517 9091 8520
rect 9033 8511 9091 8517
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 1946 8480 1952 8492
rect 1811 8452 1952 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 1946 8440 1952 8452
rect 2004 8480 2010 8492
rect 9876 8489 9904 8588
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 11609 8619 11667 8625
rect 11609 8616 11621 8619
rect 11296 8588 11621 8616
rect 11296 8576 11302 8588
rect 11609 8585 11621 8588
rect 11655 8585 11667 8619
rect 11974 8616 11980 8628
rect 11935 8588 11980 8616
rect 11609 8579 11667 8585
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 12986 8616 12992 8628
rect 12947 8588 12992 8616
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 14642 8616 14648 8628
rect 14603 8588 14648 8616
rect 14642 8576 14648 8588
rect 14700 8576 14706 8628
rect 16206 8616 16212 8628
rect 16167 8588 16212 8616
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16482 8576 16488 8628
rect 16540 8616 16546 8628
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 16540 8588 16681 8616
rect 16540 8576 16546 8588
rect 16669 8585 16681 8588
rect 16715 8585 16727 8619
rect 16669 8579 16727 8585
rect 11514 8508 11520 8560
rect 11572 8548 11578 8560
rect 11572 8520 16471 8548
rect 11572 8508 11578 8520
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 2004 8452 3433 8480
rect 2004 8440 2010 8452
rect 3421 8449 3433 8452
rect 3467 8449 3479 8483
rect 3421 8443 3479 8449
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 9640 8483 9698 8489
rect 9640 8480 9652 8483
rect 4387 8452 9652 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 9640 8449 9652 8452
rect 9686 8480 9698 8483
rect 9861 8483 9919 8489
rect 9686 8452 9812 8480
rect 9686 8449 9698 8452
rect 9640 8443 9698 8449
rect 2682 8372 2688 8424
rect 2740 8412 2746 8424
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2740 8384 2973 8412
rect 2740 8372 2746 8384
rect 2961 8381 2973 8384
rect 3007 8412 3019 8415
rect 3329 8415 3387 8421
rect 3329 8412 3341 8415
rect 3007 8384 3341 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 3329 8381 3341 8384
rect 3375 8412 3387 8415
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 3375 8384 3525 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3513 8381 3525 8384
rect 3559 8381 3571 8415
rect 3513 8375 3571 8381
rect 5261 8415 5319 8421
rect 5261 8381 5273 8415
rect 5307 8412 5319 8415
rect 5442 8412 5448 8424
rect 5307 8384 5448 8412
rect 5307 8381 5319 8384
rect 5261 8375 5319 8381
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8412 5595 8415
rect 5810 8412 5816 8424
rect 5583 8384 5816 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 5810 8372 5816 8384
rect 5868 8372 5874 8424
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 6860 8415 6918 8421
rect 6860 8412 6872 8415
rect 6788 8384 6872 8412
rect 6788 8372 6794 8384
rect 6860 8381 6872 8384
rect 6906 8412 6918 8415
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 6906 8384 7297 8412
rect 6906 8381 6918 8384
rect 6860 8375 6918 8381
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 1946 8344 1952 8356
rect 1907 8316 1952 8344
rect 1946 8304 1952 8316
rect 2004 8304 2010 8356
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8313 2099 8347
rect 2041 8307 2099 8313
rect 2056 8276 2084 8307
rect 4614 8304 4620 8356
rect 4672 8344 4678 8356
rect 6963 8347 7021 8353
rect 6963 8344 6975 8347
rect 4672 8316 6975 8344
rect 4672 8304 4678 8316
rect 6963 8313 6975 8316
rect 7009 8313 7021 8347
rect 6963 8307 7021 8313
rect 2682 8276 2688 8288
rect 2056 8248 2688 8276
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 4341 8279 4399 8285
rect 4341 8276 4353 8279
rect 3936 8248 4353 8276
rect 3936 8236 3942 8248
rect 4341 8245 4353 8248
rect 4387 8245 4399 8279
rect 5074 8276 5080 8288
rect 5035 8248 5080 8276
rect 4341 8239 4399 8245
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 6236 8248 6561 8276
rect 6236 8236 6242 8248
rect 6549 8245 6561 8248
rect 6595 8245 6607 8279
rect 6549 8239 6607 8245
rect 7837 8279 7895 8285
rect 7837 8245 7849 8279
rect 7883 8276 7895 8279
rect 8036 8276 8064 8375
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 8720 8384 9505 8412
rect 8720 8372 8726 8384
rect 9493 8381 9505 8384
rect 9539 8381 9551 8415
rect 9784 8412 9812 8452
rect 9861 8449 9873 8483
rect 9907 8480 9919 8483
rect 13170 8480 13176 8492
rect 9907 8452 13176 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 13722 8480 13728 8492
rect 13683 8452 13728 8480
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 10873 8415 10931 8421
rect 10873 8412 10885 8415
rect 9784 8384 10885 8412
rect 9493 8375 9551 8381
rect 10873 8381 10885 8384
rect 10919 8412 10931 8415
rect 10962 8412 10968 8424
rect 10919 8384 10968 8412
rect 10919 8381 10931 8384
rect 10873 8375 10931 8381
rect 9508 8344 9536 8375
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 11146 8421 11152 8424
rect 11124 8415 11152 8421
rect 11124 8412 11136 8415
rect 11059 8384 11136 8412
rect 11124 8381 11136 8384
rect 11204 8412 11210 8424
rect 11790 8412 11796 8424
rect 11204 8384 11796 8412
rect 11124 8375 11152 8381
rect 11146 8372 11152 8375
rect 11204 8372 11210 8384
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 14642 8372 14648 8424
rect 14700 8412 14706 8424
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 14700 8384 14841 8412
rect 14700 8372 14706 8384
rect 14829 8381 14841 8384
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 15381 8415 15439 8421
rect 15381 8381 15393 8415
rect 15427 8412 15439 8415
rect 15470 8412 15476 8424
rect 15427 8384 15476 8412
rect 15427 8381 15439 8384
rect 15381 8375 15439 8381
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 16443 8421 16471 8520
rect 16428 8415 16486 8421
rect 16428 8381 16440 8415
rect 16474 8412 16486 8415
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 16474 8384 17233 8412
rect 16474 8381 16486 8384
rect 16428 8375 16486 8381
rect 17221 8381 17233 8384
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 10505 8347 10563 8353
rect 10505 8344 10517 8347
rect 9508 8316 10517 8344
rect 10505 8313 10517 8316
rect 10551 8313 10563 8347
rect 10505 8307 10563 8313
rect 13357 8347 13415 8353
rect 13357 8313 13369 8347
rect 13403 8313 13415 8347
rect 13357 8307 13415 8313
rect 8570 8276 8576 8288
rect 7883 8248 8576 8276
rect 7883 8245 7895 8248
rect 7837 8239 7895 8245
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11195 8279 11253 8285
rect 11195 8276 11207 8279
rect 11112 8248 11207 8276
rect 11112 8236 11118 8248
rect 11195 8245 11207 8248
rect 11241 8245 11253 8279
rect 11195 8239 11253 8245
rect 12713 8279 12771 8285
rect 12713 8245 12725 8279
rect 12759 8276 12771 8279
rect 12894 8276 12900 8288
rect 12759 8248 12900 8276
rect 12759 8245 12771 8248
rect 12713 8239 12771 8245
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 13372 8276 13400 8307
rect 13446 8304 13452 8356
rect 13504 8344 13510 8356
rect 22094 8344 22100 8356
rect 13504 8316 13549 8344
rect 13786 8316 22100 8344
rect 13504 8304 13510 8316
rect 13786 8288 13814 8316
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 13786 8276 13820 8288
rect 13372 8248 13820 8276
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 14734 8236 14740 8288
rect 14792 8276 14798 8288
rect 14921 8279 14979 8285
rect 14921 8276 14933 8279
rect 14792 8248 14933 8276
rect 14792 8236 14798 8248
rect 14921 8245 14933 8248
rect 14967 8245 14979 8279
rect 15838 8276 15844 8288
rect 15799 8248 15844 8276
rect 14921 8239 14979 8245
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 16850 8276 16856 8288
rect 16811 8248 16856 8276
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 2096 8044 2145 8072
rect 2096 8032 2102 8044
rect 2133 8041 2145 8044
rect 2179 8041 2191 8075
rect 2682 8072 2688 8084
rect 2643 8044 2688 8072
rect 2133 8035 2191 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 3050 8072 3056 8084
rect 2963 8044 3056 8072
rect 3050 8032 3056 8044
rect 3108 8072 3114 8084
rect 5074 8072 5080 8084
rect 3108 8044 5080 8072
rect 3108 8032 3114 8044
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 7466 8072 7472 8084
rect 7427 8044 7472 8072
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 11146 8072 11152 8084
rect 11107 8044 11152 8072
rect 11146 8032 11152 8044
rect 11204 8032 11210 8084
rect 12250 8032 12256 8084
rect 12308 8072 12314 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 12308 8044 12357 8072
rect 12308 8032 12314 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12345 8035 12403 8041
rect 13725 8075 13783 8081
rect 13725 8041 13737 8075
rect 13771 8072 13783 8075
rect 13814 8072 13820 8084
rect 13771 8044 13820 8072
rect 13771 8041 13783 8044
rect 13725 8035 13783 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 15378 8072 15384 8084
rect 15339 8044 15384 8072
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 8021 8007 8079 8013
rect 8021 7973 8033 8007
rect 8067 8004 8079 8007
rect 8662 8004 8668 8016
rect 8067 7976 8668 8004
rect 8067 7973 8079 7976
rect 8021 7967 8079 7973
rect 8662 7964 8668 7976
rect 8720 7964 8726 8016
rect 1946 7896 1952 7948
rect 2004 7936 2010 7948
rect 3329 7939 3387 7945
rect 3329 7936 3341 7939
rect 2004 7908 3341 7936
rect 2004 7896 2010 7908
rect 3329 7905 3341 7908
rect 3375 7936 3387 7939
rect 4614 7936 4620 7948
rect 3375 7908 4620 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 5350 7936 5356 7948
rect 5311 7908 5356 7936
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5810 7936 5816 7948
rect 5771 7908 5816 7936
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6546 7936 6552 7948
rect 6507 7908 6552 7936
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 9858 7936 9864 7948
rect 9819 7908 9864 7936
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 11974 7936 11980 7948
rect 11887 7908 11980 7936
rect 11974 7896 11980 7908
rect 12032 7936 12038 7948
rect 12526 7936 12532 7948
rect 12032 7908 12532 7936
rect 12032 7896 12038 7908
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 15286 7936 15292 7948
rect 15247 7908 15292 7936
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15470 7896 15476 7948
rect 15528 7936 15534 7948
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 15528 7908 15853 7936
rect 15528 7896 15534 7908
rect 15841 7905 15853 7908
rect 15887 7936 15899 7939
rect 17494 7936 17500 7948
rect 15887 7908 17500 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 17494 7896 17500 7908
rect 17552 7896 17558 7948
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 1688 7840 1777 7868
rect 1688 7744 1716 7840
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 4706 7868 4712 7880
rect 4667 7840 4712 7868
rect 1765 7831 1823 7837
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7868 8447 7871
rect 8570 7868 8576 7880
rect 8435 7840 8576 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 7208 7800 7236 7831
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 10502 7868 10508 7880
rect 10463 7840 10508 7868
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 13906 7868 13912 7880
rect 13867 7840 13912 7868
rect 13906 7828 13912 7840
rect 13964 7828 13970 7880
rect 8294 7800 8300 7812
rect 7208 7772 8300 7800
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 1854 7692 1860 7744
rect 1912 7732 1918 7744
rect 3697 7735 3755 7741
rect 3697 7732 3709 7735
rect 1912 7704 3709 7732
rect 1912 7692 1918 7704
rect 3697 7701 3709 7704
rect 3743 7701 3755 7735
rect 3697 7695 3755 7701
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 8018 7732 8024 7744
rect 7156 7704 8024 7732
rect 7156 7692 7162 7704
rect 8018 7692 8024 7704
rect 8076 7732 8082 7744
rect 8159 7735 8217 7741
rect 8159 7732 8171 7735
rect 8076 7704 8171 7732
rect 8076 7692 8082 7704
rect 8159 7701 8171 7704
rect 8205 7701 8217 7735
rect 8478 7732 8484 7744
rect 8439 7704 8484 7732
rect 8159 7695 8217 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 12897 7735 12955 7741
rect 12897 7732 12909 7735
rect 11940 7704 12909 7732
rect 11940 7692 11946 7704
rect 12897 7701 12909 7704
rect 12943 7732 12955 7735
rect 13265 7735 13323 7741
rect 13265 7732 13277 7735
rect 12943 7704 13277 7732
rect 12943 7701 12955 7704
rect 12897 7695 12955 7701
rect 13265 7701 13277 7704
rect 13311 7732 13323 7735
rect 13446 7732 13452 7744
rect 13311 7704 13452 7732
rect 13311 7701 13323 7704
rect 13265 7695 13323 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 15013 7735 15071 7741
rect 15013 7732 15025 7735
rect 14884 7704 15025 7732
rect 14884 7692 14890 7704
rect 15013 7701 15025 7704
rect 15059 7701 15071 7735
rect 15013 7695 15071 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 3418 7488 3424 7540
rect 3476 7528 3482 7540
rect 4065 7531 4123 7537
rect 4065 7528 4077 7531
rect 3476 7500 4077 7528
rect 3476 7488 3482 7500
rect 4065 7497 4077 7500
rect 4111 7528 4123 7531
rect 4111 7500 5120 7528
rect 4111 7497 4123 7500
rect 4065 7491 4123 7497
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7392 2743 7395
rect 3050 7392 3056 7404
rect 2731 7364 3056 7392
rect 2731 7361 2743 7364
rect 2685 7355 2743 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 5092 7401 5120 7500
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 10597 7531 10655 7537
rect 10597 7528 10609 7531
rect 10560 7500 10609 7528
rect 10560 7488 10566 7500
rect 10597 7497 10609 7500
rect 10643 7528 10655 7531
rect 10962 7528 10968 7540
rect 10643 7500 10968 7528
rect 10643 7497 10655 7500
rect 10597 7491 10655 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 13725 7531 13783 7537
rect 13725 7497 13737 7531
rect 13771 7528 13783 7531
rect 13906 7528 13912 7540
rect 13771 7500 13912 7528
rect 13771 7497 13783 7500
rect 13725 7491 13783 7497
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 11793 7463 11851 7469
rect 11793 7460 11805 7463
rect 10060 7432 11805 7460
rect 10060 7404 10088 7432
rect 11793 7429 11805 7432
rect 11839 7460 11851 7463
rect 12161 7463 12219 7469
rect 12161 7460 12173 7463
rect 11839 7432 12173 7460
rect 11839 7429 11851 7432
rect 11793 7423 11851 7429
rect 12161 7429 12173 7432
rect 12207 7460 12219 7463
rect 12250 7460 12256 7472
rect 12207 7432 12256 7460
rect 12207 7429 12219 7432
rect 12161 7423 12219 7429
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5534 7392 5540 7404
rect 5495 7364 5540 7392
rect 5077 7355 5135 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 10042 7392 10048 7404
rect 9646 7364 10048 7392
rect 106 7284 112 7336
rect 164 7324 170 7336
rect 1432 7327 1490 7333
rect 1432 7324 1444 7327
rect 164 7296 1444 7324
rect 164 7284 170 7296
rect 1432 7293 1444 7296
rect 1478 7324 1490 7327
rect 1857 7327 1915 7333
rect 1857 7324 1869 7327
rect 1478 7296 1869 7324
rect 1478 7293 1490 7296
rect 1432 7287 1490 7293
rect 1857 7293 1869 7296
rect 1903 7293 1915 7327
rect 7742 7324 7748 7336
rect 7703 7296 7748 7324
rect 1857 7287 1915 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 9033 7327 9091 7333
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9122 7324 9128 7336
rect 9079 7296 9128 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 1535 7259 1593 7265
rect 1535 7225 1547 7259
rect 1581 7256 1593 7259
rect 2866 7256 2872 7268
rect 1581 7228 2872 7256
rect 1581 7225 1593 7228
rect 1535 7219 1593 7225
rect 2866 7216 2872 7228
rect 2924 7216 2930 7268
rect 3006 7259 3064 7265
rect 3006 7225 3018 7259
rect 3052 7225 3064 7259
rect 3006 7219 3064 7225
rect 4525 7259 4583 7265
rect 4525 7225 4537 7259
rect 4571 7256 4583 7259
rect 4893 7259 4951 7265
rect 4893 7256 4905 7259
rect 4571 7228 4905 7256
rect 4571 7225 4583 7228
rect 4525 7219 4583 7225
rect 4893 7225 4905 7228
rect 4939 7256 4951 7259
rect 5169 7259 5227 7265
rect 5169 7256 5181 7259
rect 4939 7228 5181 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 5169 7225 5181 7228
rect 5215 7256 5227 7259
rect 5350 7256 5356 7268
rect 5215 7228 5356 7256
rect 5215 7225 5227 7228
rect 5169 7219 5227 7225
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 2501 7191 2559 7197
rect 2501 7188 2513 7191
rect 2096 7160 2513 7188
rect 2096 7148 2102 7160
rect 2501 7157 2513 7160
rect 2547 7188 2559 7191
rect 3021 7188 3049 7219
rect 5350 7216 5356 7228
rect 5408 7216 5414 7268
rect 8205 7259 8263 7265
rect 8205 7225 8217 7259
rect 8251 7256 8263 7259
rect 9214 7256 9220 7268
rect 8251 7228 9220 7256
rect 8251 7225 8263 7228
rect 8205 7219 8263 7225
rect 9214 7216 9220 7228
rect 9272 7216 9278 7268
rect 9395 7259 9453 7265
rect 9395 7225 9407 7259
rect 9441 7256 9453 7259
rect 9646 7256 9674 7364
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 10870 7392 10876 7404
rect 10831 7364 10876 7392
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 11514 7392 11520 7404
rect 11475 7364 11520 7392
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7392 12495 7395
rect 12710 7392 12716 7404
rect 12483 7364 12716 7392
rect 12483 7361 12495 7364
rect 12437 7355 12495 7361
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 13924 7392 13952 7488
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13924 7364 14289 7392
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14550 7392 14556 7404
rect 14511 7364 14556 7392
rect 14277 7355 14335 7361
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 16025 7327 16083 7333
rect 16025 7293 16037 7327
rect 16071 7293 16083 7327
rect 16298 7324 16304 7336
rect 16259 7296 16304 7324
rect 16025 7287 16083 7293
rect 9441 7228 9674 7256
rect 9441 7225 9453 7228
rect 9395 7219 9453 7225
rect 3602 7188 3608 7200
rect 2547 7160 3049 7188
rect 3563 7160 3608 7188
rect 2547 7157 2559 7160
rect 2501 7151 2559 7157
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 6546 7188 6552 7200
rect 6507 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 7098 7148 7104 7200
rect 7156 7188 7162 7200
rect 7285 7191 7343 7197
rect 7285 7188 7297 7191
rect 7156 7160 7297 7188
rect 7156 7148 7162 7160
rect 7285 7157 7297 7160
rect 7331 7157 7343 7191
rect 8570 7188 8576 7200
rect 8531 7160 8576 7188
rect 7285 7151 7343 7157
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 8846 7188 8852 7200
rect 8807 7160 8852 7188
rect 8846 7148 8852 7160
rect 8904 7188 8910 7200
rect 9416 7188 9444 7219
rect 10962 7216 10968 7268
rect 11020 7256 11026 7268
rect 11020 7228 11065 7256
rect 11020 7216 11026 7228
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 12758 7259 12816 7265
rect 12758 7256 12770 7259
rect 12308 7228 12770 7256
rect 12308 7216 12314 7228
rect 12758 7225 12770 7228
rect 12804 7225 12816 7259
rect 12758 7219 12816 7225
rect 14093 7259 14151 7265
rect 14093 7225 14105 7259
rect 14139 7256 14151 7259
rect 14366 7256 14372 7268
rect 14139 7228 14372 7256
rect 14139 7225 14151 7228
rect 14093 7219 14151 7225
rect 14366 7216 14372 7228
rect 14424 7216 14430 7268
rect 15286 7216 15292 7268
rect 15344 7256 15350 7268
rect 15381 7259 15439 7265
rect 15381 7256 15393 7259
rect 15344 7228 15393 7256
rect 15344 7216 15350 7228
rect 15381 7225 15393 7228
rect 15427 7256 15439 7259
rect 15562 7256 15568 7268
rect 15427 7228 15568 7256
rect 15427 7225 15439 7228
rect 15381 7219 15439 7225
rect 15562 7216 15568 7228
rect 15620 7256 15626 7268
rect 16040 7256 16068 7287
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 16761 7259 16819 7265
rect 16761 7256 16773 7259
rect 15620 7228 16773 7256
rect 15620 7216 15626 7228
rect 16761 7225 16773 7228
rect 16807 7225 16819 7259
rect 16761 7219 16819 7225
rect 8904 7160 9444 7188
rect 8904 7148 8910 7160
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9916 7160 9965 7188
rect 9916 7148 9922 7160
rect 9953 7157 9965 7160
rect 9999 7188 10011 7191
rect 10229 7191 10287 7197
rect 10229 7188 10241 7191
rect 9999 7160 10241 7188
rect 9999 7157 10011 7160
rect 9953 7151 10011 7157
rect 10229 7157 10241 7160
rect 10275 7157 10287 7191
rect 13354 7188 13360 7200
rect 13315 7160 13360 7188
rect 10229 7151 10287 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 15838 7188 15844 7200
rect 15799 7160 15844 7188
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2314 6984 2320 6996
rect 2275 6956 2320 6984
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 2498 6944 2504 6996
rect 2556 6984 2562 6996
rect 3234 6984 3240 6996
rect 2556 6956 3240 6984
rect 2556 6944 2562 6956
rect 3234 6944 3240 6956
rect 3292 6984 3298 6996
rect 3421 6987 3479 6993
rect 3421 6984 3433 6987
rect 3292 6956 3433 6984
rect 3292 6944 3298 6956
rect 3421 6953 3433 6956
rect 3467 6953 3479 6987
rect 3421 6947 3479 6953
rect 5350 6944 5356 6996
rect 5408 6984 5414 6996
rect 5813 6987 5871 6993
rect 5813 6984 5825 6987
rect 5408 6956 5825 6984
rect 5408 6944 5414 6956
rect 5813 6953 5825 6956
rect 5859 6953 5871 6987
rect 5813 6947 5871 6953
rect 8113 6987 8171 6993
rect 8113 6953 8125 6987
rect 8159 6984 8171 6987
rect 8294 6984 8300 6996
rect 8159 6956 8300 6984
rect 8159 6953 8171 6956
rect 8113 6947 8171 6953
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 8481 6987 8539 6993
rect 8481 6953 8493 6987
rect 8527 6984 8539 6987
rect 8662 6984 8668 6996
rect 8527 6956 8668 6984
rect 8527 6953 8539 6956
rect 8481 6947 8539 6953
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 10870 6984 10876 6996
rect 10831 6956 10876 6984
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 11974 6984 11980 6996
rect 11935 6956 11980 6984
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 13081 6987 13139 6993
rect 13081 6984 13093 6987
rect 12768 6956 13093 6984
rect 12768 6944 12774 6956
rect 13081 6953 13093 6956
rect 13127 6953 13139 6987
rect 13081 6947 13139 6953
rect 14737 6987 14795 6993
rect 14737 6953 14749 6987
rect 14783 6984 14795 6987
rect 15470 6984 15476 6996
rect 14783 6956 15476 6984
rect 14783 6953 14795 6956
rect 14737 6947 14795 6953
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 17494 6984 17500 6996
rect 17455 6956 17500 6984
rect 17494 6944 17500 6956
rect 17552 6944 17558 6996
rect 24719 6987 24777 6993
rect 24719 6953 24731 6987
rect 24765 6984 24777 6987
rect 24854 6984 24860 6996
rect 24765 6956 24860 6984
rect 24765 6953 24777 6956
rect 24719 6947 24777 6953
rect 24854 6944 24860 6956
rect 24912 6944 24918 6996
rect 2590 6916 2596 6928
rect 2551 6888 2596 6916
rect 2590 6876 2596 6888
rect 2648 6876 2654 6928
rect 2866 6876 2872 6928
rect 2924 6916 2930 6928
rect 4709 6919 4767 6925
rect 4709 6916 4721 6919
rect 2924 6888 4721 6916
rect 2924 6876 2930 6888
rect 4709 6885 4721 6888
rect 4755 6916 4767 6919
rect 4798 6916 4804 6928
rect 4755 6888 4804 6916
rect 4755 6885 4767 6888
rect 4709 6879 4767 6885
rect 4798 6876 4804 6888
rect 4856 6876 4862 6928
rect 5255 6919 5313 6925
rect 5255 6885 5267 6919
rect 5301 6916 5313 6919
rect 6178 6916 6184 6928
rect 5301 6888 6184 6916
rect 5301 6885 5313 6888
rect 5255 6879 5313 6885
rect 6178 6876 6184 6888
rect 6236 6876 6242 6928
rect 6270 6876 6276 6928
rect 6328 6916 6334 6928
rect 6825 6919 6883 6925
rect 6825 6916 6837 6919
rect 6328 6888 6837 6916
rect 6328 6876 6334 6888
rect 6825 6885 6837 6888
rect 6871 6885 6883 6919
rect 9858 6916 9864 6928
rect 9819 6888 9864 6916
rect 6825 6879 6883 6885
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 10413 6919 10471 6925
rect 10413 6885 10425 6919
rect 10459 6916 10471 6919
rect 11514 6916 11520 6928
rect 10459 6888 11520 6916
rect 10459 6885 10471 6888
rect 10413 6879 10471 6885
rect 11514 6876 11520 6888
rect 11572 6876 11578 6928
rect 13354 6876 13360 6928
rect 13412 6916 13418 6928
rect 13817 6919 13875 6925
rect 13817 6916 13829 6919
rect 13412 6888 13829 6916
rect 13412 6876 13418 6888
rect 13817 6885 13829 6888
rect 13863 6885 13875 6919
rect 13817 6879 13875 6885
rect 14369 6919 14427 6925
rect 14369 6885 14381 6919
rect 14415 6916 14427 6919
rect 14550 6916 14556 6928
rect 14415 6888 14556 6916
rect 14415 6885 14427 6888
rect 14369 6879 14427 6885
rect 14550 6876 14556 6888
rect 14608 6876 14614 6928
rect 14826 6876 14832 6928
rect 14884 6916 14890 6928
rect 27614 6916 27620 6928
rect 14884 6888 17043 6916
rect 14884 6876 14890 6888
rect 9122 6848 9128 6860
rect 9083 6820 9128 6848
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 15451 6857 15479 6888
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 11940 6820 12173 6848
rect 11940 6808 11946 6820
rect 12161 6817 12173 6820
rect 12207 6817 12219 6851
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 12161 6811 12219 6817
rect 15028 6820 15301 6848
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6780 1455 6783
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 1443 6752 2513 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 2501 6749 2513 6752
rect 2547 6780 2559 6783
rect 2958 6780 2964 6792
rect 2547 6752 2964 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6780 3203 6783
rect 3510 6780 3516 6792
rect 3191 6752 3516 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 4890 6780 4896 6792
rect 4851 6752 4896 6780
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 6730 6780 6736 6792
rect 6691 6752 6736 6780
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6780 8631 6783
rect 9582 6780 9588 6792
rect 8619 6752 9588 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 13722 6780 13728 6792
rect 13683 6752 13728 6780
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 15028 6789 15056 6820
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15436 6851 15494 6857
rect 15436 6817 15448 6851
rect 15482 6817 15494 6851
rect 16850 6848 16856 6860
rect 16811 6820 16856 6848
rect 15436 6811 15494 6817
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 17015 6857 17043 6888
rect 24647 6888 27620 6916
rect 24647 6860 24675 6888
rect 27614 6876 27620 6888
rect 27672 6876 27678 6928
rect 17000 6851 17058 6857
rect 17000 6817 17012 6851
rect 17046 6848 17058 6851
rect 17310 6848 17316 6860
rect 17046 6820 17316 6848
rect 17046 6817 17058 6820
rect 17000 6811 17058 6817
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 24647 6857 24676 6860
rect 24632 6851 24676 6857
rect 24632 6848 24644 6851
rect 24583 6820 24644 6848
rect 24632 6817 24644 6820
rect 24632 6811 24676 6817
rect 24670 6808 24676 6811
rect 24728 6808 24734 6860
rect 15013 6783 15071 6789
rect 15013 6780 15025 6783
rect 14200 6752 15025 6780
rect 7282 6712 7288 6724
rect 7243 6684 7288 6712
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 14200 6712 14228 6752
rect 15013 6749 15025 6752
rect 15059 6749 15071 6783
rect 15013 6743 15071 6749
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6780 15715 6783
rect 17221 6783 17279 6789
rect 17221 6780 17233 6783
rect 15703 6752 17233 6780
rect 15703 6749 15715 6752
rect 15657 6743 15715 6749
rect 17221 6749 17233 6752
rect 17267 6749 17279 6783
rect 17221 6743 17279 6749
rect 8720 6684 14228 6712
rect 8720 6672 8726 6684
rect 15286 6672 15292 6724
rect 15344 6712 15350 6724
rect 15672 6712 15700 6743
rect 15344 6684 15700 6712
rect 15764 6684 17172 6712
rect 15344 6672 15350 6684
rect 15764 6656 15792 6684
rect 1949 6647 2007 6653
rect 1949 6613 1961 6647
rect 1995 6644 2007 6647
rect 2038 6644 2044 6656
rect 1995 6616 2044 6644
rect 1995 6613 2007 6616
rect 1949 6607 2007 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 7742 6644 7748 6656
rect 7703 6616 7748 6644
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 12342 6644 12348 6656
rect 12303 6616 12348 6644
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 13449 6647 13507 6653
rect 13449 6644 13461 6647
rect 12768 6616 13461 6644
rect 12768 6604 12774 6616
rect 13449 6613 13461 6616
rect 13495 6613 13507 6647
rect 13449 6607 13507 6613
rect 15565 6647 15623 6653
rect 15565 6613 15577 6647
rect 15611 6644 15623 6647
rect 15746 6644 15752 6656
rect 15611 6616 15752 6644
rect 15611 6613 15623 6616
rect 15565 6607 15623 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 15933 6647 15991 6653
rect 15933 6613 15945 6647
rect 15979 6644 15991 6647
rect 16298 6644 16304 6656
rect 15979 6616 16304 6644
rect 15979 6613 15991 6616
rect 15933 6607 15991 6613
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 17144 6653 17172 6684
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17218 6644 17224 6656
rect 17175 6616 17224 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2958 6440 2964 6452
rect 2919 6412 2964 6440
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 4617 6443 4675 6449
rect 4617 6409 4629 6443
rect 4663 6440 4675 6443
rect 4706 6440 4712 6452
rect 4663 6412 4712 6440
rect 4663 6409 4675 6412
rect 4617 6403 4675 6409
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 6270 6440 6276 6452
rect 6231 6412 6276 6440
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9769 6443 9827 6449
rect 9769 6440 9781 6443
rect 9272 6412 9781 6440
rect 9272 6400 9278 6412
rect 9769 6409 9781 6412
rect 9815 6440 9827 6443
rect 10134 6440 10140 6452
rect 9815 6412 10140 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11882 6440 11888 6452
rect 11843 6412 11888 6440
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12342 6440 12348 6452
rect 12299 6412 12348 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 13633 6443 13691 6449
rect 13633 6440 13645 6443
rect 13412 6412 13645 6440
rect 13412 6400 13418 6412
rect 13633 6409 13645 6412
rect 13679 6440 13691 6443
rect 13679 6412 14136 6440
rect 13679 6409 13691 6412
rect 13633 6403 13691 6409
rect 4249 6375 4307 6381
rect 4249 6341 4261 6375
rect 4295 6372 4307 6375
rect 4890 6372 4896 6384
rect 4295 6344 4896 6372
rect 4295 6341 4307 6344
rect 4249 6335 4307 6341
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 6178 6332 6184 6384
rect 6236 6372 6242 6384
rect 8021 6375 8079 6381
rect 8021 6372 8033 6375
rect 6236 6344 8033 6372
rect 6236 6332 6242 6344
rect 8021 6341 8033 6344
rect 8067 6341 8079 6375
rect 8021 6335 8079 6341
rect 2222 6304 2228 6316
rect 1872 6276 2228 6304
rect 1872 6245 1900 6276
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 3234 6304 3240 6316
rect 3195 6276 3240 6304
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 3510 6304 3516 6316
rect 3471 6276 3516 6304
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 4798 6304 4804 6316
rect 4759 6276 4804 6304
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6304 5503 6307
rect 5534 6304 5540 6316
rect 5491 6276 5540 6304
rect 5491 6273 5503 6276
rect 5445 6267 5503 6273
rect 5534 6264 5540 6276
rect 5592 6304 5598 6316
rect 6730 6304 6736 6316
rect 5592 6276 6736 6304
rect 5592 6264 5598 6276
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6205 1915 6239
rect 1857 6199 1915 6205
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6236 2191 6239
rect 2314 6236 2320 6248
rect 2179 6208 2320 6236
rect 2179 6205 2191 6208
rect 2133 6199 2191 6205
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 5460 6208 7021 6236
rect 3329 6171 3387 6177
rect 3329 6137 3341 6171
rect 3375 6168 3387 6171
rect 3602 6168 3608 6180
rect 3375 6140 3608 6168
rect 3375 6137 3387 6140
rect 3329 6131 3387 6137
rect 3602 6128 3608 6140
rect 3660 6128 3666 6180
rect 4798 6128 4804 6180
rect 4856 6168 4862 6180
rect 4893 6171 4951 6177
rect 4893 6168 4905 6171
rect 4856 6140 4905 6168
rect 4856 6128 4862 6140
rect 4893 6137 4905 6140
rect 4939 6137 4951 6171
rect 4893 6131 4951 6137
rect 1670 6100 1676 6112
rect 1631 6072 1676 6100
rect 1670 6060 1676 6072
rect 1728 6060 1734 6112
rect 2590 6060 2596 6112
rect 2648 6100 2654 6112
rect 2685 6103 2743 6109
rect 2685 6100 2697 6103
rect 2648 6072 2697 6100
rect 2648 6060 2654 6072
rect 2685 6069 2697 6072
rect 2731 6100 2743 6103
rect 3142 6100 3148 6112
rect 2731 6072 3148 6100
rect 2731 6069 2743 6072
rect 2685 6063 2743 6069
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 5460 6100 5488 6208
rect 7009 6205 7021 6208
rect 7055 6236 7067 6239
rect 7653 6239 7711 6245
rect 7653 6236 7665 6239
rect 7055 6208 7665 6236
rect 7055 6205 7067 6208
rect 7009 6199 7067 6205
rect 7653 6205 7665 6208
rect 7699 6205 7711 6239
rect 7653 6199 7711 6205
rect 5902 6128 5908 6180
rect 5960 6168 5966 6180
rect 6549 6171 6607 6177
rect 6549 6168 6561 6171
rect 5960 6140 6561 6168
rect 5960 6128 5966 6140
rect 6549 6137 6561 6140
rect 6595 6168 6607 6171
rect 6825 6171 6883 6177
rect 6825 6168 6837 6171
rect 6595 6140 6837 6168
rect 6595 6137 6607 6140
rect 6549 6131 6607 6137
rect 6825 6137 6837 6140
rect 6871 6137 6883 6171
rect 8036 6168 8064 6335
rect 9766 6264 9772 6316
rect 9824 6304 9830 6316
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 9824 6276 10333 6304
rect 9824 6264 9830 6276
rect 10321 6273 10333 6276
rect 10367 6304 10379 6307
rect 11333 6307 11391 6313
rect 11333 6304 11345 6307
rect 10367 6276 11345 6304
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 11333 6273 11345 6276
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 13357 6307 13415 6313
rect 13357 6273 13369 6307
rect 13403 6304 13415 6307
rect 13722 6304 13728 6316
rect 13403 6276 13728 6304
rect 13403 6273 13415 6276
rect 13357 6267 13415 6273
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 14108 6245 14136 6412
rect 14366 6400 14372 6452
rect 14424 6440 14430 6452
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 14424 6412 14473 6440
rect 14424 6400 14430 6412
rect 14461 6409 14473 6412
rect 14507 6409 14519 6443
rect 14461 6403 14519 6409
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 15473 6443 15531 6449
rect 15473 6440 15485 6443
rect 14700 6412 15485 6440
rect 14700 6400 14706 6412
rect 15473 6409 15485 6412
rect 15519 6440 15531 6443
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 15519 6412 15577 6440
rect 15519 6409 15531 6412
rect 15473 6403 15531 6409
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15565 6403 15623 6409
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 17589 6443 17647 6449
rect 17589 6440 17601 6443
rect 16908 6412 17601 6440
rect 16908 6400 16914 6412
rect 17589 6409 17601 6412
rect 17635 6409 17647 6443
rect 24670 6440 24676 6452
rect 24631 6412 24676 6440
rect 17589 6403 17647 6409
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 17218 6372 17224 6384
rect 17179 6344 17224 6372
rect 17218 6332 17224 6344
rect 17276 6332 17282 6384
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 15212 6276 16865 6304
rect 15212 6248 15240 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 18690 6264 18696 6316
rect 18748 6264 18754 6316
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6236 8263 6239
rect 14093 6239 14151 6245
rect 8251 6208 9536 6236
rect 8251 6205 8263 6208
rect 8205 6199 8263 6205
rect 8526 6171 8584 6177
rect 8526 6168 8538 6171
rect 8036 6140 8538 6168
rect 6825 6131 6883 6137
rect 8526 6137 8538 6140
rect 8572 6168 8584 6171
rect 8846 6168 8852 6180
rect 8572 6140 8852 6168
rect 8572 6137 8584 6140
rect 8526 6131 8584 6137
rect 8846 6128 8852 6140
rect 8904 6128 8910 6180
rect 9508 6112 9536 6208
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 14277 6239 14335 6245
rect 14277 6236 14289 6239
rect 14139 6208 14289 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 14277 6205 14289 6208
rect 14323 6205 14335 6239
rect 15194 6236 15200 6248
rect 15155 6208 15200 6236
rect 14277 6199 14335 6205
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 15473 6239 15531 6245
rect 15473 6205 15485 6239
rect 15519 6236 15531 6239
rect 15654 6236 15660 6248
rect 15519 6208 15660 6236
rect 15519 6205 15531 6208
rect 15473 6199 15531 6205
rect 15654 6196 15660 6208
rect 15712 6236 15718 6248
rect 15749 6239 15807 6245
rect 15749 6236 15761 6239
rect 15712 6208 15761 6236
rect 15712 6196 15718 6208
rect 15749 6205 15761 6208
rect 15795 6205 15807 6239
rect 16298 6236 16304 6248
rect 16259 6208 16304 6236
rect 15749 6199 15807 6205
rect 16298 6196 16304 6208
rect 16356 6196 16362 6248
rect 18708 6236 18736 6264
rect 18912 6239 18970 6245
rect 18912 6236 18924 6239
rect 18708 6208 18924 6236
rect 18912 6205 18924 6208
rect 18958 6236 18970 6239
rect 19337 6239 19395 6245
rect 19337 6236 19349 6239
rect 18958 6208 19349 6236
rect 18958 6205 18970 6208
rect 18912 6199 18970 6205
rect 19337 6205 19349 6208
rect 19383 6205 19395 6239
rect 19337 6199 19395 6205
rect 10042 6168 10048 6180
rect 10003 6140 10048 6168
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 10134 6128 10140 6180
rect 10192 6168 10198 6180
rect 10192 6140 10237 6168
rect 10192 6128 10198 6140
rect 12158 6128 12164 6180
rect 12216 6168 12222 6180
rect 12710 6168 12716 6180
rect 12216 6140 12716 6168
rect 12216 6128 12222 6140
rect 12710 6128 12716 6140
rect 12768 6128 12774 6180
rect 12805 6171 12863 6177
rect 12805 6137 12817 6171
rect 12851 6137 12863 6171
rect 12805 6131 12863 6137
rect 4120 6072 5488 6100
rect 5813 6103 5871 6109
rect 4120 6060 4126 6072
rect 5813 6069 5825 6103
rect 5859 6100 5871 6103
rect 6178 6100 6184 6112
rect 5859 6072 6184 6100
rect 5859 6069 5871 6072
rect 5813 6063 5871 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6362 6060 6368 6112
rect 6420 6100 6426 6112
rect 7098 6100 7104 6112
rect 6420 6072 7104 6100
rect 6420 6060 6426 6072
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 9122 6100 9128 6112
rect 9083 6072 9128 6100
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9490 6100 9496 6112
rect 9451 6072 9496 6100
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 10060 6100 10088 6128
rect 10965 6103 11023 6109
rect 10965 6100 10977 6103
rect 10060 6072 10977 6100
rect 10965 6069 10977 6072
rect 11011 6069 11023 6103
rect 10965 6063 11023 6069
rect 12342 6060 12348 6112
rect 12400 6100 12406 6112
rect 12820 6100 12848 6131
rect 15838 6100 15844 6112
rect 12400 6072 12848 6100
rect 15799 6072 15844 6100
rect 12400 6060 12406 6072
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 19015 6103 19073 6109
rect 19015 6069 19027 6103
rect 19061 6100 19073 6103
rect 19242 6100 19248 6112
rect 19061 6072 19248 6100
rect 19061 6069 19073 6072
rect 19015 6063 19073 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1535 5899 1593 5905
rect 1535 5865 1547 5899
rect 1581 5896 1593 5899
rect 1854 5896 1860 5908
rect 1581 5868 1860 5896
rect 1581 5865 1593 5868
rect 1535 5859 1593 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 2222 5896 2228 5908
rect 2004 5868 2228 5896
rect 2004 5856 2010 5868
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3602 5896 3608 5908
rect 3559 5868 3608 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 5261 5899 5319 5905
rect 5261 5865 5273 5899
rect 5307 5896 5319 5899
rect 5534 5896 5540 5908
rect 5307 5868 5540 5896
rect 5307 5865 5319 5868
rect 5261 5859 5319 5865
rect 5534 5856 5540 5868
rect 5592 5896 5598 5908
rect 6270 5896 6276 5908
rect 5592 5868 6276 5896
rect 5592 5856 5598 5868
rect 6270 5856 6276 5868
rect 6328 5896 6334 5908
rect 6641 5899 6699 5905
rect 6641 5896 6653 5899
rect 6328 5868 6653 5896
rect 6328 5856 6334 5868
rect 6641 5865 6653 5868
rect 6687 5865 6699 5899
rect 6641 5859 6699 5865
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 7285 5899 7343 5905
rect 7285 5896 7297 5899
rect 6788 5868 7297 5896
rect 6788 5856 6794 5868
rect 7285 5865 7297 5868
rect 7331 5865 7343 5899
rect 7285 5859 7343 5865
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 9122 5896 9128 5908
rect 7800 5868 9128 5896
rect 7800 5856 7806 5868
rect 5902 5828 5908 5840
rect 4126 5800 5908 5828
rect 1210 5720 1216 5772
rect 1268 5760 1274 5772
rect 1432 5763 1490 5769
rect 1432 5760 1444 5763
rect 1268 5732 1444 5760
rect 1268 5720 1274 5732
rect 1432 5729 1444 5732
rect 1478 5729 1490 5763
rect 3050 5760 3056 5772
rect 3011 5732 3056 5760
rect 1432 5723 1490 5729
rect 3050 5720 3056 5732
rect 3108 5760 3114 5772
rect 4126 5760 4154 5800
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 6083 5831 6141 5837
rect 6083 5797 6095 5831
rect 6129 5828 6141 5831
rect 6178 5828 6184 5840
rect 6129 5800 6184 5828
rect 6129 5797 6141 5800
rect 6083 5791 6141 5797
rect 6178 5788 6184 5800
rect 6236 5788 6242 5840
rect 8220 5837 8248 5868
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 9858 5896 9864 5908
rect 9819 5868 9864 5896
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 13722 5896 13728 5908
rect 13683 5868 13728 5896
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 14737 5899 14795 5905
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 14826 5896 14832 5908
rect 14783 5868 14832 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 14826 5856 14832 5868
rect 14884 5856 14890 5908
rect 15562 5896 15568 5908
rect 15523 5868 15568 5896
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 16298 5896 16304 5908
rect 16259 5868 16304 5896
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 17310 5896 17316 5908
rect 17271 5868 17316 5896
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 8205 5831 8263 5837
rect 8205 5797 8217 5831
rect 8251 5797 8263 5831
rect 8205 5791 8263 5797
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 9766 5828 9772 5840
rect 8803 5800 9772 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 9766 5788 9772 5800
rect 9824 5788 9830 5840
rect 10045 5831 10103 5837
rect 10045 5797 10057 5831
rect 10091 5828 10103 5831
rect 12710 5828 12716 5840
rect 10091 5800 12716 5828
rect 10091 5797 10103 5800
rect 10045 5791 10103 5797
rect 12710 5788 12716 5800
rect 12768 5788 12774 5840
rect 12802 5788 12808 5840
rect 12860 5828 12866 5840
rect 14461 5831 14519 5837
rect 12860 5800 12905 5828
rect 12860 5788 12866 5800
rect 14461 5797 14473 5831
rect 14507 5828 14519 5831
rect 14507 5800 20944 5828
rect 14507 5797 14519 5800
rect 14461 5791 14519 5797
rect 20916 5772 20944 5800
rect 4706 5760 4712 5772
rect 3108 5732 4154 5760
rect 4667 5732 4712 5760
rect 3108 5720 3114 5732
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 4893 5763 4951 5769
rect 4893 5729 4905 5763
rect 4939 5760 4951 5763
rect 7190 5760 7196 5772
rect 4939 5732 7196 5760
rect 4939 5729 4951 5732
rect 4893 5723 4951 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 9030 5760 9036 5772
rect 8991 5732 9036 5760
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 11238 5760 11244 5772
rect 11199 5732 11244 5760
rect 11238 5720 11244 5732
rect 11296 5720 11302 5772
rect 11330 5720 11336 5772
rect 11388 5760 11394 5772
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 11388 5732 11529 5760
rect 11388 5720 11394 5732
rect 11517 5729 11529 5732
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 14252 5763 14310 5769
rect 14252 5729 14264 5763
rect 14298 5760 14310 5763
rect 14550 5760 14556 5772
rect 14298 5732 14556 5760
rect 14298 5729 14310 5732
rect 14252 5723 14310 5729
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 15654 5760 15660 5772
rect 15615 5732 15660 5760
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 20898 5760 20904 5772
rect 20811 5732 20904 5760
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 2406 5692 2412 5704
rect 2367 5664 2412 5692
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 5718 5692 5724 5704
rect 5679 5664 5724 5692
rect 5718 5652 5724 5664
rect 5776 5692 5782 5704
rect 5994 5692 6000 5704
rect 5776 5664 6000 5692
rect 5776 5652 5782 5664
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7892 5664 8125 5692
rect 7892 5652 7898 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 9766 5692 9772 5704
rect 8812 5664 9772 5692
rect 8812 5652 8818 5664
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 11790 5692 11796 5704
rect 11751 5664 11796 5692
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 12989 5695 13047 5701
rect 12989 5692 13001 5695
rect 12124 5664 13001 5692
rect 12124 5652 12130 5664
rect 12989 5661 13001 5664
rect 13035 5692 13047 5695
rect 13446 5692 13452 5704
rect 13035 5664 13452 5692
rect 13035 5661 13047 5664
rect 12989 5655 13047 5661
rect 13446 5652 13452 5664
rect 13504 5652 13510 5704
rect 15562 5652 15568 5704
rect 15620 5692 15626 5704
rect 16853 5695 16911 5701
rect 16853 5692 16865 5695
rect 15620 5664 16865 5692
rect 15620 5652 15626 5664
rect 16853 5661 16865 5664
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 15105 5627 15163 5633
rect 15105 5593 15117 5627
rect 15151 5624 15163 5627
rect 15746 5624 15752 5636
rect 15151 5596 15752 5624
rect 15151 5593 15163 5596
rect 15105 5587 15163 5593
rect 15746 5584 15752 5596
rect 15804 5584 15810 5636
rect 2222 5556 2228 5568
rect 2183 5528 2228 5556
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 6914 5556 6920 5568
rect 6875 5528 6920 5556
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 10778 5556 10784 5568
rect 10739 5528 10784 5556
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 12434 5556 12440 5568
rect 12395 5528 12440 5556
rect 12434 5516 12440 5528
rect 12492 5516 12498 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 14458 5556 14464 5568
rect 12584 5528 14464 5556
rect 12584 5516 12590 5528
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 21085 5559 21143 5565
rect 21085 5525 21097 5559
rect 21131 5556 21143 5559
rect 22830 5556 22836 5568
rect 21131 5528 22836 5556
rect 21131 5525 21143 5528
rect 21085 5519 21143 5525
rect 22830 5516 22836 5528
rect 22888 5516 22894 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2958 5352 2964 5364
rect 2919 5324 2964 5352
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 8803 5355 8861 5361
rect 8803 5352 8815 5355
rect 6420 5324 8815 5352
rect 6420 5312 6426 5324
rect 8803 5321 8815 5324
rect 8849 5352 8861 5355
rect 9030 5352 9036 5364
rect 8849 5324 9036 5352
rect 8849 5321 8861 5324
rect 8803 5315 8861 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9309 5355 9367 5361
rect 9309 5321 9321 5355
rect 9355 5352 9367 5355
rect 10778 5352 10784 5364
rect 9355 5324 10784 5352
rect 9355 5321 9367 5324
rect 9309 5315 9367 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 12250 5352 12256 5364
rect 12211 5324 12256 5352
rect 12250 5312 12256 5324
rect 12308 5352 12314 5364
rect 12618 5352 12624 5364
rect 12308 5324 12624 5352
rect 12308 5312 12314 5324
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 13633 5355 13691 5361
rect 13633 5352 13645 5355
rect 12768 5324 13645 5352
rect 12768 5312 12774 5324
rect 13633 5321 13645 5324
rect 13679 5321 13691 5355
rect 13633 5315 13691 5321
rect 13909 5355 13967 5361
rect 13909 5321 13921 5355
rect 13955 5352 13967 5355
rect 15286 5352 15292 5364
rect 13955 5324 15292 5352
rect 13955 5321 13967 5324
rect 13909 5315 13967 5321
rect 15286 5312 15292 5324
rect 15344 5352 15350 5364
rect 15381 5355 15439 5361
rect 15381 5352 15393 5355
rect 15344 5324 15393 5352
rect 15344 5312 15350 5324
rect 15381 5321 15393 5324
rect 15427 5352 15439 5355
rect 15654 5352 15660 5364
rect 15427 5324 15660 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 20898 5352 20904 5364
rect 20859 5324 20904 5352
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 8205 5287 8263 5293
rect 8205 5253 8217 5287
rect 8251 5284 8263 5287
rect 8294 5284 8300 5296
rect 8251 5256 8300 5284
rect 8251 5253 8263 5256
rect 8205 5247 8263 5253
rect 8294 5244 8300 5256
rect 8352 5284 8358 5296
rect 8941 5287 8999 5293
rect 8941 5284 8953 5287
rect 8352 5256 8953 5284
rect 8352 5244 8358 5256
rect 8941 5253 8953 5256
rect 8987 5253 8999 5287
rect 8941 5247 8999 5253
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 9677 5287 9735 5293
rect 9677 5284 9689 5287
rect 9180 5256 9689 5284
rect 9180 5244 9186 5256
rect 9677 5253 9689 5256
rect 9723 5253 9735 5287
rect 9677 5247 9735 5253
rect 1762 5176 1768 5228
rect 1820 5216 1826 5228
rect 2041 5219 2099 5225
rect 2041 5216 2053 5219
rect 1820 5188 2053 5216
rect 1820 5176 1826 5188
rect 2041 5185 2053 5188
rect 2087 5185 2099 5219
rect 3142 5216 3148 5228
rect 3103 5188 3148 5216
rect 2041 5179 2099 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 6914 5216 6920 5228
rect 6875 5188 6920 5216
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7282 5216 7288 5228
rect 7243 5188 7288 5216
rect 7282 5176 7288 5188
rect 7340 5216 7346 5228
rect 7650 5216 7656 5228
rect 7340 5188 7656 5216
rect 7340 5176 7346 5188
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 8435 5188 9045 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 9033 5185 9045 5188
rect 9079 5216 9091 5219
rect 9214 5216 9220 5228
rect 9079 5188 9220 5216
rect 9079 5185 9091 5188
rect 9033 5179 9091 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 10796 5216 10824 5312
rect 11440 5256 12572 5284
rect 10796 5188 11284 5216
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 1946 5148 1952 5160
rect 1903 5120 1952 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 1946 5108 1952 5120
rect 2004 5108 2010 5160
rect 2133 5151 2191 5157
rect 2133 5117 2145 5151
rect 2179 5148 2191 5151
rect 2958 5148 2964 5160
rect 2179 5120 2964 5148
rect 2179 5117 2191 5120
rect 2133 5111 2191 5117
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 3602 5148 3608 5160
rect 3563 5120 3608 5148
rect 3602 5108 3608 5120
rect 3660 5148 3666 5160
rect 4157 5151 4215 5157
rect 4157 5148 4169 5151
rect 3660 5120 4169 5148
rect 3660 5108 3666 5120
rect 4157 5117 4169 5120
rect 4203 5117 4215 5151
rect 5534 5148 5540 5160
rect 5495 5120 5540 5148
rect 4157 5111 4215 5117
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 8665 5151 8723 5157
rect 8665 5117 8677 5151
rect 8711 5148 8723 5151
rect 8938 5148 8944 5160
rect 8711 5120 8944 5148
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 8938 5108 8944 5120
rect 8996 5108 9002 5160
rect 11256 5157 11284 5188
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 11057 5151 11115 5157
rect 11057 5148 11069 5151
rect 10735 5120 11069 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 11057 5117 11069 5120
rect 11103 5117 11115 5151
rect 11057 5111 11115 5117
rect 11241 5151 11299 5157
rect 11241 5117 11253 5151
rect 11287 5148 11299 5151
rect 11330 5148 11336 5160
rect 11287 5120 11336 5148
rect 11287 5117 11299 5120
rect 11241 5111 11299 5117
rect 2685 5083 2743 5089
rect 2685 5049 2697 5083
rect 2731 5080 2743 5083
rect 3050 5080 3056 5092
rect 2731 5052 3056 5080
rect 2731 5049 2743 5052
rect 2685 5043 2743 5049
rect 3050 5040 3056 5052
rect 3108 5040 3114 5092
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 5951 5052 6561 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 6549 5049 6561 5052
rect 6595 5080 6607 5083
rect 7009 5083 7067 5089
rect 7009 5080 7021 5083
rect 6595 5052 7021 5080
rect 6595 5049 6607 5052
rect 6549 5043 6607 5049
rect 7009 5049 7021 5052
rect 7055 5049 7067 5083
rect 7009 5043 7067 5049
rect 8294 5040 8300 5092
rect 8352 5080 8358 5092
rect 10704 5080 10732 5111
rect 8352 5052 10732 5080
rect 11072 5080 11100 5111
rect 11330 5108 11336 5120
rect 11388 5108 11394 5160
rect 11440 5080 11468 5256
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5216 11575 5219
rect 12434 5216 12440 5228
rect 11563 5188 12440 5216
rect 11563 5185 11575 5188
rect 11517 5179 11575 5185
rect 12434 5176 12440 5188
rect 12492 5176 12498 5228
rect 12544 5216 12572 5256
rect 13354 5244 13360 5296
rect 13412 5284 13418 5296
rect 20073 5287 20131 5293
rect 13412 5256 15884 5284
rect 13412 5244 13418 5256
rect 12894 5216 12900 5228
rect 12544 5188 12900 5216
rect 12894 5176 12900 5188
rect 12952 5216 12958 5228
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 12952 5188 14105 5216
rect 12952 5176 12958 5188
rect 14093 5185 14105 5188
rect 14139 5216 14151 5219
rect 15470 5216 15476 5228
rect 14139 5188 15476 5216
rect 14139 5185 14151 5188
rect 14093 5179 14151 5185
rect 14476 5157 14504 5188
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 13449 5151 13507 5157
rect 13449 5148 13461 5151
rect 11072 5052 11468 5080
rect 11808 5120 13461 5148
rect 8352 5040 8358 5052
rect 3068 5012 3096 5040
rect 3602 5012 3608 5024
rect 3068 4984 3608 5012
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 4617 5015 4675 5021
rect 4617 4981 4629 5015
rect 4663 5012 4675 5015
rect 4706 5012 4712 5024
rect 4663 4984 4712 5012
rect 4663 4981 4675 4984
rect 4617 4975 4675 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 4985 5015 5043 5021
rect 4985 4981 4997 5015
rect 5031 5012 5043 5015
rect 5350 5012 5356 5024
rect 5031 4984 5356 5012
rect 5031 4981 5043 4984
rect 4985 4975 5043 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 6880 4984 8401 5012
rect 6880 4972 6886 4984
rect 8389 4981 8401 4984
rect 8435 5012 8447 5015
rect 8481 5015 8539 5021
rect 8481 5012 8493 5015
rect 8435 4984 8493 5012
rect 8435 4981 8447 4984
rect 8389 4975 8447 4981
rect 8481 4981 8493 4984
rect 8527 4981 8539 5015
rect 8481 4975 8539 4981
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 11238 5012 11244 5024
rect 10744 4984 11244 5012
rect 10744 4972 10750 4984
rect 11238 4972 11244 4984
rect 11296 5012 11302 5024
rect 11808 5021 11836 5120
rect 13449 5117 13461 5120
rect 13495 5117 13507 5151
rect 13449 5111 13507 5117
rect 14461 5151 14519 5157
rect 14461 5117 14473 5151
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 14737 5151 14795 5157
rect 14737 5117 14749 5151
rect 14783 5148 14795 5151
rect 15378 5148 15384 5160
rect 14783 5120 15384 5148
rect 14783 5117 14795 5120
rect 14737 5111 14795 5117
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 15856 5157 15884 5256
rect 20073 5253 20085 5287
rect 20119 5284 20131 5287
rect 21542 5284 21548 5296
rect 20119 5256 21548 5284
rect 20119 5253 20131 5256
rect 20073 5247 20131 5253
rect 21542 5244 21548 5256
rect 21600 5244 21606 5296
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 15887 5120 16773 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 16761 5117 16773 5120
rect 16807 5117 16819 5151
rect 16761 5111 16819 5117
rect 17862 5108 17868 5160
rect 17920 5148 17926 5160
rect 18084 5151 18142 5157
rect 18084 5148 18096 5151
rect 17920 5120 18096 5148
rect 17920 5108 17926 5120
rect 18084 5117 18096 5120
rect 18130 5148 18142 5151
rect 18509 5151 18567 5157
rect 18509 5148 18521 5151
rect 18130 5120 18521 5148
rect 18130 5117 18142 5120
rect 18084 5111 18142 5117
rect 18509 5117 18521 5120
rect 18555 5117 18567 5151
rect 18509 5111 18567 5117
rect 19242 5108 19248 5160
rect 19300 5148 19306 5160
rect 19889 5151 19947 5157
rect 19889 5148 19901 5151
rect 19300 5120 19901 5148
rect 19300 5108 19306 5120
rect 19889 5117 19901 5120
rect 19935 5148 19947 5151
rect 20441 5151 20499 5157
rect 20441 5148 20453 5151
rect 19935 5120 20453 5148
rect 19935 5117 19947 5120
rect 19889 5111 19947 5117
rect 20441 5117 20453 5120
rect 20487 5117 20499 5151
rect 20441 5111 20499 5117
rect 12618 5040 12624 5092
rect 12676 5080 12682 5092
rect 12758 5083 12816 5089
rect 12758 5080 12770 5083
rect 12676 5052 12770 5080
rect 12676 5040 12682 5052
rect 12758 5049 12770 5052
rect 12804 5049 12816 5083
rect 12758 5043 12816 5049
rect 12894 5040 12900 5092
rect 12952 5080 12958 5092
rect 15749 5083 15807 5089
rect 15749 5080 15761 5083
rect 12952 5052 15761 5080
rect 12952 5040 12958 5052
rect 15749 5049 15761 5052
rect 15795 5049 15807 5083
rect 15749 5043 15807 5049
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 11296 4984 11805 5012
rect 11296 4972 11302 4984
rect 11793 4981 11805 4984
rect 11839 4981 11851 5015
rect 13354 5012 13360 5024
rect 13315 4984 13360 5012
rect 11793 4975 11851 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13449 5015 13507 5021
rect 13449 4981 13461 5015
rect 13495 5012 13507 5015
rect 13909 5015 13967 5021
rect 13909 5012 13921 5015
rect 13495 4984 13921 5012
rect 13495 4981 13507 4984
rect 13449 4975 13507 4981
rect 13909 4981 13921 4984
rect 13955 4981 13967 5015
rect 14274 5012 14280 5024
rect 14235 4984 14280 5012
rect 13909 4975 13967 4981
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 18187 5015 18245 5021
rect 18187 4981 18199 5015
rect 18233 5012 18245 5015
rect 18414 5012 18420 5024
rect 18233 4984 18420 5012
rect 18233 4981 18245 4984
rect 18187 4975 18245 4981
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1210 4768 1216 4820
rect 1268 4808 1274 4820
rect 2225 4811 2283 4817
rect 2225 4808 2237 4811
rect 1268 4780 2237 4808
rect 1268 4768 1274 4780
rect 2225 4777 2237 4780
rect 2271 4777 2283 4811
rect 2225 4771 2283 4777
rect 3053 4811 3111 4817
rect 3053 4777 3065 4811
rect 3099 4808 3111 4811
rect 4430 4808 4436 4820
rect 3099 4780 4436 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 4430 4768 4436 4780
rect 4488 4768 4494 4820
rect 4982 4808 4988 4820
rect 4943 4780 4988 4808
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5994 4808 6000 4820
rect 5955 4780 6000 4808
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 8018 4808 8024 4820
rect 6098 4780 8024 4808
rect 1946 4740 1952 4752
rect 1907 4712 1952 4740
rect 1946 4700 1952 4712
rect 2004 4700 2010 4752
rect 2406 4740 2412 4752
rect 2367 4712 2412 4740
rect 2406 4700 2412 4712
rect 2464 4740 2470 4752
rect 2958 4740 2964 4752
rect 2464 4712 2964 4740
rect 2464 4700 2470 4712
rect 2958 4700 2964 4712
rect 3016 4740 3022 4752
rect 3421 4743 3479 4749
rect 3421 4740 3433 4743
rect 3016 4712 3433 4740
rect 3016 4700 3022 4712
rect 3421 4709 3433 4712
rect 3467 4709 3479 4743
rect 5442 4740 5448 4752
rect 3421 4703 3479 4709
rect 5184 4712 5448 4740
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 5184 4681 5212 4712
rect 5442 4700 5448 4712
rect 5500 4740 5506 4752
rect 6098 4740 6126 4780
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 9030 4808 9036 4820
rect 8991 4780 9036 4808
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 9861 4811 9919 4817
rect 9861 4808 9873 4811
rect 9824 4780 9873 4808
rect 9824 4768 9830 4780
rect 9861 4777 9873 4780
rect 9907 4777 9919 4811
rect 11330 4808 11336 4820
rect 11291 4780 11336 4808
rect 9861 4771 9919 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 12802 4808 12808 4820
rect 12759 4780 12808 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 14550 4808 14556 4820
rect 14511 4780 14556 4808
rect 14550 4768 14556 4780
rect 14608 4768 14614 4820
rect 14734 4768 14740 4820
rect 14792 4808 14798 4820
rect 15381 4811 15439 4817
rect 15381 4808 15393 4811
rect 14792 4780 15393 4808
rect 14792 4768 14798 4780
rect 15381 4777 15393 4780
rect 15427 4777 15439 4811
rect 15381 4771 15439 4777
rect 5500 4712 6126 4740
rect 5500 4700 5506 4712
rect 6178 4700 6184 4752
rect 6236 4740 6242 4752
rect 6457 4743 6515 4749
rect 6457 4740 6469 4743
rect 6236 4712 6469 4740
rect 6236 4700 6242 4712
rect 6457 4709 6469 4712
rect 6503 4740 6515 4743
rect 8662 4740 8668 4752
rect 6503 4712 8668 4740
rect 6503 4709 6515 4712
rect 6457 4703 6515 4709
rect 8662 4700 8668 4712
rect 8720 4700 8726 4752
rect 10502 4740 10508 4752
rect 10463 4712 10508 4740
rect 10502 4700 10508 4712
rect 10560 4700 10566 4752
rect 12250 4700 12256 4752
rect 12308 4740 12314 4752
rect 13265 4743 13323 4749
rect 13265 4740 13277 4743
rect 12308 4712 13277 4740
rect 12308 4700 12314 4712
rect 13265 4709 13277 4712
rect 13311 4740 13323 4743
rect 13354 4740 13360 4752
rect 13311 4712 13360 4740
rect 13311 4709 13323 4712
rect 13265 4703 13323 4709
rect 13354 4700 13360 4712
rect 13412 4700 13418 4752
rect 15838 4740 15844 4752
rect 15304 4712 15844 4740
rect 15304 4684 15332 4712
rect 15838 4700 15844 4712
rect 15896 4700 15902 4752
rect 1535 4675 1593 4681
rect 1535 4641 1547 4675
rect 1581 4672 1593 4675
rect 5169 4675 5227 4681
rect 1581 4644 3280 4672
rect 1581 4641 1593 4644
rect 1535 4635 1593 4641
rect 106 4564 112 4616
rect 164 4604 170 4616
rect 2774 4604 2780 4616
rect 164 4576 2544 4604
rect 2735 4576 2780 4604
rect 164 4564 170 4576
rect 2516 4536 2544 4576
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 2574 4539 2632 4545
rect 2574 4536 2586 4539
rect 2516 4508 2586 4536
rect 2574 4505 2586 4508
rect 2620 4536 2632 4539
rect 3142 4536 3148 4548
rect 2620 4508 3148 4536
rect 2620 4505 2632 4508
rect 2574 4499 2632 4505
rect 3142 4496 3148 4508
rect 3200 4496 3206 4548
rect 3252 4536 3280 4644
rect 5169 4641 5181 4675
rect 5215 4641 5227 4675
rect 5350 4672 5356 4684
rect 5311 4644 5356 4672
rect 5169 4635 5227 4641
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 6822 4681 6828 4684
rect 6796 4675 6828 4681
rect 6796 4641 6808 4675
rect 6796 4635 6828 4641
rect 6822 4632 6828 4635
rect 6880 4632 6886 4684
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8294 4672 8300 4684
rect 8076 4644 8300 4672
rect 8076 4632 8082 4644
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8478 4672 8484 4684
rect 8439 4644 8484 4672
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 11882 4632 11888 4684
rect 11940 4672 11946 4684
rect 11977 4675 12035 4681
rect 11977 4672 11989 4675
rect 11940 4644 11989 4672
rect 11940 4632 11946 4644
rect 11977 4641 11989 4644
rect 12023 4672 12035 4675
rect 12526 4672 12532 4684
rect 12023 4644 12532 4672
rect 12023 4641 12035 4644
rect 11977 4635 12035 4641
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 15286 4672 15292 4684
rect 15247 4644 15292 4672
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 15378 4632 15384 4684
rect 15436 4672 15442 4684
rect 15749 4675 15807 4681
rect 15749 4672 15761 4675
rect 15436 4644 15761 4672
rect 15436 4632 15442 4644
rect 15749 4641 15761 4644
rect 15795 4641 15807 4675
rect 15749 4635 15807 4641
rect 16853 4675 16911 4681
rect 16853 4641 16865 4675
rect 16899 4672 16911 4675
rect 17218 4672 17224 4684
rect 16899 4644 17224 4672
rect 16899 4641 16911 4644
rect 16853 4635 16911 4641
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 18414 4632 18420 4684
rect 18472 4672 18478 4684
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 18472 4644 18705 4672
rect 18472 4632 18478 4644
rect 18693 4641 18705 4644
rect 18739 4641 18751 4675
rect 18693 4635 18751 4641
rect 8754 4604 8760 4616
rect 8715 4576 8760 4604
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 9640 4576 10425 4604
rect 9640 4564 9646 4576
rect 10413 4573 10425 4576
rect 10459 4604 10471 4607
rect 10870 4604 10876 4616
rect 10459 4576 10876 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 11057 4607 11115 4613
rect 11057 4573 11069 4607
rect 11103 4604 11115 4607
rect 11238 4604 11244 4616
rect 11103 4576 11244 4604
rect 11103 4573 11115 4576
rect 11057 4567 11115 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 13173 4607 13231 4613
rect 13173 4604 13185 4607
rect 13044 4576 13185 4604
rect 13044 4564 13050 4576
rect 13173 4573 13185 4576
rect 13219 4573 13231 4607
rect 13446 4604 13452 4616
rect 13407 4576 13452 4604
rect 13173 4567 13231 4573
rect 13446 4564 13452 4576
rect 13504 4564 13510 4616
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14366 4604 14372 4616
rect 14323 4576 14372 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14366 4564 14372 4576
rect 14424 4604 14430 4616
rect 15396 4604 15424 4632
rect 14424 4576 15424 4604
rect 14424 4564 14430 4576
rect 10042 4536 10048 4548
rect 3252 4508 10048 4536
rect 10042 4496 10048 4508
rect 10100 4496 10106 4548
rect 12161 4539 12219 4545
rect 12161 4505 12173 4539
rect 12207 4536 12219 4539
rect 13630 4536 13636 4548
rect 12207 4508 13636 4536
rect 12207 4505 12219 4508
rect 12161 4499 12219 4505
rect 13630 4496 13636 4508
rect 13688 4496 13694 4548
rect 15286 4496 15292 4548
rect 15344 4536 15350 4548
rect 17037 4539 17095 4545
rect 17037 4536 17049 4539
rect 15344 4508 17049 4536
rect 15344 4496 15350 4508
rect 17037 4505 17049 4508
rect 17083 4505 17095 4539
rect 17037 4499 17095 4505
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 2685 4471 2743 4477
rect 2685 4468 2697 4471
rect 2372 4440 2697 4468
rect 2372 4428 2378 4440
rect 2685 4437 2697 4440
rect 2731 4437 2743 4471
rect 2685 4431 2743 4437
rect 3050 4428 3056 4480
rect 3108 4468 3114 4480
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 3108 4440 3801 4468
rect 3108 4428 3114 4440
rect 3789 4437 3801 4440
rect 3835 4468 3847 4471
rect 4338 4468 4344 4480
rect 3835 4440 4344 4468
rect 3835 4437 3847 4440
rect 3789 4431 3847 4437
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 4614 4468 4620 4480
rect 4575 4440 4620 4468
rect 4614 4428 4620 4440
rect 4672 4468 4678 4480
rect 6362 4468 6368 4480
rect 4672 4440 6368 4468
rect 4672 4428 4678 4440
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 6595 4471 6653 4477
rect 6595 4468 6607 4471
rect 6512 4440 6607 4468
rect 6512 4428 6518 4440
rect 6595 4437 6607 4440
rect 6641 4437 6653 4471
rect 6730 4468 6736 4480
rect 6691 4440 6736 4468
rect 6595 4431 6653 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 6917 4471 6975 4477
rect 6917 4437 6929 4471
rect 6963 4468 6975 4471
rect 7006 4468 7012 4480
rect 6963 4440 7012 4468
rect 6963 4437 6975 4440
rect 6917 4431 6975 4437
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 7834 4468 7840 4480
rect 7795 4440 7840 4468
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 16390 4468 16396 4480
rect 16351 4440 16396 4468
rect 16390 4428 16396 4440
rect 16448 4428 16454 4480
rect 18874 4468 18880 4480
rect 18835 4440 18880 4468
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1578 4224 1584 4276
rect 1636 4264 1642 4276
rect 1673 4267 1731 4273
rect 1673 4264 1685 4267
rect 1636 4236 1685 4264
rect 1636 4224 1642 4236
rect 1673 4233 1685 4236
rect 1719 4233 1731 4267
rect 1673 4227 1731 4233
rect 3053 4267 3111 4273
rect 3053 4233 3065 4267
rect 3099 4264 3111 4267
rect 3234 4264 3240 4276
rect 3099 4236 3240 4264
rect 3099 4233 3111 4236
rect 3053 4227 3111 4233
rect 3234 4224 3240 4236
rect 3292 4264 3298 4276
rect 3786 4264 3792 4276
rect 3292 4236 3792 4264
rect 3292 4224 3298 4236
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 4062 4264 4068 4276
rect 4023 4236 4068 4264
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 6362 4264 6368 4276
rect 5368 4236 6368 4264
rect 2314 4156 2320 4208
rect 2372 4196 2378 4208
rect 4246 4196 4252 4208
rect 2372 4168 4252 4196
rect 2372 4156 2378 4168
rect 4246 4156 4252 4168
rect 4304 4196 4310 4208
rect 4433 4199 4491 4205
rect 4433 4196 4445 4199
rect 4304 4168 4445 4196
rect 4304 4156 4310 4168
rect 4433 4165 4445 4168
rect 4479 4165 4491 4199
rect 4433 4159 4491 4165
rect 4614 4156 4620 4208
rect 4672 4196 4678 4208
rect 4755 4199 4813 4205
rect 4755 4196 4767 4199
rect 4672 4168 4767 4196
rect 4672 4156 4678 4168
rect 4755 4165 4767 4168
rect 4801 4165 4813 4199
rect 4890 4196 4896 4208
rect 4851 4168 4896 4196
rect 4755 4159 4813 4165
rect 4890 4156 4896 4168
rect 4948 4196 4954 4208
rect 5368 4196 5396 4236
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 6454 4224 6460 4276
rect 6512 4264 6518 4276
rect 6641 4267 6699 4273
rect 6641 4264 6653 4267
rect 6512 4236 6653 4264
rect 6512 4224 6518 4236
rect 6641 4233 6653 4236
rect 6687 4233 6699 4267
rect 6641 4227 6699 4233
rect 10502 4224 10508 4276
rect 10560 4264 10566 4276
rect 10781 4267 10839 4273
rect 10781 4264 10793 4267
rect 10560 4236 10793 4264
rect 10560 4224 10566 4236
rect 10781 4233 10793 4236
rect 10827 4264 10839 4267
rect 17034 4264 17040 4276
rect 10827 4236 17040 4264
rect 10827 4233 10839 4236
rect 10781 4227 10839 4233
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 18414 4224 18420 4276
rect 18472 4264 18478 4276
rect 18877 4267 18935 4273
rect 18877 4264 18889 4267
rect 18472 4236 18889 4264
rect 18472 4224 18478 4236
rect 18877 4233 18889 4236
rect 18923 4233 18935 4267
rect 18877 4227 18935 4233
rect 4948 4168 5396 4196
rect 4948 4156 4954 4168
rect 5442 4156 5448 4208
rect 5500 4196 5506 4208
rect 5629 4199 5687 4205
rect 5629 4196 5641 4199
rect 5500 4168 5641 4196
rect 5500 4156 5506 4168
rect 5629 4165 5641 4168
rect 5675 4165 5687 4199
rect 9401 4199 9459 4205
rect 9401 4196 9413 4199
rect 5629 4159 5687 4165
rect 6380 4168 9413 4196
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4264 4100 4997 4128
rect 1486 4060 1492 4072
rect 1447 4032 1492 4060
rect 1486 4020 1492 4032
rect 1544 4020 1550 4072
rect 2958 4060 2964 4072
rect 2919 4032 2964 4060
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 3510 4060 3516 4072
rect 3200 4032 3516 4060
rect 3200 4020 3206 4032
rect 3510 4020 3516 4032
rect 3568 4060 3574 4072
rect 3697 4063 3755 4069
rect 3697 4060 3709 4063
rect 3568 4032 3709 4060
rect 3568 4020 3574 4032
rect 3697 4029 3709 4032
rect 3743 4060 3755 4063
rect 4062 4060 4068 4072
rect 3743 4032 4068 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 2372 3896 2421 3924
rect 2372 3884 2378 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 2774 3924 2780 3936
rect 2735 3896 2780 3924
rect 2409 3887 2467 3893
rect 2774 3884 2780 3896
rect 2832 3924 2838 3936
rect 4264 3924 4292 4100
rect 4985 4097 4997 4100
rect 5031 4128 5043 4131
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5031 4100 5549 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 6178 4128 6184 4140
rect 6139 4100 6184 4128
rect 5537 4091 5595 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 4338 4020 4344 4072
rect 4396 4060 4402 4072
rect 6380 4060 6408 4168
rect 9401 4165 9413 4168
rect 9447 4196 9459 4199
rect 9493 4199 9551 4205
rect 9493 4196 9505 4199
rect 9447 4168 9505 4196
rect 9447 4165 9459 4168
rect 9401 4159 9459 4165
rect 9493 4165 9505 4168
rect 9539 4165 9551 4199
rect 10686 4196 10692 4208
rect 9493 4159 9551 4165
rect 9646 4168 10692 4196
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4128 6883 4131
rect 6914 4128 6920 4140
rect 6871 4100 6920 4128
rect 6871 4097 6883 4100
rect 6825 4091 6883 4097
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 9646 4128 9674 4168
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 11057 4199 11115 4205
rect 11057 4196 11069 4199
rect 10928 4168 11069 4196
rect 10928 4156 10934 4168
rect 11057 4165 11069 4168
rect 11103 4165 11115 4199
rect 11882 4196 11888 4208
rect 11843 4168 11888 4196
rect 11057 4159 11115 4165
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 12250 4196 12256 4208
rect 12211 4168 12256 4196
rect 12250 4156 12256 4168
rect 12308 4156 12314 4208
rect 14093 4199 14151 4205
rect 14093 4165 14105 4199
rect 14139 4196 14151 4199
rect 14642 4196 14648 4208
rect 14139 4168 14648 4196
rect 14139 4165 14151 4168
rect 14093 4159 14151 4165
rect 14642 4156 14648 4168
rect 14700 4156 14706 4208
rect 16761 4199 16819 4205
rect 16761 4196 16773 4199
rect 14936 4168 16773 4196
rect 9766 4128 9772 4140
rect 8128 4100 9674 4128
rect 9727 4100 9772 4128
rect 8128 4069 8156 4100
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12802 4128 12808 4140
rect 11848 4100 12808 4128
rect 11848 4088 11854 4100
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 14936 4137 14964 4168
rect 16761 4165 16773 4168
rect 16807 4165 16819 4199
rect 16761 4159 16819 4165
rect 14921 4131 14979 4137
rect 14921 4128 14933 4131
rect 13044 4100 14933 4128
rect 13044 4088 13050 4100
rect 14921 4097 14933 4100
rect 14967 4097 14979 4131
rect 14921 4091 14979 4097
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4128 16267 4131
rect 16390 4128 16396 4140
rect 16255 4100 16396 4128
rect 16255 4097 16267 4100
rect 16209 4091 16267 4097
rect 16390 4088 16396 4100
rect 16448 4128 16454 4140
rect 18187 4131 18245 4137
rect 18187 4128 18199 4131
rect 16448 4100 18199 4128
rect 16448 4088 16454 4100
rect 18187 4097 18199 4100
rect 18233 4097 18245 4131
rect 18187 4091 18245 4097
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 4396 4032 6408 4060
rect 7944 4032 8125 4060
rect 4396 4020 4402 4032
rect 4614 3992 4620 4004
rect 4575 3964 4620 3992
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 5537 3995 5595 4001
rect 5537 3961 5549 3995
rect 5583 3992 5595 3995
rect 6822 3992 6828 4004
rect 5583 3964 6828 3992
rect 5583 3961 5595 3964
rect 5537 3955 5595 3961
rect 6822 3952 6828 3964
rect 6880 3992 6886 4004
rect 7285 3995 7343 4001
rect 7285 3992 7297 3995
rect 6880 3964 7297 3992
rect 6880 3952 6886 3964
rect 7285 3961 7297 3964
rect 7331 3961 7343 3995
rect 7285 3955 7343 3961
rect 4338 3924 4344 3936
rect 2832 3896 4344 3924
rect 2832 3884 2838 3896
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 5261 3927 5319 3933
rect 5261 3924 5273 3927
rect 5132 3896 5273 3924
rect 5132 3884 5138 3896
rect 5261 3893 5273 3896
rect 5307 3924 5319 3927
rect 5350 3924 5356 3936
rect 5307 3896 5356 3924
rect 5307 3893 5319 3896
rect 5261 3887 5319 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 7944 3933 7972 4032
rect 8113 4029 8125 4032
rect 8159 4029 8171 4063
rect 8113 4023 8171 4029
rect 8478 4020 8484 4072
rect 8536 4060 8542 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8536 4032 8677 4060
rect 8536 4020 8542 4032
rect 8665 4029 8677 4032
rect 8711 4060 8723 4063
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8711 4032 9137 4060
rect 8711 4029 8723 4032
rect 8665 4023 8723 4029
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 11238 4060 11244 4072
rect 11199 4032 11244 4060
rect 9125 4023 9183 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 12618 4060 12624 4072
rect 12579 4032 12624 4060
rect 12618 4020 12624 4032
rect 12676 4060 12682 4072
rect 13725 4063 13783 4069
rect 12676 4032 13169 4060
rect 12676 4020 12682 4032
rect 8846 3992 8852 4004
rect 8807 3964 8852 3992
rect 8846 3952 8852 3964
rect 8904 3952 8910 4004
rect 9401 3995 9459 4001
rect 9401 3961 9413 3995
rect 9447 3992 9459 3995
rect 9858 3992 9864 4004
rect 9447 3964 9864 3992
rect 9447 3961 9459 3964
rect 9401 3955 9459 3961
rect 9858 3952 9864 3964
rect 9916 3952 9922 4004
rect 10413 3995 10471 4001
rect 10413 3961 10425 3995
rect 10459 3992 10471 3995
rect 11514 3992 11520 4004
rect 10459 3964 11520 3992
rect 10459 3961 10471 3964
rect 10413 3955 10471 3961
rect 11514 3952 11520 3964
rect 11572 3952 11578 4004
rect 13141 4001 13169 4032
rect 13725 4029 13737 4063
rect 13771 4060 13783 4063
rect 18084 4063 18142 4069
rect 18084 4060 18096 4063
rect 13771 4032 14504 4060
rect 13771 4029 13783 4032
rect 13725 4023 13783 4029
rect 13126 3995 13184 4001
rect 13126 3961 13138 3995
rect 13172 3992 13184 3995
rect 13354 3992 13360 4004
rect 13172 3964 13360 3992
rect 13172 3961 13184 3964
rect 13126 3955 13184 3961
rect 13354 3952 13360 3964
rect 13412 3952 13418 4004
rect 6641 3927 6699 3933
rect 6641 3924 6653 3927
rect 6512 3896 6653 3924
rect 6512 3884 6518 3896
rect 6641 3893 6653 3896
rect 6687 3893 6699 3927
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 7887 3896 7941 3924
rect 6641 3887 6699 3893
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 7929 3887 7987 3893
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 10042 3924 10048 3936
rect 8996 3896 10048 3924
rect 8996 3884 9002 3896
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 11379 3927 11437 3933
rect 11379 3893 11391 3927
rect 11425 3924 11437 3927
rect 12342 3924 12348 3936
rect 11425 3896 12348 3924
rect 11425 3893 11437 3896
rect 11379 3887 11437 3893
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 14366 3924 14372 3936
rect 14327 3896 14372 3924
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 14476 3924 14504 4032
rect 17512 4032 18096 4060
rect 14642 3992 14648 4004
rect 14603 3964 14648 3992
rect 14642 3952 14648 3964
rect 14700 3952 14706 4004
rect 14737 3995 14795 4001
rect 14737 3961 14749 3995
rect 14783 3992 14795 3995
rect 15746 3992 15752 4004
rect 14783 3964 15752 3992
rect 14783 3961 14795 3964
rect 14737 3955 14795 3961
rect 14752 3924 14780 3955
rect 15746 3952 15752 3964
rect 15804 3952 15810 4004
rect 16025 3995 16083 4001
rect 16025 3961 16037 3995
rect 16071 3992 16083 3995
rect 16298 3992 16304 4004
rect 16071 3964 16304 3992
rect 16071 3961 16083 3964
rect 16025 3955 16083 3961
rect 16298 3952 16304 3964
rect 16356 3952 16362 4004
rect 16390 3952 16396 4004
rect 16448 3992 16454 4004
rect 17512 3992 17540 4032
rect 18084 4029 18096 4032
rect 18130 4060 18142 4063
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 18130 4032 18521 4060
rect 18130 4029 18142 4032
rect 18084 4023 18142 4029
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 19128 4063 19186 4069
rect 19128 4029 19140 4063
rect 19174 4060 19186 4063
rect 19174 4029 19196 4060
rect 19128 4023 19196 4029
rect 16448 3964 17540 3992
rect 16448 3952 16454 3964
rect 17586 3952 17592 4004
rect 17644 3992 17650 4004
rect 19168 3992 19196 4023
rect 19521 3995 19579 4001
rect 19521 3992 19533 3995
rect 17644 3964 19533 3992
rect 17644 3952 17650 3964
rect 19521 3961 19533 3964
rect 19567 3961 19579 3995
rect 19521 3955 19579 3961
rect 14476 3896 14780 3924
rect 15657 3927 15715 3933
rect 15657 3893 15669 3927
rect 15703 3924 15715 3927
rect 15838 3924 15844 3936
rect 15703 3896 15844 3924
rect 15703 3893 15715 3896
rect 15657 3887 15715 3893
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 17218 3924 17224 3936
rect 17131 3896 17224 3924
rect 17218 3884 17224 3896
rect 17276 3924 17282 3936
rect 17402 3924 17408 3936
rect 17276 3896 17408 3924
rect 17276 3884 17282 3896
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 17494 3884 17500 3936
rect 17552 3924 17558 3936
rect 19199 3927 19257 3933
rect 19199 3924 19211 3927
rect 17552 3896 19211 3924
rect 17552 3884 17558 3896
rect 19199 3893 19211 3896
rect 19245 3893 19257 3927
rect 19199 3887 19257 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1394 3680 1400 3732
rect 1452 3720 1458 3732
rect 1857 3723 1915 3729
rect 1857 3720 1869 3723
rect 1452 3692 1869 3720
rect 1452 3680 1458 3692
rect 1857 3689 1869 3692
rect 1903 3689 1915 3723
rect 3510 3720 3516 3732
rect 3471 3692 3516 3720
rect 1857 3683 1915 3689
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 4203 3723 4261 3729
rect 4203 3720 4215 3723
rect 3752 3692 4215 3720
rect 3752 3680 3758 3692
rect 4203 3689 4215 3692
rect 4249 3689 4261 3723
rect 4203 3683 4261 3689
rect 4614 3680 4620 3732
rect 4672 3720 4678 3732
rect 5077 3723 5135 3729
rect 5077 3720 5089 3723
rect 4672 3692 5089 3720
rect 4672 3680 4678 3692
rect 5077 3689 5089 3692
rect 5123 3720 5135 3723
rect 6178 3720 6184 3732
rect 5123 3692 6184 3720
rect 5123 3689 5135 3692
rect 5077 3683 5135 3689
rect 6178 3680 6184 3692
rect 6236 3680 6242 3732
rect 6454 3720 6460 3732
rect 6415 3692 6460 3720
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 8018 3720 8024 3732
rect 7979 3692 8024 3720
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8478 3720 8484 3732
rect 8439 3692 8484 3720
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 9398 3720 9404 3732
rect 8812 3692 9404 3720
rect 8812 3680 8818 3692
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10597 3723 10655 3729
rect 10597 3720 10609 3723
rect 9916 3692 10609 3720
rect 9916 3680 9922 3692
rect 10597 3689 10609 3692
rect 10643 3689 10655 3723
rect 12802 3720 12808 3732
rect 12763 3692 12808 3720
rect 10597 3683 10655 3689
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 13354 3720 13360 3732
rect 13315 3692 13360 3720
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 13955 3692 15516 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 3881 3655 3939 3661
rect 3881 3621 3893 3655
rect 3927 3652 3939 3655
rect 4982 3652 4988 3664
rect 3927 3624 4988 3652
rect 3927 3621 3939 3624
rect 3881 3615 3939 3621
rect 4982 3612 4988 3624
rect 5040 3612 5046 3664
rect 5166 3612 5172 3664
rect 5224 3652 5230 3664
rect 5582 3655 5640 3661
rect 5582 3652 5594 3655
rect 5224 3624 5594 3652
rect 5224 3612 5230 3624
rect 5582 3621 5594 3624
rect 5628 3621 5640 3655
rect 7190 3652 7196 3664
rect 7103 3624 7196 3652
rect 5582 3615 5640 3621
rect 7190 3612 7196 3624
rect 7248 3652 7254 3664
rect 7834 3652 7840 3664
rect 7248 3624 7840 3652
rect 7248 3612 7254 3624
rect 7834 3612 7840 3624
rect 7892 3612 7898 3664
rect 10042 3661 10048 3664
rect 10039 3652 10048 3661
rect 10003 3624 10048 3652
rect 10039 3615 10048 3624
rect 10042 3612 10048 3615
rect 10100 3612 10106 3664
rect 11514 3652 11520 3664
rect 11475 3624 11520 3652
rect 11514 3612 11520 3624
rect 11572 3612 11578 3664
rect 11606 3612 11612 3664
rect 11664 3652 11670 3664
rect 12529 3655 12587 3661
rect 11664 3624 11709 3652
rect 11664 3612 11670 3624
rect 12529 3621 12541 3655
rect 12575 3652 12587 3655
rect 12986 3652 12992 3664
rect 12575 3624 12992 3652
rect 12575 3621 12587 3624
rect 12529 3615 12587 3621
rect 12986 3612 12992 3624
rect 13044 3612 13050 3664
rect 15488 3661 15516 3692
rect 15746 3680 15752 3732
rect 15804 3720 15810 3732
rect 15804 3692 19104 3720
rect 15804 3680 15810 3692
rect 15473 3655 15531 3661
rect 15473 3621 15485 3655
rect 15519 3652 15531 3655
rect 15654 3652 15660 3664
rect 15519 3624 15660 3652
rect 15519 3621 15531 3624
rect 15473 3615 15531 3621
rect 15654 3612 15660 3624
rect 15712 3652 15718 3664
rect 15712 3624 16068 3652
rect 15712 3612 15718 3624
rect 1302 3544 1308 3596
rect 1360 3584 1366 3596
rect 1432 3587 1490 3593
rect 1432 3584 1444 3587
rect 1360 3556 1444 3584
rect 1360 3544 1366 3556
rect 1432 3553 1444 3556
rect 1478 3553 1490 3587
rect 1432 3547 1490 3553
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 2222 3584 2228 3596
rect 1636 3556 2228 3584
rect 1636 3544 1642 3556
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 3050 3584 3056 3596
rect 3011 3556 3056 3584
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 4132 3587 4190 3593
rect 4132 3553 4144 3587
rect 4178 3584 4190 3587
rect 4522 3584 4528 3596
rect 4178 3556 4528 3584
rect 4178 3553 4190 3556
rect 4132 3547 4190 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 6181 3587 6239 3593
rect 6181 3584 6193 3587
rect 4764 3556 6193 3584
rect 4764 3544 4770 3556
rect 6181 3553 6193 3556
rect 6227 3584 6239 3587
rect 6546 3584 6552 3596
rect 6227 3556 6552 3584
rect 6227 3553 6239 3556
rect 6181 3547 6239 3553
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 8570 3584 8576 3596
rect 8531 3556 8576 3584
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 16040 3584 16068 3624
rect 16298 3612 16304 3664
rect 16356 3652 16362 3664
rect 18417 3655 18475 3661
rect 18417 3652 18429 3655
rect 16356 3624 18429 3652
rect 16356 3612 16362 3624
rect 18417 3621 18429 3624
rect 18463 3621 18475 3655
rect 18417 3615 18475 3621
rect 19076 3596 19104 3692
rect 16945 3587 17003 3593
rect 16945 3584 16957 3587
rect 16040 3556 16957 3584
rect 16945 3553 16957 3556
rect 16991 3584 17003 3587
rect 17310 3584 17316 3596
rect 16991 3556 17316 3584
rect 16991 3553 17003 3556
rect 16945 3547 17003 3553
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 19058 3584 19064 3596
rect 19019 3556 19064 3584
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 4890 3516 4896 3528
rect 3191 3488 4896 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5258 3516 5264 3528
rect 5171 3488 5264 3516
rect 5258 3476 5264 3488
rect 5316 3516 5322 3528
rect 6638 3516 6644 3528
rect 5316 3488 6644 3516
rect 5316 3476 5322 3488
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 7098 3516 7104 3528
rect 7059 3488 7104 3516
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 7558 3516 7564 3528
rect 7519 3488 7564 3516
rect 7558 3476 7564 3488
rect 7616 3476 7622 3528
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 8904 3488 9689 3516
rect 8904 3476 8910 3488
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 11793 3519 11851 3525
rect 11793 3516 11805 3519
rect 9677 3479 9735 3485
rect 11624 3488 11805 3516
rect 1535 3451 1593 3457
rect 1535 3417 1547 3451
rect 1581 3448 1593 3451
rect 1581 3420 4016 3448
rect 1581 3417 1593 3420
rect 1535 3411 1593 3417
rect 3988 3380 4016 3420
rect 4338 3408 4344 3460
rect 4396 3448 4402 3460
rect 4617 3451 4675 3457
rect 4617 3448 4629 3451
rect 4396 3420 4629 3448
rect 4396 3408 4402 3420
rect 4617 3417 4629 3420
rect 4663 3417 4675 3451
rect 4617 3411 4675 3417
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 11333 3451 11391 3457
rect 11333 3448 11345 3451
rect 11296 3420 11345 3448
rect 11296 3408 11302 3420
rect 11333 3417 11345 3420
rect 11379 3448 11391 3451
rect 11624 3448 11652 3488
rect 11793 3485 11805 3488
rect 11839 3485 11851 3519
rect 12986 3516 12992 3528
rect 12947 3488 12992 3516
rect 11793 3479 11851 3485
rect 12986 3476 12992 3488
rect 13044 3516 13050 3528
rect 14274 3516 14280 3528
rect 13044 3488 14280 3516
rect 13044 3476 13050 3488
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 15378 3516 15384 3528
rect 15339 3488 15384 3516
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 15470 3476 15476 3528
rect 15528 3516 15534 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 15528 3488 16865 3516
rect 15528 3476 15534 3488
rect 16853 3485 16865 3488
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 11379 3420 11652 3448
rect 11379 3417 11391 3420
rect 11333 3411 11391 3417
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 15933 3451 15991 3457
rect 15933 3448 15945 3451
rect 14884 3420 15945 3448
rect 14884 3408 14890 3420
rect 15933 3417 15945 3420
rect 15979 3417 15991 3451
rect 15933 3411 15991 3417
rect 16393 3451 16451 3457
rect 16393 3417 16405 3451
rect 16439 3448 16451 3451
rect 16482 3448 16488 3460
rect 16439 3420 16488 3448
rect 16439 3417 16451 3420
rect 16393 3411 16451 3417
rect 4430 3380 4436 3392
rect 3988 3352 4436 3380
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 6917 3383 6975 3389
rect 6917 3349 6929 3383
rect 6963 3380 6975 3383
rect 7190 3380 7196 3392
rect 6963 3352 7196 3380
rect 6963 3349 6975 3352
rect 6917 3343 6975 3349
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 8478 3340 8484 3392
rect 8536 3380 8542 3392
rect 8711 3383 8769 3389
rect 8711 3380 8723 3383
rect 8536 3352 8723 3380
rect 8536 3340 8542 3352
rect 8711 3349 8723 3352
rect 8757 3380 8769 3383
rect 9033 3383 9091 3389
rect 9033 3380 9045 3383
rect 8757 3352 9045 3380
rect 8757 3349 8769 3352
rect 8711 3343 8769 3349
rect 9033 3349 9045 3352
rect 9079 3349 9091 3383
rect 9033 3343 9091 3349
rect 14645 3383 14703 3389
rect 14645 3349 14657 3383
rect 14691 3380 14703 3383
rect 15746 3380 15752 3392
rect 14691 3352 15752 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 15948 3380 15976 3411
rect 16482 3408 16488 3420
rect 16540 3448 16546 3460
rect 20254 3448 20260 3460
rect 16540 3420 20260 3448
rect 16540 3408 16546 3420
rect 20254 3408 20260 3420
rect 20312 3408 20318 3460
rect 17954 3380 17960 3392
rect 15948 3352 17960 3380
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 18046 3340 18052 3392
rect 18104 3380 18110 3392
rect 19518 3380 19524 3392
rect 18104 3352 19524 3380
rect 18104 3340 18110 3352
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1302 3136 1308 3188
rect 1360 3176 1366 3188
rect 2501 3179 2559 3185
rect 2501 3176 2513 3179
rect 1360 3148 2513 3176
rect 1360 3136 1366 3148
rect 2501 3145 2513 3148
rect 2547 3145 2559 3179
rect 2958 3176 2964 3188
rect 2919 3148 2964 3176
rect 2501 3139 2559 3145
rect 2516 3108 2544 3139
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 4893 3179 4951 3185
rect 4893 3145 4905 3179
rect 4939 3176 4951 3179
rect 5166 3176 5172 3188
rect 4939 3148 5172 3176
rect 4939 3145 4951 3148
rect 4893 3139 4951 3145
rect 5166 3136 5172 3148
rect 5224 3176 5230 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 5224 3148 6193 3176
rect 5224 3136 5230 3148
rect 6181 3145 6193 3148
rect 6227 3176 6239 3179
rect 6270 3176 6276 3188
rect 6227 3148 6276 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 6546 3176 6552 3188
rect 6507 3148 6552 3176
rect 6546 3136 6552 3148
rect 6604 3176 6610 3188
rect 7006 3176 7012 3188
rect 6604 3148 7012 3176
rect 6604 3136 6610 3148
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 7834 3176 7840 3188
rect 7795 3148 7840 3176
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8846 3176 8852 3188
rect 8807 3148 8852 3176
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 8938 3136 8944 3188
rect 8996 3176 9002 3188
rect 9217 3179 9275 3185
rect 9217 3176 9229 3179
rect 8996 3148 9229 3176
rect 8996 3136 9002 3148
rect 9217 3145 9229 3148
rect 9263 3176 9275 3179
rect 11054 3176 11060 3188
rect 9263 3148 9674 3176
rect 11015 3148 11060 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 4338 3108 4344 3120
rect 2516 3080 4344 3108
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 4522 3108 4528 3120
rect 4435 3080 4528 3108
rect 4522 3068 4528 3080
rect 4580 3108 4586 3120
rect 5994 3108 6000 3120
rect 4580 3080 6000 3108
rect 4580 3068 4586 3080
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 7098 3068 7104 3120
rect 7156 3108 7162 3120
rect 8205 3111 8263 3117
rect 8205 3108 8217 3111
rect 7156 3080 8217 3108
rect 7156 3068 7162 3080
rect 8205 3077 8217 3080
rect 8251 3077 8263 3111
rect 8205 3071 8263 3077
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2130 3040 2136 3052
rect 1903 3012 2136 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3040 4215 3043
rect 5258 3040 5264 3052
rect 4203 3012 5264 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 6362 3000 6368 3052
rect 6420 3040 6426 3052
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 6420 3012 8401 3040
rect 6420 3000 6426 3012
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 9398 3040 9404 3052
rect 9359 3012 9404 3040
rect 8389 3003 8447 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 842 2932 848 2984
rect 900 2972 906 2984
rect 1486 2972 1492 2984
rect 900 2944 1492 2972
rect 900 2932 906 2944
rect 1486 2932 1492 2944
rect 1544 2932 1550 2984
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2406 2972 2412 2984
rect 2271 2944 2412 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2941 3571 2975
rect 3878 2972 3884 2984
rect 3839 2944 3884 2972
rect 3513 2935 3571 2941
rect 1854 2864 1860 2916
rect 1912 2904 1918 2916
rect 3237 2907 3295 2913
rect 3237 2904 3249 2907
rect 1912 2876 3249 2904
rect 1912 2864 1918 2876
rect 3237 2873 3249 2876
rect 3283 2904 3295 2907
rect 3528 2904 3556 2935
rect 3878 2932 3884 2944
rect 3936 2972 3942 2984
rect 4982 2972 4988 2984
rect 3936 2944 4154 2972
rect 4943 2944 4988 2972
rect 3936 2932 3942 2944
rect 3283 2876 3556 2904
rect 4126 2904 4154 2944
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5074 2904 5080 2916
rect 4126 2876 5080 2904
rect 3283 2873 3295 2876
rect 3237 2867 3295 2873
rect 5074 2864 5080 2876
rect 5132 2864 5138 2916
rect 5166 2864 5172 2916
rect 5224 2904 5230 2916
rect 5306 2907 5364 2913
rect 5306 2904 5318 2907
rect 5224 2876 5318 2904
rect 5224 2864 5230 2876
rect 5306 2873 5318 2876
rect 5352 2873 5364 2907
rect 6730 2904 6736 2916
rect 5306 2867 5364 2873
rect 5920 2876 6736 2904
rect 4982 2796 4988 2848
rect 5040 2836 5046 2848
rect 5920 2845 5948 2876
rect 6730 2864 6736 2876
rect 6788 2864 6794 2916
rect 6917 2907 6975 2913
rect 6917 2873 6929 2907
rect 6963 2873 6975 2907
rect 6917 2867 6975 2873
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5040 2808 5917 2836
rect 5040 2796 5046 2808
rect 5905 2805 5917 2808
rect 5951 2805 5963 2839
rect 6932 2836 6960 2867
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 7558 2904 7564 2916
rect 7064 2876 7109 2904
rect 7519 2876 7564 2904
rect 7064 2864 7070 2876
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 9646 2904 9674 3148
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12986 3176 12992 3188
rect 12299 3148 12992 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13081 3179 13139 3185
rect 13081 3145 13093 3179
rect 13127 3176 13139 3179
rect 13354 3176 13360 3188
rect 13127 3148 13360 3176
rect 13127 3145 13139 3148
rect 13081 3139 13139 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 13596 3148 14565 3176
rect 13596 3136 13602 3148
rect 14553 3145 14565 3148
rect 14599 3176 14611 3179
rect 14829 3179 14887 3185
rect 14829 3176 14841 3179
rect 14599 3148 14841 3176
rect 14599 3145 14611 3148
rect 14553 3139 14611 3145
rect 14829 3145 14841 3148
rect 14875 3145 14887 3179
rect 14829 3139 14887 3145
rect 15013 3179 15071 3185
rect 15013 3145 15025 3179
rect 15059 3176 15071 3179
rect 15378 3176 15384 3188
rect 15059 3148 15384 3176
rect 15059 3145 15071 3148
rect 15013 3139 15071 3145
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15654 3176 15660 3188
rect 15615 3148 15660 3176
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16209 3179 16267 3185
rect 16209 3145 16221 3179
rect 16255 3176 16267 3179
rect 16574 3176 16580 3188
rect 16255 3148 16580 3176
rect 16255 3145 16267 3148
rect 16209 3139 16267 3145
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 17310 3176 17316 3188
rect 17271 3148 17316 3176
rect 17310 3136 17316 3148
rect 17368 3136 17374 3188
rect 17402 3136 17408 3188
rect 17460 3176 17466 3188
rect 19751 3179 19809 3185
rect 19751 3176 19763 3179
rect 17460 3148 19763 3176
rect 17460 3136 17466 3148
rect 19751 3145 19763 3148
rect 19797 3145 19809 3179
rect 19751 3139 19809 3145
rect 10321 3111 10379 3117
rect 10321 3077 10333 3111
rect 10367 3108 10379 3111
rect 11606 3108 11612 3120
rect 10367 3080 11612 3108
rect 10367 3077 10379 3080
rect 10321 3071 10379 3077
rect 11606 3068 11612 3080
rect 11664 3068 11670 3120
rect 12710 3068 12716 3120
rect 12768 3108 12774 3120
rect 15289 3111 15347 3117
rect 15289 3108 15301 3111
rect 12768 3080 15301 3108
rect 12768 3068 12774 3080
rect 15289 3077 15301 3080
rect 15335 3077 15347 3111
rect 15396 3108 15424 3136
rect 15396 3080 16712 3108
rect 15289 3071 15347 3077
rect 16684 3052 16712 3080
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 19058 3108 19064 3120
rect 18012 3080 18276 3108
rect 19019 3080 19064 3108
rect 18012 3068 18018 3080
rect 14734 3040 14740 3052
rect 13372 3012 14740 3040
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 13372 2981 13400 3012
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 16393 3043 16451 3049
rect 16393 3009 16405 3043
rect 16439 3040 16451 3043
rect 16482 3040 16488 3052
rect 16439 3012 16488 3040
rect 16439 3009 16451 3012
rect 16393 3003 16451 3009
rect 16482 3000 16488 3012
rect 16540 3000 16546 3052
rect 16666 3040 16672 3052
rect 16579 3012 16672 3040
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 17034 3000 17040 3052
rect 17092 3040 17098 3052
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17092 3012 18061 3040
rect 17092 3000 17098 3012
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 11149 2975 11207 2981
rect 11149 2972 11161 2975
rect 11112 2944 11161 2972
rect 11112 2932 11118 2944
rect 11149 2941 11161 2944
rect 11195 2941 11207 2975
rect 11149 2935 11207 2941
rect 12713 2975 12771 2981
rect 12713 2941 12725 2975
rect 12759 2972 12771 2975
rect 13357 2975 13415 2981
rect 13357 2972 13369 2975
rect 12759 2944 13369 2972
rect 12759 2941 12771 2944
rect 12713 2935 12771 2941
rect 13357 2941 13369 2944
rect 13403 2941 13415 2975
rect 13357 2935 13415 2941
rect 14829 2975 14887 2981
rect 14829 2941 14841 2975
rect 14875 2972 14887 2975
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 14875 2944 15117 2972
rect 14875 2941 14887 2944
rect 14829 2935 14887 2941
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 18141 2975 18199 2981
rect 18141 2941 18153 2975
rect 18187 2941 18199 2975
rect 18248 2972 18276 3080
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 19648 2975 19706 2981
rect 19648 2972 19660 2975
rect 18248 2944 19660 2972
rect 18141 2935 18199 2941
rect 19648 2941 19660 2944
rect 19694 2972 19706 2975
rect 20073 2975 20131 2981
rect 20073 2972 20085 2975
rect 19694 2944 20085 2972
rect 19694 2941 19706 2944
rect 19648 2935 19706 2941
rect 20073 2941 20085 2944
rect 20119 2941 20131 2975
rect 20073 2935 20131 2941
rect 20692 2975 20750 2981
rect 20692 2941 20704 2975
rect 20738 2972 20750 2975
rect 24372 2975 24430 2981
rect 20738 2944 21220 2972
rect 20738 2941 20750 2944
rect 20692 2935 20750 2941
rect 9722 2907 9780 2913
rect 9722 2904 9734 2907
rect 9646 2876 9734 2904
rect 9722 2873 9734 2876
rect 9768 2904 9780 2907
rect 9950 2904 9956 2916
rect 9768 2876 9956 2904
rect 9768 2873 9780 2876
rect 9722 2867 9780 2873
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 13446 2864 13452 2916
rect 13504 2904 13510 2916
rect 13678 2907 13736 2913
rect 13678 2904 13690 2907
rect 13504 2876 13690 2904
rect 13504 2864 13510 2876
rect 13678 2873 13690 2876
rect 13724 2873 13736 2907
rect 13678 2867 13736 2873
rect 13786 2876 16344 2904
rect 7190 2836 7196 2848
rect 6932 2808 7196 2836
rect 5905 2799 5963 2805
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 10686 2796 10692 2848
rect 10744 2836 10750 2848
rect 11333 2839 11391 2845
rect 11333 2836 11345 2839
rect 10744 2808 11345 2836
rect 10744 2796 10750 2808
rect 11333 2805 11345 2808
rect 11379 2805 11391 2839
rect 11333 2799 11391 2805
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 11793 2839 11851 2845
rect 11793 2836 11805 2839
rect 11664 2808 11805 2836
rect 11664 2796 11670 2808
rect 11793 2805 11805 2808
rect 11839 2836 11851 2839
rect 13786 2836 13814 2876
rect 11839 2808 13814 2836
rect 14277 2839 14335 2845
rect 11839 2805 11851 2808
rect 11793 2799 11851 2805
rect 14277 2805 14289 2839
rect 14323 2836 14335 2839
rect 15930 2836 15936 2848
rect 14323 2808 15936 2836
rect 14323 2805 14335 2808
rect 14277 2799 14335 2805
rect 15930 2796 15936 2808
rect 15988 2796 15994 2848
rect 16316 2836 16344 2876
rect 16482 2864 16488 2916
rect 16540 2904 16546 2916
rect 17773 2907 17831 2913
rect 17773 2904 17785 2907
rect 16540 2876 16585 2904
rect 17144 2876 17785 2904
rect 16540 2864 16546 2876
rect 17144 2836 17172 2876
rect 17773 2873 17785 2876
rect 17819 2904 17831 2907
rect 18156 2904 18184 2935
rect 21192 2913 21220 2944
rect 24372 2941 24384 2975
rect 24418 2972 24430 2975
rect 24418 2944 24900 2972
rect 24418 2941 24430 2944
rect 24372 2935 24430 2941
rect 17819 2876 18184 2904
rect 21177 2907 21235 2913
rect 17819 2873 17831 2876
rect 17773 2867 17831 2873
rect 21177 2873 21189 2907
rect 21223 2904 21235 2907
rect 23842 2904 23848 2916
rect 21223 2876 23848 2904
rect 21223 2873 21235 2876
rect 21177 2867 21235 2873
rect 23842 2864 23848 2876
rect 23900 2864 23906 2916
rect 16316 2808 17172 2836
rect 20162 2796 20168 2848
rect 20220 2836 20226 2848
rect 20763 2839 20821 2845
rect 20763 2836 20775 2839
rect 20220 2808 20775 2836
rect 20220 2796 20226 2808
rect 20763 2805 20775 2808
rect 20809 2805 20821 2839
rect 20763 2799 20821 2805
rect 20898 2796 20904 2848
rect 20956 2836 20962 2848
rect 24872 2845 24900 2944
rect 24443 2839 24501 2845
rect 24443 2836 24455 2839
rect 20956 2808 24455 2836
rect 20956 2796 20962 2808
rect 24443 2805 24455 2808
rect 24489 2805 24501 2839
rect 24443 2799 24501 2805
rect 24857 2839 24915 2845
rect 24857 2805 24869 2839
rect 24903 2836 24915 2839
rect 25958 2836 25964 2848
rect 24903 2808 25964 2836
rect 24903 2805 24915 2808
rect 24857 2799 24915 2805
rect 25958 2796 25964 2808
rect 26016 2796 26022 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1535 2635 1593 2641
rect 1535 2601 1547 2635
rect 1581 2632 1593 2635
rect 3418 2632 3424 2644
rect 1581 2604 3424 2632
rect 1581 2601 1593 2604
rect 1535 2595 1593 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 3878 2632 3884 2644
rect 3559 2604 3884 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 4522 2632 4528 2644
rect 4483 2604 4528 2632
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 5350 2592 5356 2644
rect 5408 2632 5414 2644
rect 6362 2632 6368 2644
rect 5408 2604 6368 2632
rect 5408 2592 5414 2604
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 6638 2632 6644 2644
rect 6599 2604 6644 2632
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 7558 2632 7564 2644
rect 7024 2604 7564 2632
rect 4982 2564 4988 2576
rect 3804 2536 4988 2564
rect 3804 2505 3832 2536
rect 4982 2524 4988 2536
rect 5040 2524 5046 2576
rect 7024 2573 7052 2604
rect 7558 2592 7564 2604
rect 7616 2632 7622 2644
rect 8297 2635 8355 2641
rect 8297 2632 8309 2635
rect 7616 2604 8309 2632
rect 7616 2592 7622 2604
rect 8297 2601 8309 2604
rect 8343 2601 8355 2635
rect 9490 2632 9496 2644
rect 9451 2604 9496 2632
rect 8297 2595 8355 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 9950 2632 9956 2644
rect 9911 2604 9956 2632
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 12342 2632 12348 2644
rect 12303 2604 12348 2632
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 13354 2632 13360 2644
rect 13315 2604 13360 2632
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 15930 2632 15936 2644
rect 15891 2604 15936 2632
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 16206 2592 16212 2644
rect 16264 2632 16270 2644
rect 18049 2635 18107 2641
rect 18049 2632 18061 2635
rect 16264 2604 18061 2632
rect 16264 2592 16270 2604
rect 5445 2567 5503 2573
rect 5445 2564 5457 2567
rect 5092 2536 5457 2564
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2496 1522 2499
rect 3053 2499 3111 2505
rect 1510 2468 2360 2496
rect 1510 2465 1522 2468
rect 1464 2459 1522 2465
rect 2332 2369 2360 2468
rect 3053 2465 3065 2499
rect 3099 2496 3111 2499
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 3099 2468 3801 2496
rect 3099 2465 3111 2468
rect 3053 2459 3111 2465
rect 3789 2465 3801 2468
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 4316 2499 4374 2505
rect 4316 2465 4328 2499
rect 4362 2496 4374 2499
rect 4798 2496 4804 2508
rect 4362 2468 4804 2496
rect 4362 2465 4374 2468
rect 4316 2459 4374 2465
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 5092 2437 5120 2536
rect 5445 2533 5457 2536
rect 5491 2533 5503 2567
rect 5445 2527 5503 2533
rect 7009 2567 7067 2573
rect 7009 2533 7021 2567
rect 7055 2533 7067 2567
rect 7009 2527 7067 2533
rect 7098 2524 7104 2576
rect 7156 2564 7162 2576
rect 7929 2567 7987 2573
rect 7929 2564 7941 2567
rect 7156 2536 7941 2564
rect 7156 2524 7162 2536
rect 7929 2533 7941 2536
rect 7975 2533 7987 2567
rect 9508 2564 9536 2592
rect 10505 2567 10563 2573
rect 10505 2564 10517 2567
rect 9508 2536 10517 2564
rect 7929 2527 7987 2533
rect 10505 2533 10517 2536
rect 10551 2533 10563 2567
rect 10505 2527 10563 2533
rect 11057 2567 11115 2573
rect 11057 2533 11069 2567
rect 11103 2564 11115 2567
rect 11514 2564 11520 2576
rect 11103 2536 11520 2564
rect 11103 2533 11115 2536
rect 11057 2527 11115 2533
rect 11514 2524 11520 2536
rect 11572 2564 11578 2576
rect 11701 2567 11759 2573
rect 11701 2564 11713 2567
rect 11572 2536 11713 2564
rect 11572 2524 11578 2536
rect 11701 2533 11713 2536
rect 11747 2533 11759 2567
rect 11701 2527 11759 2533
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 12360 2496 12388 2592
rect 14001 2567 14059 2573
rect 14001 2533 14013 2567
rect 14047 2564 14059 2567
rect 14921 2567 14979 2573
rect 14921 2564 14933 2567
rect 14047 2536 14933 2564
rect 14047 2533 14059 2536
rect 14001 2527 14059 2533
rect 14921 2533 14933 2536
rect 14967 2564 14979 2567
rect 15470 2564 15476 2576
rect 14967 2536 15476 2564
rect 14967 2533 14979 2536
rect 14921 2527 14979 2533
rect 15470 2524 15476 2536
rect 15528 2524 15534 2576
rect 16316 2573 16344 2604
rect 18049 2601 18061 2604
rect 18095 2632 18107 2635
rect 20162 2632 20168 2644
rect 18095 2604 18460 2632
rect 18095 2601 18107 2604
rect 18049 2595 18107 2601
rect 16301 2567 16359 2573
rect 16301 2533 16313 2567
rect 16347 2533 16359 2567
rect 16301 2527 16359 2533
rect 16574 2524 16580 2576
rect 16632 2564 16638 2576
rect 18325 2567 18383 2573
rect 18325 2564 18337 2567
rect 16632 2536 18337 2564
rect 16632 2524 16638 2536
rect 18325 2533 18337 2536
rect 18371 2533 18383 2567
rect 18325 2527 18383 2533
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12360 2468 12633 2496
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 14553 2499 14611 2505
rect 14553 2465 14565 2499
rect 14599 2496 14611 2499
rect 14826 2496 14832 2508
rect 14599 2468 14832 2496
rect 14599 2465 14611 2468
rect 14553 2459 14611 2465
rect 14826 2456 14832 2468
rect 14884 2456 14890 2508
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2496 15347 2499
rect 15562 2496 15568 2508
rect 15335 2468 15568 2496
rect 15335 2465 15347 2468
rect 15289 2459 15347 2465
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2428 3203 2431
rect 5077 2431 5135 2437
rect 5077 2428 5089 2431
rect 3191 2400 5089 2428
rect 3191 2397 3203 2400
rect 3145 2391 3203 2397
rect 5077 2397 5089 2400
rect 5123 2397 5135 2431
rect 5350 2428 5356 2440
rect 5311 2400 5356 2428
rect 5077 2391 5135 2397
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 10413 2431 10471 2437
rect 5828 2400 6960 2428
rect 2317 2363 2375 2369
rect 2317 2329 2329 2363
rect 2363 2360 2375 2363
rect 5828 2360 5856 2400
rect 2363 2332 5856 2360
rect 6932 2360 6960 2400
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 11425 2431 11483 2437
rect 11425 2428 11437 2431
rect 10459 2400 11437 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 11425 2397 11437 2400
rect 11471 2428 11483 2431
rect 13909 2431 13967 2437
rect 11471 2400 13814 2428
rect 11471 2397 11483 2400
rect 11425 2391 11483 2397
rect 7282 2360 7288 2372
rect 6932 2332 7288 2360
rect 2363 2329 2375 2332
rect 2317 2323 2375 2329
rect 7282 2320 7288 2332
rect 7340 2320 7346 2372
rect 7561 2363 7619 2369
rect 7561 2329 7573 2363
rect 7607 2329 7619 2363
rect 7561 2323 7619 2329
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 9214 2360 9220 2372
rect 8711 2332 9220 2360
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 1949 2295 2007 2301
rect 1949 2261 1961 2295
rect 1995 2292 2007 2295
rect 2406 2292 2412 2304
rect 1995 2264 2412 2292
rect 1995 2261 2007 2264
rect 1949 2255 2007 2261
rect 2406 2252 2412 2264
rect 2464 2252 2470 2304
rect 4798 2292 4804 2304
rect 4759 2264 4804 2292
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 6089 2295 6147 2301
rect 6089 2261 6101 2295
rect 6135 2292 6147 2295
rect 7576 2292 7604 2323
rect 9214 2320 9220 2332
rect 9272 2320 9278 2372
rect 11606 2320 11612 2372
rect 11664 2360 11670 2372
rect 12805 2363 12863 2369
rect 12805 2360 12817 2363
rect 11664 2332 12817 2360
rect 11664 2320 11670 2332
rect 12805 2329 12817 2332
rect 12851 2329 12863 2363
rect 12805 2323 12863 2329
rect 8570 2292 8576 2304
rect 6135 2264 8576 2292
rect 6135 2261 6147 2264
rect 6089 2255 6147 2261
rect 8570 2252 8576 2264
rect 8628 2292 8634 2304
rect 9033 2295 9091 2301
rect 9033 2292 9045 2295
rect 8628 2264 9045 2292
rect 8628 2252 8634 2264
rect 9033 2261 9045 2264
rect 9079 2261 9091 2295
rect 13786 2292 13814 2400
rect 13909 2397 13921 2431
rect 13955 2428 13967 2431
rect 15304 2428 15332 2459
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 18432 2505 18460 2604
rect 18524 2604 20168 2632
rect 18417 2499 18475 2505
rect 18417 2465 18429 2499
rect 18463 2465 18475 2499
rect 18417 2459 18475 2465
rect 13955 2400 15332 2428
rect 16209 2431 16267 2437
rect 13955 2397 13967 2400
rect 13909 2391 13967 2397
rect 16209 2397 16221 2431
rect 16255 2397 16267 2431
rect 16666 2428 16672 2440
rect 16627 2400 16672 2428
rect 16209 2391 16267 2397
rect 16224 2360 16252 2391
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2428 17279 2431
rect 18524 2428 18552 2604
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 20254 2592 20260 2644
rect 20312 2632 20318 2644
rect 21315 2635 21373 2641
rect 21315 2632 21327 2635
rect 20312 2604 21327 2632
rect 20312 2592 20318 2604
rect 21315 2601 21327 2604
rect 21361 2601 21373 2635
rect 21315 2595 21373 2601
rect 23477 2567 23535 2573
rect 23477 2564 23489 2567
rect 23007 2536 23489 2564
rect 19518 2456 19524 2508
rect 19576 2496 19582 2508
rect 23007 2505 23035 2536
rect 23477 2533 23489 2536
rect 23523 2564 23535 2567
rect 24854 2564 24860 2576
rect 23523 2536 24860 2564
rect 23523 2533 23535 2536
rect 23477 2527 23535 2533
rect 24854 2524 24860 2536
rect 24912 2524 24918 2576
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19576 2468 19901 2496
rect 19576 2456 19582 2468
rect 19889 2465 19901 2468
rect 19935 2496 19947 2499
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 19935 2468 20453 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 20441 2459 20499 2465
rect 21244 2499 21302 2505
rect 21244 2465 21256 2499
rect 21290 2465 21302 2499
rect 21244 2459 21302 2465
rect 22992 2499 23050 2505
rect 22992 2465 23004 2499
rect 23038 2465 23050 2499
rect 22992 2459 23050 2465
rect 24648 2499 24706 2505
rect 24648 2465 24660 2499
rect 24694 2496 24706 2499
rect 24694 2468 25176 2496
rect 24694 2465 24706 2468
rect 24648 2459 24706 2465
rect 17267 2400 18552 2428
rect 17267 2397 17279 2400
rect 17221 2391 17279 2397
rect 17236 2360 17264 2391
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 21259 2428 21287 2459
rect 21637 2431 21695 2437
rect 21637 2428 21649 2431
rect 18748 2400 21649 2428
rect 18748 2388 18754 2400
rect 21637 2397 21649 2400
rect 21683 2397 21695 2431
rect 21637 2391 21695 2397
rect 24719 2363 24777 2369
rect 24719 2360 24731 2363
rect 16224 2332 17264 2360
rect 23446 2332 24731 2360
rect 17494 2292 17500 2304
rect 13786 2264 17500 2292
rect 9033 2255 9091 2261
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 19702 2252 19708 2304
rect 19760 2292 19766 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 19760 2264 20085 2292
rect 19760 2252 19766 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 21450 2252 21456 2304
rect 21508 2292 21514 2304
rect 23063 2295 23121 2301
rect 23063 2292 23075 2295
rect 21508 2264 23075 2292
rect 21508 2252 21514 2264
rect 23063 2261 23075 2264
rect 23109 2261 23121 2295
rect 23063 2255 23121 2261
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 23446 2292 23474 2332
rect 24719 2329 24731 2332
rect 24765 2329 24777 2363
rect 24719 2323 24777 2329
rect 25148 2301 25176 2468
rect 23256 2264 23474 2292
rect 25133 2295 25191 2301
rect 23256 2252 23262 2264
rect 25133 2261 25145 2295
rect 25179 2292 25191 2295
rect 27062 2292 27068 2304
rect 25179 2264 27068 2292
rect 25179 2261 25191 2264
rect 25133 2255 25191 2261
rect 27062 2252 27068 2264
rect 27120 2252 27126 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 4338 76 4344 128
rect 4396 116 4402 128
rect 8386 116 8392 128
rect 4396 88 8392 116
rect 4396 76 4402 88
rect 8386 76 8392 88
rect 8444 76 8450 128
rect 18874 76 18880 128
rect 18932 116 18938 128
rect 20622 116 20628 128
rect 18932 88 20628 116
rect 18932 76 18938 88
rect 20622 76 20628 88
rect 20680 76 20686 128
<< via1 >>
rect 7748 27480 7800 27532
rect 8852 27480 8904 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 16856 24352 16908 24404
rect 2872 24216 2924 24268
rect 11980 24259 12032 24268
rect 11980 24225 11998 24259
rect 11998 24225 12032 24259
rect 11980 24216 12032 24225
rect 12532 24216 12584 24268
rect 13452 24216 13504 24268
rect 15844 24216 15896 24268
rect 24676 24259 24728 24268
rect 24676 24225 24694 24259
rect 24694 24225 24728 24259
rect 24676 24216 24728 24225
rect 26884 24216 26936 24268
rect 12716 24080 12768 24132
rect 3608 24012 3660 24064
rect 12348 24012 12400 24064
rect 12624 24012 12676 24064
rect 20628 24012 20680 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2872 23851 2924 23860
rect 2872 23817 2881 23851
rect 2881 23817 2915 23851
rect 2915 23817 2924 23851
rect 2872 23808 2924 23817
rect 3148 23851 3200 23860
rect 3148 23817 3157 23851
rect 3157 23817 3191 23851
rect 3191 23817 3200 23851
rect 3148 23808 3200 23817
rect 4804 23851 4856 23860
rect 4804 23817 4813 23851
rect 4813 23817 4847 23851
rect 4847 23817 4856 23851
rect 4804 23808 4856 23817
rect 7012 23851 7064 23860
rect 7012 23817 7021 23851
rect 7021 23817 7055 23851
rect 7055 23817 7064 23851
rect 7012 23808 7064 23817
rect 10876 23808 10928 23860
rect 11980 23851 12032 23860
rect 11980 23817 11989 23851
rect 11989 23817 12023 23851
rect 12023 23817 12032 23851
rect 11980 23808 12032 23817
rect 13452 23851 13504 23860
rect 13452 23817 13461 23851
rect 13461 23817 13495 23851
rect 13495 23817 13504 23851
rect 13452 23808 13504 23817
rect 14832 23808 14884 23860
rect 15844 23851 15896 23860
rect 15844 23817 15853 23851
rect 15853 23817 15887 23851
rect 15887 23817 15896 23851
rect 15844 23808 15896 23817
rect 16488 23808 16540 23860
rect 18880 23808 18932 23860
rect 3424 23740 3476 23792
rect 8300 23672 8352 23724
rect 940 23604 992 23656
rect 1308 23468 1360 23520
rect 4804 23604 4856 23656
rect 7472 23604 7524 23656
rect 12808 23715 12860 23724
rect 12808 23681 12817 23715
rect 12817 23681 12851 23715
rect 12851 23681 12860 23715
rect 12808 23672 12860 23681
rect 10140 23647 10192 23656
rect 10140 23613 10149 23647
rect 10149 23613 10183 23647
rect 10183 23613 10192 23647
rect 10140 23604 10192 23613
rect 16856 23647 16908 23656
rect 16856 23613 16865 23647
rect 16865 23613 16899 23647
rect 16899 23613 16908 23647
rect 16856 23604 16908 23613
rect 20904 23808 20956 23860
rect 22836 23808 22888 23860
rect 24676 23808 24728 23860
rect 25228 23851 25280 23860
rect 25228 23817 25237 23851
rect 25237 23817 25271 23851
rect 25271 23817 25280 23851
rect 25228 23808 25280 23817
rect 24860 23740 24912 23792
rect 25228 23604 25280 23656
rect 4068 23468 4120 23520
rect 8852 23468 8904 23520
rect 12440 23468 12492 23520
rect 12716 23536 12768 23588
rect 14924 23579 14976 23588
rect 14924 23545 14933 23579
rect 14933 23545 14967 23579
rect 14967 23545 14976 23579
rect 14924 23536 14976 23545
rect 15568 23579 15620 23588
rect 14740 23511 14792 23520
rect 14740 23477 14749 23511
rect 14749 23477 14783 23511
rect 14783 23477 14792 23511
rect 15568 23545 15577 23579
rect 15577 23545 15611 23579
rect 15611 23545 15620 23579
rect 15568 23536 15620 23545
rect 14740 23468 14792 23477
rect 20076 23468 20128 23520
rect 22744 23468 22796 23520
rect 24584 23468 24636 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 7472 23264 7524 23316
rect 12256 23264 12308 23316
rect 14924 23307 14976 23316
rect 12624 23196 12676 23248
rect 14924 23273 14933 23307
rect 14933 23273 14967 23307
rect 14967 23273 14976 23307
rect 14924 23264 14976 23273
rect 15476 23239 15528 23248
rect 15476 23205 15485 23239
rect 15485 23205 15519 23239
rect 15519 23205 15528 23239
rect 15476 23196 15528 23205
rect 11612 23128 11664 23180
rect 13084 23060 13136 23112
rect 13268 23103 13320 23112
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 13268 23060 13320 23069
rect 15384 23103 15436 23112
rect 15384 23069 15393 23103
rect 15393 23069 15427 23103
rect 15427 23069 15436 23103
rect 15384 23060 15436 23069
rect 15568 23060 15620 23112
rect 8484 22967 8536 22976
rect 8484 22933 8493 22967
rect 8493 22933 8527 22967
rect 8527 22933 8536 22967
rect 8484 22924 8536 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 13084 22720 13136 22772
rect 14740 22763 14792 22772
rect 14740 22729 14749 22763
rect 14749 22729 14783 22763
rect 14783 22729 14792 22763
rect 14740 22720 14792 22729
rect 15384 22720 15436 22772
rect 20076 22720 20128 22772
rect 12348 22584 12400 22636
rect 12256 22516 12308 22568
rect 2044 22423 2096 22432
rect 2044 22389 2053 22423
rect 2053 22389 2087 22423
rect 2087 22389 2096 22423
rect 2044 22380 2096 22389
rect 7840 22380 7892 22432
rect 8484 22380 8536 22432
rect 13268 22448 13320 22500
rect 14188 22380 14240 22432
rect 15476 22559 15528 22568
rect 15476 22525 15485 22559
rect 15485 22525 15519 22559
rect 15519 22525 15528 22559
rect 15476 22516 15528 22525
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 12440 22108 12492 22160
rect 12532 21972 12584 22024
rect 11428 21904 11480 21956
rect 12808 21972 12860 22024
rect 11612 21879 11664 21888
rect 11612 21845 11621 21879
rect 11621 21845 11655 21879
rect 11655 21845 11664 21879
rect 11612 21836 11664 21845
rect 12072 21836 12124 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 12532 21632 12584 21684
rect 12440 21539 12492 21548
rect 12440 21505 12449 21539
rect 12449 21505 12483 21539
rect 12483 21505 12492 21539
rect 12440 21496 12492 21505
rect 12348 21428 12400 21480
rect 12532 21471 12584 21480
rect 12532 21437 12541 21471
rect 12541 21437 12575 21471
rect 12575 21437 12584 21471
rect 12532 21428 12584 21437
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 11888 20748 11940 20800
rect 12532 20748 12584 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 1768 20340 1820 20392
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 14280 20000 14332 20052
rect 15568 20000 15620 20052
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 1216 19252 1268 19304
rect 25136 19252 25188 19304
rect 1400 19116 1452 19168
rect 22100 19116 22152 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1768 18955 1820 18964
rect 1768 18921 1777 18955
rect 1777 18921 1811 18955
rect 1811 18921 1820 18955
rect 1768 18912 1820 18921
rect 2044 18912 2096 18964
rect 1676 18776 1728 18828
rect 2964 18776 3016 18828
rect 2412 18572 2464 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 10140 18368 10192 18420
rect 2412 18207 2464 18216
rect 2412 18173 2421 18207
rect 2421 18173 2455 18207
rect 2455 18173 2464 18207
rect 2412 18164 2464 18173
rect 10140 18164 10192 18216
rect 3792 18096 3844 18148
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 2964 18071 3016 18080
rect 2964 18037 2973 18071
rect 2973 18037 3007 18071
rect 3007 18037 3016 18071
rect 2964 18028 3016 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 4068 17824 4120 17876
rect 7748 17867 7800 17876
rect 7748 17833 7757 17867
rect 7757 17833 7791 17867
rect 7791 17833 7800 17867
rect 7748 17824 7800 17833
rect 9588 17756 9640 17808
rect 2136 17731 2188 17740
rect 2136 17697 2145 17731
rect 2145 17697 2179 17731
rect 2179 17697 2188 17731
rect 2136 17688 2188 17697
rect 2412 17731 2464 17740
rect 2412 17697 2421 17731
rect 2421 17697 2455 17731
rect 2455 17697 2464 17731
rect 2412 17688 2464 17697
rect 3700 17688 3752 17740
rect 4620 17688 4672 17740
rect 7380 17688 7432 17740
rect 2320 17663 2372 17672
rect 2320 17629 2329 17663
rect 2329 17629 2363 17663
rect 2363 17629 2372 17663
rect 2320 17620 2372 17629
rect 10140 17663 10192 17672
rect 9128 17552 9180 17604
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 11152 17552 11204 17604
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 2688 17484 2740 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 4620 17323 4672 17332
rect 4620 17289 4629 17323
rect 4629 17289 4663 17323
rect 4663 17289 4672 17323
rect 4620 17280 4672 17289
rect 9128 17323 9180 17332
rect 9128 17289 9137 17323
rect 9137 17289 9171 17323
rect 9171 17289 9180 17323
rect 9128 17280 9180 17289
rect 7380 17212 7432 17264
rect 9772 17144 9824 17196
rect 10140 17187 10192 17196
rect 10140 17153 10149 17187
rect 10149 17153 10183 17187
rect 10183 17153 10192 17187
rect 10140 17144 10192 17153
rect 11152 17187 11204 17196
rect 11152 17153 11161 17187
rect 11161 17153 11195 17187
rect 11195 17153 11204 17187
rect 11152 17144 11204 17153
rect 2136 17076 2188 17128
rect 1492 17008 1544 17060
rect 2872 17076 2924 17128
rect 3976 17076 4028 17128
rect 7656 17119 7708 17128
rect 7656 17085 7665 17119
rect 7665 17085 7699 17119
rect 7699 17085 7708 17119
rect 7656 17076 7708 17085
rect 3240 16983 3292 16992
rect 3240 16949 3249 16983
rect 3249 16949 3283 16983
rect 3283 16949 3292 16983
rect 3240 16940 3292 16949
rect 3700 16983 3752 16992
rect 3700 16949 3709 16983
rect 3709 16949 3743 16983
rect 3743 16949 3752 16983
rect 3700 16940 3752 16949
rect 6184 17008 6236 17060
rect 7564 16983 7616 16992
rect 7564 16949 7573 16983
rect 7573 16949 7607 16983
rect 7607 16949 7616 16983
rect 7564 16940 7616 16949
rect 9588 16940 9640 16992
rect 9772 17051 9824 17060
rect 9772 17017 9781 17051
rect 9781 17017 9815 17051
rect 9815 17017 9824 17051
rect 9772 17008 9824 17017
rect 11336 17008 11388 17060
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 3700 16736 3752 16788
rect 7380 16736 7432 16788
rect 9588 16736 9640 16788
rect 7564 16668 7616 16720
rect 9496 16668 9548 16720
rect 10692 16668 10744 16720
rect 1676 16600 1728 16652
rect 3976 16600 4028 16652
rect 4988 16600 5040 16652
rect 6276 16643 6328 16652
rect 6276 16609 6285 16643
rect 6285 16609 6319 16643
rect 6319 16609 6328 16643
rect 6276 16600 6328 16609
rect 11336 16643 11388 16652
rect 11336 16609 11345 16643
rect 11345 16609 11379 16643
rect 11379 16609 11388 16643
rect 11336 16600 11388 16609
rect 1768 16575 1820 16584
rect 1768 16541 1777 16575
rect 1777 16541 1811 16575
rect 1811 16541 1820 16575
rect 1768 16532 1820 16541
rect 5448 16532 5500 16584
rect 6644 16532 6696 16584
rect 8208 16532 8260 16584
rect 9036 16532 9088 16584
rect 7932 16507 7984 16516
rect 7932 16473 7941 16507
rect 7941 16473 7975 16507
rect 7975 16473 7984 16507
rect 7932 16464 7984 16473
rect 2872 16439 2924 16448
rect 2872 16405 2881 16439
rect 2881 16405 2915 16439
rect 2915 16405 2924 16439
rect 2872 16396 2924 16405
rect 3884 16396 3936 16448
rect 4344 16439 4396 16448
rect 4344 16405 4353 16439
rect 4353 16405 4387 16439
rect 4387 16405 4396 16439
rect 4344 16396 4396 16405
rect 5080 16439 5132 16448
rect 5080 16405 5089 16439
rect 5089 16405 5123 16439
rect 5123 16405 5132 16439
rect 5080 16396 5132 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1768 16192 1820 16244
rect 3148 16235 3200 16244
rect 3148 16201 3157 16235
rect 3157 16201 3191 16235
rect 3191 16201 3200 16235
rect 3148 16192 3200 16201
rect 4988 16192 5040 16244
rect 6644 16235 6696 16244
rect 6644 16201 6653 16235
rect 6653 16201 6687 16235
rect 6687 16201 6696 16235
rect 6644 16192 6696 16201
rect 7564 16192 7616 16244
rect 11336 16192 11388 16244
rect 9036 16124 9088 16176
rect 6276 16099 6328 16108
rect 1768 15852 1820 15904
rect 2688 15920 2740 15972
rect 6276 16065 6285 16099
rect 6285 16065 6319 16099
rect 6319 16065 6328 16099
rect 7932 16099 7984 16108
rect 6276 16056 6328 16065
rect 7932 16065 7941 16099
rect 7941 16065 7975 16099
rect 7975 16065 7984 16099
rect 7932 16056 7984 16065
rect 9772 16056 9824 16108
rect 10692 16056 10744 16108
rect 3148 15988 3200 16040
rect 5080 16031 5132 16040
rect 5080 15997 5089 16031
rect 5089 15997 5123 16031
rect 5123 15997 5132 16031
rect 5080 15988 5132 15997
rect 4436 15963 4488 15972
rect 4436 15929 4445 15963
rect 4445 15929 4479 15963
rect 4479 15929 4488 15963
rect 4436 15920 4488 15929
rect 7472 15963 7524 15972
rect 7472 15929 7481 15963
rect 7481 15929 7515 15963
rect 7515 15929 7524 15963
rect 7472 15920 7524 15929
rect 7656 15920 7708 15972
rect 3056 15852 3108 15904
rect 4344 15852 4396 15904
rect 5264 15852 5316 15904
rect 5448 15895 5500 15904
rect 5448 15861 5457 15895
rect 5457 15861 5491 15895
rect 5491 15861 5500 15895
rect 5448 15852 5500 15861
rect 9496 15895 9548 15904
rect 9496 15861 9505 15895
rect 9505 15861 9539 15895
rect 9539 15861 9548 15895
rect 9496 15852 9548 15861
rect 9772 15963 9824 15972
rect 9772 15929 9781 15963
rect 9781 15929 9815 15963
rect 9815 15929 9824 15963
rect 9772 15920 9824 15929
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 8208 15691 8260 15700
rect 8208 15657 8217 15691
rect 8217 15657 8251 15691
rect 8251 15657 8260 15691
rect 8208 15648 8260 15657
rect 1860 15580 1912 15632
rect 6828 15623 6880 15632
rect 6828 15589 6837 15623
rect 6837 15589 6871 15623
rect 6871 15589 6880 15623
rect 6828 15580 6880 15589
rect 7472 15580 7524 15632
rect 9496 15580 9548 15632
rect 4988 15555 5040 15564
rect 4988 15521 4997 15555
rect 4997 15521 5031 15555
rect 5031 15521 5040 15555
rect 4988 15512 5040 15521
rect 9772 15555 9824 15564
rect 9772 15521 9781 15555
rect 9781 15521 9815 15555
rect 9815 15521 9824 15555
rect 9772 15512 9824 15521
rect 11612 15555 11664 15564
rect 11612 15521 11621 15555
rect 11621 15521 11655 15555
rect 11655 15521 11664 15555
rect 11612 15512 11664 15521
rect 1308 15444 1360 15496
rect 3148 15444 3200 15496
rect 6184 15444 6236 15496
rect 10784 15444 10836 15496
rect 2964 15308 3016 15360
rect 3884 15351 3936 15360
rect 3884 15317 3893 15351
rect 3893 15317 3927 15351
rect 3927 15317 3936 15351
rect 3884 15308 3936 15317
rect 4620 15351 4672 15360
rect 4620 15317 4629 15351
rect 4629 15317 4663 15351
rect 4663 15317 4672 15351
rect 4620 15308 4672 15317
rect 7748 15351 7800 15360
rect 7748 15317 7757 15351
rect 7757 15317 7791 15351
rect 7791 15317 7800 15351
rect 7748 15308 7800 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 3148 15147 3200 15156
rect 3148 15113 3157 15147
rect 3157 15113 3191 15147
rect 3191 15113 3200 15147
rect 3148 15104 3200 15113
rect 3608 15147 3660 15156
rect 3608 15113 3617 15147
rect 3617 15113 3651 15147
rect 3651 15113 3660 15147
rect 3608 15104 3660 15113
rect 4436 15104 4488 15156
rect 4988 15104 5040 15156
rect 6184 15147 6236 15156
rect 6184 15113 6193 15147
rect 6193 15113 6227 15147
rect 6227 15113 6236 15147
rect 6184 15104 6236 15113
rect 11612 15147 11664 15156
rect 11612 15113 11621 15147
rect 11621 15113 11655 15147
rect 11655 15113 11664 15147
rect 11612 15104 11664 15113
rect 25136 15147 25188 15156
rect 25136 15113 25145 15147
rect 25145 15113 25179 15147
rect 25179 15113 25188 15147
rect 25136 15104 25188 15113
rect 2688 15079 2740 15088
rect 2688 15045 2697 15079
rect 2697 15045 2731 15079
rect 2731 15045 2740 15079
rect 2688 15036 2740 15045
rect 3056 15036 3108 15088
rect 2964 14968 3016 15020
rect 3608 14968 3660 15020
rect 4712 15011 4764 15020
rect 4712 14977 4721 15011
rect 4721 14977 4755 15011
rect 4755 14977 4764 15011
rect 4712 14968 4764 14977
rect 6828 15036 6880 15088
rect 11244 15079 11296 15088
rect 7472 14968 7524 15020
rect 11244 15045 11253 15079
rect 11253 15045 11287 15079
rect 11287 15045 11296 15079
rect 11244 15036 11296 15045
rect 11152 14968 11204 15020
rect 1676 14832 1728 14884
rect 2228 14875 2280 14884
rect 2228 14841 2237 14875
rect 2237 14841 2271 14875
rect 2271 14841 2280 14875
rect 2228 14832 2280 14841
rect 4436 14832 4488 14884
rect 1860 14807 1912 14816
rect 1860 14773 1869 14807
rect 1869 14773 1903 14807
rect 1903 14773 1912 14807
rect 1860 14764 1912 14773
rect 7748 14832 7800 14884
rect 10784 14875 10836 14884
rect 10784 14841 10793 14875
rect 10793 14841 10827 14875
rect 10827 14841 10836 14875
rect 10784 14832 10836 14841
rect 8208 14764 8260 14816
rect 12256 14832 12308 14884
rect 25136 14900 25188 14952
rect 12164 14807 12216 14816
rect 12164 14773 12173 14807
rect 12173 14773 12207 14807
rect 12207 14773 12216 14807
rect 12164 14764 12216 14773
rect 12532 14807 12584 14816
rect 12532 14773 12541 14807
rect 12541 14773 12575 14807
rect 12575 14773 12584 14807
rect 12532 14764 12584 14773
rect 25136 14764 25188 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 7012 14560 7064 14612
rect 7656 14603 7708 14612
rect 7656 14569 7665 14603
rect 7665 14569 7699 14603
rect 7699 14569 7708 14603
rect 7656 14560 7708 14569
rect 9772 14560 9824 14612
rect 9864 14560 9916 14612
rect 11336 14560 11388 14612
rect 13084 14603 13136 14612
rect 13084 14569 13093 14603
rect 13093 14569 13127 14603
rect 13127 14569 13136 14603
rect 13084 14560 13136 14569
rect 2780 14492 2832 14544
rect 4620 14492 4672 14544
rect 11612 14535 11664 14544
rect 11612 14501 11621 14535
rect 11621 14501 11655 14535
rect 11655 14501 11664 14535
rect 11612 14492 11664 14501
rect 23848 14492 23900 14544
rect 1584 14424 1636 14476
rect 12992 14467 13044 14476
rect 12992 14433 13001 14467
rect 13001 14433 13035 14467
rect 13035 14433 13044 14467
rect 12992 14424 13044 14433
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 2964 14399 3016 14408
rect 2964 14365 2973 14399
rect 2973 14365 3007 14399
rect 3007 14365 3016 14399
rect 2964 14356 3016 14365
rect 4068 14356 4120 14408
rect 4528 14356 4580 14408
rect 8024 14356 8076 14408
rect 9496 14356 9548 14408
rect 11520 14399 11572 14408
rect 11520 14365 11529 14399
rect 11529 14365 11563 14399
rect 11563 14365 11572 14399
rect 11520 14356 11572 14365
rect 14464 14424 14516 14476
rect 11244 14288 11296 14340
rect 1768 14220 1820 14272
rect 2044 14220 2096 14272
rect 4712 14220 4764 14272
rect 6368 14220 6420 14272
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 12256 14220 12308 14272
rect 24860 14356 24912 14408
rect 25136 14288 25188 14340
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 2228 14016 2280 14068
rect 4068 14059 4120 14068
rect 2320 13880 2372 13932
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 4620 14016 4672 14068
rect 7748 14059 7800 14068
rect 7748 14025 7757 14059
rect 7757 14025 7791 14059
rect 7791 14025 7800 14059
rect 7748 14016 7800 14025
rect 8024 14059 8076 14068
rect 8024 14025 8033 14059
rect 8033 14025 8067 14059
rect 8067 14025 8076 14059
rect 8024 14016 8076 14025
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 11612 14016 11664 14068
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 12992 14016 13044 14068
rect 14188 14059 14240 14068
rect 14188 14025 14197 14059
rect 14197 14025 14231 14059
rect 14231 14025 14240 14059
rect 14188 14016 14240 14025
rect 25136 14059 25188 14068
rect 25136 14025 25145 14059
rect 25145 14025 25179 14059
rect 25179 14025 25188 14059
rect 25136 14016 25188 14025
rect 4528 13948 4580 14000
rect 4712 13880 4764 13932
rect 7104 13880 7156 13932
rect 8944 13880 8996 13932
rect 4896 13744 4948 13796
rect 10784 13880 10836 13932
rect 13084 13880 13136 13932
rect 13360 13812 13412 13864
rect 24676 13880 24728 13932
rect 2044 13676 2096 13728
rect 2780 13676 2832 13728
rect 6644 13719 6696 13728
rect 6644 13685 6653 13719
rect 6653 13685 6687 13719
rect 6687 13685 6696 13719
rect 6644 13676 6696 13685
rect 7012 13676 7064 13728
rect 9772 13744 9824 13796
rect 9864 13676 9916 13728
rect 24860 13787 24912 13796
rect 13176 13719 13228 13728
rect 13176 13685 13185 13719
rect 13185 13685 13219 13719
rect 13219 13685 13228 13719
rect 13176 13676 13228 13685
rect 23848 13676 23900 13728
rect 24032 13719 24084 13728
rect 24032 13685 24041 13719
rect 24041 13685 24075 13719
rect 24075 13685 24084 13719
rect 24860 13753 24869 13787
rect 24869 13753 24903 13787
rect 24903 13753 24912 13787
rect 24860 13744 24912 13753
rect 24032 13676 24084 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 4896 13472 4948 13524
rect 8024 13472 8076 13524
rect 9772 13515 9824 13524
rect 9772 13481 9781 13515
rect 9781 13481 9815 13515
rect 9815 13481 9824 13515
rect 9772 13472 9824 13481
rect 10784 13515 10836 13524
rect 10784 13481 10793 13515
rect 10793 13481 10827 13515
rect 10827 13481 10836 13515
rect 10784 13472 10836 13481
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 12256 13515 12308 13524
rect 12256 13481 12265 13515
rect 12265 13481 12299 13515
rect 12299 13481 12308 13515
rect 12256 13472 12308 13481
rect 13360 13515 13412 13524
rect 13360 13481 13369 13515
rect 13369 13481 13403 13515
rect 13403 13481 13412 13515
rect 13360 13472 13412 13481
rect 24032 13515 24084 13524
rect 24032 13481 24041 13515
rect 24041 13481 24075 13515
rect 24075 13481 24084 13515
rect 24032 13472 24084 13481
rect 2044 13404 2096 13456
rect 5080 13404 5132 13456
rect 7748 13379 7800 13388
rect 7748 13345 7757 13379
rect 7757 13345 7791 13379
rect 7791 13345 7800 13379
rect 7748 13336 7800 13345
rect 9680 13379 9732 13388
rect 1952 13268 2004 13320
rect 2596 13268 2648 13320
rect 4344 13268 4396 13320
rect 6184 13268 6236 13320
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 7380 13268 7432 13320
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 9680 13336 9732 13345
rect 8944 13268 8996 13320
rect 12164 13336 12216 13388
rect 13544 13379 13596 13388
rect 13544 13345 13553 13379
rect 13553 13345 13587 13379
rect 13587 13345 13596 13379
rect 13544 13336 13596 13345
rect 23848 13379 23900 13388
rect 23848 13345 23857 13379
rect 23857 13345 23891 13379
rect 23891 13345 23900 13379
rect 23848 13336 23900 13345
rect 2504 13200 2556 13252
rect 2780 13175 2832 13184
rect 2780 13141 2789 13175
rect 2789 13141 2823 13175
rect 2823 13141 2832 13175
rect 2780 13132 2832 13141
rect 3516 13132 3568 13184
rect 7104 13175 7156 13184
rect 7104 13141 7113 13175
rect 7113 13141 7147 13175
rect 7147 13141 7156 13175
rect 7104 13132 7156 13141
rect 9128 13132 9180 13184
rect 9496 13132 9548 13184
rect 11152 13175 11204 13184
rect 11152 13141 11161 13175
rect 11161 13141 11195 13175
rect 11195 13141 11204 13175
rect 11152 13132 11204 13141
rect 14372 13132 14424 13184
rect 24860 13175 24912 13184
rect 24860 13141 24869 13175
rect 24869 13141 24903 13175
rect 24903 13141 24912 13175
rect 24860 13132 24912 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 5172 12928 5224 12980
rect 6276 12928 6328 12980
rect 7748 12928 7800 12980
rect 3792 12860 3844 12912
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 6000 12792 6052 12844
rect 2780 12724 2832 12776
rect 3056 12724 3108 12776
rect 4160 12724 4212 12776
rect 7380 12767 7432 12776
rect 1952 12588 2004 12640
rect 4620 12656 4672 12708
rect 7380 12733 7389 12767
rect 7389 12733 7423 12767
rect 7423 12733 7432 12767
rect 7380 12724 7432 12733
rect 18604 12860 18656 12912
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 12532 12792 12584 12844
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 23848 12835 23900 12844
rect 23848 12801 23857 12835
rect 23857 12801 23891 12835
rect 23891 12801 23900 12835
rect 23848 12792 23900 12801
rect 8944 12767 8996 12776
rect 8944 12733 8953 12767
rect 8953 12733 8987 12767
rect 8987 12733 8996 12767
rect 8944 12724 8996 12733
rect 10968 12767 11020 12776
rect 9680 12699 9732 12708
rect 9680 12665 9689 12699
rect 9689 12665 9723 12699
rect 9723 12665 9732 12699
rect 9680 12656 9732 12665
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 12164 12724 12216 12776
rect 6644 12588 6696 12640
rect 7104 12631 7156 12640
rect 7104 12597 7113 12631
rect 7113 12597 7147 12631
rect 7147 12597 7156 12631
rect 7104 12588 7156 12597
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 11704 12588 11756 12640
rect 12900 12656 12952 12708
rect 13544 12656 13596 12708
rect 14372 12699 14424 12708
rect 14372 12665 14381 12699
rect 14381 12665 14415 12699
rect 14415 12665 14424 12699
rect 14372 12656 14424 12665
rect 15752 12656 15804 12708
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2596 12427 2648 12436
rect 2596 12393 2605 12427
rect 2605 12393 2639 12427
rect 2639 12393 2648 12427
rect 2596 12384 2648 12393
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 5172 12384 5224 12436
rect 10968 12384 11020 12436
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 13176 12427 13228 12436
rect 13176 12393 13185 12427
rect 13185 12393 13219 12427
rect 13219 12393 13228 12427
rect 13176 12384 13228 12393
rect 14280 12384 14332 12436
rect 1676 12291 1728 12300
rect 1676 12257 1685 12291
rect 1685 12257 1719 12291
rect 1719 12257 1728 12291
rect 1676 12248 1728 12257
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 5080 12291 5132 12300
rect 3240 12180 3292 12232
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 6092 12248 6144 12300
rect 7380 12316 7432 12368
rect 8944 12316 8996 12368
rect 8668 12248 8720 12300
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 5448 12180 5500 12232
rect 6552 12223 6604 12232
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 6552 12180 6604 12189
rect 8576 12180 8628 12232
rect 10600 12180 10652 12232
rect 11336 12248 11388 12300
rect 12900 12248 12952 12300
rect 14372 12248 14424 12300
rect 15752 12291 15804 12300
rect 15752 12257 15761 12291
rect 15761 12257 15795 12291
rect 15795 12257 15804 12291
rect 15752 12248 15804 12257
rect 11796 12180 11848 12232
rect 12164 12180 12216 12232
rect 13912 12180 13964 12232
rect 6184 12112 6236 12164
rect 7288 12112 7340 12164
rect 12992 12112 13044 12164
rect 2044 12087 2096 12096
rect 2044 12053 2053 12087
rect 2053 12053 2087 12087
rect 2087 12053 2096 12087
rect 2044 12044 2096 12053
rect 4160 12044 4212 12096
rect 5264 12044 5316 12096
rect 6460 12087 6512 12096
rect 6460 12053 6469 12087
rect 6469 12053 6503 12087
rect 6503 12053 6512 12087
rect 6460 12044 6512 12053
rect 8300 12087 8352 12096
rect 8300 12053 8309 12087
rect 8309 12053 8343 12087
rect 8343 12053 8352 12087
rect 8300 12044 8352 12053
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 3240 11840 3292 11892
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 8576 11883 8628 11892
rect 8576 11849 8585 11883
rect 8585 11849 8619 11883
rect 8619 11849 8628 11883
rect 8576 11840 8628 11849
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 10140 11883 10192 11892
rect 10140 11849 10149 11883
rect 10149 11849 10183 11883
rect 10183 11849 10192 11883
rect 10140 11840 10192 11849
rect 11888 11840 11940 11892
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 15752 11883 15804 11892
rect 15752 11849 15761 11883
rect 15761 11849 15795 11883
rect 15795 11849 15804 11883
rect 15752 11840 15804 11849
rect 24216 11840 24268 11892
rect 1768 11772 1820 11824
rect 7840 11772 7892 11824
rect 8024 11772 8076 11824
rect 12808 11772 12860 11824
rect 14556 11772 14608 11824
rect 3792 11704 3844 11756
rect 7196 11704 7248 11756
rect 10600 11747 10652 11756
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 10600 11704 10652 11713
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 11888 11679 11940 11688
rect 5080 11636 5132 11645
rect 2504 11611 2556 11620
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 2504 11577 2513 11611
rect 2513 11577 2547 11611
rect 2547 11577 2556 11611
rect 2504 11568 2556 11577
rect 11888 11645 11897 11679
rect 11897 11645 11931 11679
rect 11931 11645 11940 11679
rect 11888 11636 11940 11645
rect 14096 11704 14148 11756
rect 1676 11500 1728 11509
rect 2320 11500 2372 11552
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3148 11500 3200 11509
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 5356 11500 5408 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 6092 11500 6144 11552
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 7288 11500 7340 11552
rect 7840 11568 7892 11620
rect 8300 11500 8352 11552
rect 9772 11500 9824 11552
rect 11520 11568 11572 11620
rect 11152 11500 11204 11552
rect 13544 11568 13596 11620
rect 13912 11611 13964 11620
rect 13912 11577 13921 11611
rect 13921 11577 13955 11611
rect 13955 11577 13964 11611
rect 13912 11568 13964 11577
rect 13176 11543 13228 11552
rect 13176 11509 13185 11543
rect 13185 11509 13219 11543
rect 13219 11509 13228 11543
rect 13176 11500 13228 11509
rect 27620 11500 27672 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 3148 11296 3200 11348
rect 4068 11296 4120 11348
rect 7196 11339 7248 11348
rect 7196 11305 7205 11339
rect 7205 11305 7239 11339
rect 7239 11305 7248 11339
rect 7196 11296 7248 11305
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 10968 11296 11020 11348
rect 12808 11296 12860 11348
rect 13084 11296 13136 11348
rect 2044 11228 2096 11280
rect 2504 11271 2556 11280
rect 2504 11237 2513 11271
rect 2513 11237 2547 11271
rect 2547 11237 2556 11271
rect 2504 11228 2556 11237
rect 3976 11160 4028 11212
rect 5264 11160 5316 11212
rect 5908 11228 5960 11280
rect 7472 11271 7524 11280
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 7472 11237 7481 11271
rect 7481 11237 7515 11271
rect 7515 11237 7524 11271
rect 7472 11228 7524 11237
rect 8024 11271 8076 11280
rect 8024 11237 8033 11271
rect 8033 11237 8067 11271
rect 8067 11237 8076 11271
rect 8024 11228 8076 11237
rect 11152 11228 11204 11280
rect 13268 11271 13320 11280
rect 13268 11237 13277 11271
rect 13277 11237 13311 11271
rect 13311 11237 13320 11271
rect 13268 11228 13320 11237
rect 7012 11092 7064 11144
rect 9404 11092 9456 11144
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 9036 11024 9088 11076
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 12716 11024 12768 11076
rect 13176 11024 13228 11076
rect 1676 10999 1728 11008
rect 1676 10965 1685 10999
rect 1685 10965 1719 10999
rect 1719 10965 1728 10999
rect 1676 10956 1728 10965
rect 3700 10956 3752 11008
rect 5356 10956 5408 11008
rect 6460 10999 6512 11008
rect 6460 10965 6469 10999
rect 6469 10965 6503 10999
rect 6503 10965 6512 10999
rect 6460 10956 6512 10965
rect 9772 10956 9824 11008
rect 11244 10999 11296 11008
rect 11244 10965 11253 10999
rect 11253 10965 11287 10999
rect 11287 10965 11296 10999
rect 11244 10956 11296 10965
rect 13084 10999 13136 11008
rect 13084 10965 13093 10999
rect 13093 10965 13127 10999
rect 13127 10965 13136 10999
rect 13084 10956 13136 10965
rect 13820 10956 13872 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1676 10752 1728 10804
rect 3976 10752 4028 10804
rect 11244 10752 11296 10804
rect 14464 10795 14516 10804
rect 6276 10684 6328 10736
rect 8852 10727 8904 10736
rect 8852 10693 8861 10727
rect 8861 10693 8895 10727
rect 8895 10693 8904 10727
rect 8852 10684 8904 10693
rect 9772 10684 9824 10736
rect 14464 10761 14473 10795
rect 14473 10761 14507 10795
rect 14507 10761 14516 10795
rect 14464 10752 14516 10761
rect 13820 10684 13872 10736
rect 14280 10727 14332 10736
rect 14280 10693 14289 10727
rect 14289 10693 14323 10727
rect 14323 10693 14332 10727
rect 14280 10684 14332 10693
rect 2504 10616 2556 10668
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 4804 10616 4856 10668
rect 6460 10616 6512 10668
rect 7656 10616 7708 10668
rect 8576 10616 8628 10668
rect 10048 10616 10100 10668
rect 11428 10616 11480 10668
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 1768 10548 1820 10600
rect 5724 10591 5776 10600
rect 3700 10523 3752 10532
rect 3700 10489 3709 10523
rect 3709 10489 3743 10523
rect 3743 10489 3752 10523
rect 3700 10480 3752 10489
rect 1952 10455 2004 10464
rect 1952 10421 1961 10455
rect 1961 10421 1995 10455
rect 1995 10421 2004 10455
rect 1952 10412 2004 10421
rect 2136 10412 2188 10464
rect 5724 10557 5733 10591
rect 5733 10557 5767 10591
rect 5767 10557 5776 10591
rect 5724 10548 5776 10557
rect 7472 10548 7524 10600
rect 8300 10548 8352 10600
rect 5080 10523 5132 10532
rect 5080 10489 5089 10523
rect 5089 10489 5123 10523
rect 5123 10489 5132 10523
rect 5080 10480 5132 10489
rect 7288 10480 7340 10532
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 10692 10548 10744 10557
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 8576 10523 8628 10532
rect 8576 10489 8585 10523
rect 8585 10489 8619 10523
rect 8619 10489 8628 10523
rect 8576 10480 8628 10489
rect 12532 10523 12584 10532
rect 12532 10489 12541 10523
rect 12541 10489 12575 10523
rect 12575 10489 12584 10523
rect 12532 10480 12584 10489
rect 12624 10523 12676 10532
rect 12624 10489 12633 10523
rect 12633 10489 12667 10523
rect 12667 10489 12676 10523
rect 13176 10523 13228 10532
rect 12624 10480 12676 10489
rect 13176 10489 13185 10523
rect 13185 10489 13219 10523
rect 13219 10489 13228 10523
rect 13176 10480 13228 10489
rect 5264 10412 5316 10464
rect 5448 10412 5500 10464
rect 6184 10412 6236 10464
rect 6644 10455 6696 10464
rect 6644 10421 6653 10455
rect 6653 10421 6687 10455
rect 6687 10421 6696 10455
rect 6644 10412 6696 10421
rect 8024 10455 8076 10464
rect 8024 10421 8033 10455
rect 8033 10421 8067 10455
rect 8067 10421 8076 10455
rect 8024 10412 8076 10421
rect 8852 10412 8904 10464
rect 11152 10412 11204 10464
rect 12716 10412 12768 10464
rect 13728 10480 13780 10532
rect 14004 10523 14056 10532
rect 14004 10489 14013 10523
rect 14013 10489 14047 10523
rect 14047 10489 14056 10523
rect 14004 10480 14056 10489
rect 13636 10412 13688 10464
rect 14372 10412 14424 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2044 10251 2096 10260
rect 2044 10217 2053 10251
rect 2053 10217 2087 10251
rect 2087 10217 2096 10251
rect 2044 10208 2096 10217
rect 2872 10208 2924 10260
rect 3608 10208 3660 10260
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 6000 10208 6052 10260
rect 7656 10251 7708 10260
rect 2136 10072 2188 10124
rect 3884 10140 3936 10192
rect 4252 10183 4304 10192
rect 4252 10149 4261 10183
rect 4261 10149 4295 10183
rect 4295 10149 4304 10183
rect 4252 10140 4304 10149
rect 5080 10140 5132 10192
rect 2688 10047 2740 10056
rect 2688 10013 2697 10047
rect 2697 10013 2731 10047
rect 2731 10013 2740 10047
rect 2688 10004 2740 10013
rect 4436 10004 4488 10056
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 8668 10208 8720 10260
rect 11428 10208 11480 10260
rect 13268 10208 13320 10260
rect 13728 10208 13780 10260
rect 14004 10208 14056 10260
rect 15384 10208 15436 10260
rect 6460 10183 6512 10192
rect 6460 10149 6469 10183
rect 6469 10149 6503 10183
rect 6503 10149 6512 10183
rect 6460 10140 6512 10149
rect 7012 10183 7064 10192
rect 7012 10149 7021 10183
rect 7021 10149 7055 10183
rect 7055 10149 7064 10183
rect 7012 10140 7064 10149
rect 7840 10183 7892 10192
rect 7840 10149 7849 10183
rect 7849 10149 7883 10183
rect 7883 10149 7892 10183
rect 7840 10140 7892 10149
rect 11520 10183 11572 10192
rect 11520 10149 11529 10183
rect 11529 10149 11563 10183
rect 11563 10149 11572 10183
rect 11520 10140 11572 10149
rect 11612 10183 11664 10192
rect 11612 10149 11621 10183
rect 11621 10149 11655 10183
rect 11655 10149 11664 10183
rect 11612 10140 11664 10149
rect 12624 10140 12676 10192
rect 8300 10115 8352 10124
rect 8300 10081 8309 10115
rect 8309 10081 8343 10115
rect 8343 10081 8352 10115
rect 8300 10072 8352 10081
rect 9864 10115 9916 10124
rect 9864 10081 9873 10115
rect 9873 10081 9907 10115
rect 9907 10081 9916 10115
rect 9864 10072 9916 10081
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 13084 10115 13136 10124
rect 13084 10081 13093 10115
rect 13093 10081 13127 10115
rect 13127 10081 13136 10115
rect 13084 10072 13136 10081
rect 13176 10072 13228 10124
rect 15292 10115 15344 10124
rect 15292 10081 15336 10115
rect 15336 10081 15344 10115
rect 15292 10072 15344 10081
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 15568 10004 15620 10056
rect 6276 9936 6328 9988
rect 2044 9868 2096 9920
rect 2596 9911 2648 9920
rect 2596 9877 2605 9911
rect 2605 9877 2639 9911
rect 2639 9877 2648 9911
rect 2596 9868 2648 9877
rect 5356 9911 5408 9920
rect 5356 9877 5365 9911
rect 5365 9877 5399 9911
rect 5399 9877 5408 9911
rect 5356 9868 5408 9877
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9404 9868 9456 9877
rect 10692 9911 10744 9920
rect 10692 9877 10701 9911
rect 10701 9877 10735 9911
rect 10735 9877 10744 9911
rect 10692 9868 10744 9877
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 14464 9868 14516 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2596 9664 2648 9716
rect 3700 9664 3752 9716
rect 4252 9664 4304 9716
rect 4436 9707 4488 9716
rect 4436 9673 4445 9707
rect 4445 9673 4479 9707
rect 4479 9673 4488 9707
rect 4436 9664 4488 9673
rect 9864 9664 9916 9716
rect 10692 9664 10744 9716
rect 11888 9664 11940 9716
rect 12256 9707 12308 9716
rect 12256 9673 12265 9707
rect 12265 9673 12299 9707
rect 12299 9673 12308 9707
rect 12256 9664 12308 9673
rect 13084 9664 13136 9716
rect 15292 9707 15344 9716
rect 15292 9673 15301 9707
rect 15301 9673 15335 9707
rect 15335 9673 15344 9707
rect 15292 9664 15344 9673
rect 8392 9596 8444 9648
rect 8852 9639 8904 9648
rect 8852 9605 8861 9639
rect 8861 9605 8895 9639
rect 8895 9605 8904 9639
rect 8852 9596 8904 9605
rect 10968 9596 11020 9648
rect 13820 9596 13872 9648
rect 14832 9596 14884 9648
rect 1492 9528 1544 9580
rect 3516 9528 3568 9580
rect 6460 9528 6512 9580
rect 7012 9528 7064 9580
rect 8576 9528 8628 9580
rect 10140 9528 10192 9580
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10692 9528 10744 9580
rect 1584 9392 1636 9444
rect 2320 9392 2372 9444
rect 2412 9367 2464 9376
rect 2412 9333 2421 9367
rect 2421 9333 2455 9367
rect 2455 9333 2464 9367
rect 2412 9324 2464 9333
rect 3240 9367 3292 9376
rect 3240 9333 3249 9367
rect 3249 9333 3283 9367
rect 3283 9333 3292 9367
rect 3240 9324 3292 9333
rect 6460 9392 6512 9444
rect 6828 9324 6880 9376
rect 9404 9460 9456 9512
rect 9036 9392 9088 9444
rect 8024 9367 8076 9376
rect 8024 9333 8033 9367
rect 8033 9333 8067 9367
rect 8067 9333 8076 9367
rect 8024 9324 8076 9333
rect 8392 9367 8444 9376
rect 8392 9333 8401 9367
rect 8401 9333 8435 9367
rect 8435 9333 8444 9367
rect 8392 9324 8444 9333
rect 10048 9324 10100 9376
rect 11152 9392 11204 9444
rect 12256 9460 12308 9512
rect 14648 9528 14700 9580
rect 12992 9503 13044 9512
rect 12992 9469 13001 9503
rect 13001 9469 13035 9503
rect 13035 9469 13044 9503
rect 12992 9460 13044 9469
rect 11612 9435 11664 9444
rect 11612 9401 11621 9435
rect 11621 9401 11655 9435
rect 11655 9401 11664 9435
rect 17040 9503 17092 9512
rect 17040 9469 17049 9503
rect 17049 9469 17083 9503
rect 17083 9469 17092 9503
rect 17040 9460 17092 9469
rect 14004 9435 14056 9444
rect 11612 9392 11664 9401
rect 14004 9401 14013 9435
rect 14013 9401 14047 9435
rect 14047 9401 14056 9435
rect 14004 9392 14056 9401
rect 12532 9367 12584 9376
rect 12532 9333 12541 9367
rect 12541 9333 12575 9367
rect 12575 9333 12584 9367
rect 12532 9324 12584 9333
rect 18052 9324 18104 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 3516 9163 3568 9172
rect 3516 9129 3525 9163
rect 3525 9129 3559 9163
rect 3559 9129 3568 9163
rect 3516 9120 3568 9129
rect 4436 9120 4488 9172
rect 4528 9120 4580 9172
rect 6460 9163 6512 9172
rect 6460 9129 6469 9163
rect 6469 9129 6503 9163
rect 6503 9129 6512 9163
rect 6460 9120 6512 9129
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 8300 9163 8352 9172
rect 8300 9129 8309 9163
rect 8309 9129 8343 9163
rect 8343 9129 8352 9163
rect 8300 9120 8352 9129
rect 9036 9163 9088 9172
rect 9036 9129 9045 9163
rect 9045 9129 9079 9163
rect 9079 9129 9088 9163
rect 9036 9120 9088 9129
rect 10140 9120 10192 9172
rect 10692 9163 10744 9172
rect 10692 9129 10701 9163
rect 10701 9129 10735 9163
rect 10735 9129 10744 9163
rect 10692 9120 10744 9129
rect 11520 9120 11572 9172
rect 12716 9163 12768 9172
rect 12716 9129 12725 9163
rect 12725 9129 12759 9163
rect 12759 9129 12768 9163
rect 12716 9120 12768 9129
rect 1952 9095 2004 9104
rect 1952 9061 1961 9095
rect 1961 9061 1995 9095
rect 1995 9061 2004 9095
rect 1952 9052 2004 9061
rect 4896 9052 4948 9104
rect 5264 9027 5316 9036
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 2780 8959 2832 8968
rect 2780 8925 2789 8959
rect 2789 8925 2823 8959
rect 2823 8925 2832 8959
rect 2780 8916 2832 8925
rect 2136 8848 2188 8900
rect 5264 8993 5273 9027
rect 5273 8993 5307 9027
rect 5307 8993 5316 9027
rect 5264 8984 5316 8993
rect 6184 9052 6236 9104
rect 6644 9052 6696 9104
rect 11244 9095 11296 9104
rect 11244 9061 11253 9095
rect 11253 9061 11287 9095
rect 11287 9061 11296 9095
rect 11244 9052 11296 9061
rect 15476 9052 15528 9104
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 2044 8780 2096 8832
rect 3240 8780 3292 8832
rect 4436 8780 4488 8832
rect 5356 8916 5408 8968
rect 11888 8984 11940 9036
rect 12900 9027 12952 9036
rect 12900 8993 12909 9027
rect 12909 8993 12943 9027
rect 12943 8993 12952 9027
rect 12900 8984 12952 8993
rect 12992 8984 13044 9036
rect 13176 8984 13228 9036
rect 13636 8984 13688 9036
rect 7472 8916 7524 8968
rect 10876 8916 10928 8968
rect 11980 8916 12032 8968
rect 15384 8984 15436 9036
rect 16856 8984 16908 9036
rect 16212 8916 16264 8968
rect 11796 8848 11848 8900
rect 15844 8848 15896 8900
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 10140 8780 10192 8832
rect 12992 8780 13044 8832
rect 14832 8780 14884 8832
rect 15752 8823 15804 8832
rect 15752 8789 15761 8823
rect 15761 8789 15795 8823
rect 15795 8789 15804 8823
rect 15752 8780 15804 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2228 8576 2280 8628
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 5264 8576 5316 8628
rect 8484 8576 8536 8628
rect 10140 8619 10192 8628
rect 2504 8551 2556 8560
rect 2504 8517 2513 8551
rect 2513 8517 2547 8551
rect 2547 8517 2556 8551
rect 2504 8508 2556 8517
rect 5448 8508 5500 8560
rect 8300 8508 8352 8560
rect 9772 8551 9824 8560
rect 9772 8517 9781 8551
rect 9781 8517 9815 8551
rect 9815 8517 9824 8551
rect 9772 8508 9824 8517
rect 1952 8440 2004 8492
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 11244 8576 11296 8628
rect 11980 8619 12032 8628
rect 11980 8585 11989 8619
rect 11989 8585 12023 8619
rect 12023 8585 12032 8619
rect 11980 8576 12032 8585
rect 12992 8619 13044 8628
rect 12992 8585 13001 8619
rect 13001 8585 13035 8619
rect 13035 8585 13044 8619
rect 12992 8576 13044 8585
rect 14648 8619 14700 8628
rect 14648 8585 14657 8619
rect 14657 8585 14691 8619
rect 14691 8585 14700 8619
rect 14648 8576 14700 8585
rect 16212 8619 16264 8628
rect 16212 8585 16221 8619
rect 16221 8585 16255 8619
rect 16255 8585 16264 8619
rect 16212 8576 16264 8585
rect 16488 8576 16540 8628
rect 11520 8508 11572 8560
rect 2688 8372 2740 8424
rect 5448 8372 5500 8424
rect 5816 8372 5868 8424
rect 6736 8372 6788 8424
rect 1952 8347 2004 8356
rect 1952 8313 1961 8347
rect 1961 8313 1995 8347
rect 1995 8313 2004 8347
rect 1952 8304 2004 8313
rect 4620 8304 4672 8356
rect 2688 8236 2740 8288
rect 3884 8236 3936 8288
rect 5080 8279 5132 8288
rect 5080 8245 5089 8279
rect 5089 8245 5123 8279
rect 5123 8245 5132 8279
rect 5080 8236 5132 8245
rect 6184 8236 6236 8288
rect 8668 8372 8720 8424
rect 13176 8440 13228 8492
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 10968 8372 11020 8424
rect 11152 8415 11204 8424
rect 11152 8381 11170 8415
rect 11170 8381 11204 8415
rect 11152 8372 11204 8381
rect 11796 8372 11848 8424
rect 14648 8372 14700 8424
rect 15476 8372 15528 8424
rect 8576 8236 8628 8288
rect 11060 8236 11112 8288
rect 12900 8236 12952 8288
rect 13452 8347 13504 8356
rect 13452 8313 13461 8347
rect 13461 8313 13495 8347
rect 13495 8313 13504 8347
rect 13452 8304 13504 8313
rect 22100 8304 22152 8356
rect 13820 8236 13872 8288
rect 14740 8236 14792 8288
rect 15844 8279 15896 8288
rect 15844 8245 15853 8279
rect 15853 8245 15887 8279
rect 15887 8245 15896 8279
rect 15844 8236 15896 8245
rect 16856 8279 16908 8288
rect 16856 8245 16865 8279
rect 16865 8245 16899 8279
rect 16899 8245 16908 8279
rect 16856 8236 16908 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2044 8032 2096 8084
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 5080 8032 5132 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 11152 8075 11204 8084
rect 11152 8041 11161 8075
rect 11161 8041 11195 8075
rect 11195 8041 11204 8075
rect 11152 8032 11204 8041
rect 12256 8032 12308 8084
rect 13820 8032 13872 8084
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 8668 7964 8720 8016
rect 1952 7896 2004 7948
rect 4620 7896 4672 7948
rect 5356 7939 5408 7948
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 5356 7896 5408 7905
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 6552 7939 6604 7948
rect 6552 7905 6561 7939
rect 6561 7905 6595 7939
rect 6595 7905 6604 7939
rect 6552 7896 6604 7905
rect 9864 7939 9916 7948
rect 9864 7905 9873 7939
rect 9873 7905 9907 7939
rect 9907 7905 9916 7939
rect 9864 7896 9916 7905
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 12532 7896 12584 7948
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 15476 7896 15528 7948
rect 17500 7896 17552 7948
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 8576 7828 8628 7880
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 13912 7871 13964 7880
rect 13912 7837 13921 7871
rect 13921 7837 13955 7871
rect 13955 7837 13964 7871
rect 13912 7828 13964 7837
rect 8300 7803 8352 7812
rect 8300 7769 8309 7803
rect 8309 7769 8343 7803
rect 8343 7769 8352 7803
rect 8300 7760 8352 7769
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 1860 7692 1912 7744
rect 7104 7692 7156 7744
rect 8024 7692 8076 7744
rect 8484 7735 8536 7744
rect 8484 7701 8493 7735
rect 8493 7701 8527 7735
rect 8527 7701 8536 7735
rect 8484 7692 8536 7701
rect 11888 7692 11940 7744
rect 13452 7692 13504 7744
rect 14832 7692 14884 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 3424 7488 3476 7540
rect 3056 7352 3108 7404
rect 10508 7488 10560 7540
rect 10968 7488 11020 7540
rect 13912 7488 13964 7540
rect 12256 7420 12308 7472
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 112 7284 164 7336
rect 7748 7327 7800 7336
rect 7748 7293 7757 7327
rect 7757 7293 7791 7327
rect 7791 7293 7800 7327
rect 7748 7284 7800 7293
rect 9128 7284 9180 7336
rect 2872 7216 2924 7268
rect 2044 7148 2096 7200
rect 5356 7216 5408 7268
rect 9220 7216 9272 7268
rect 10048 7352 10100 7404
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 12716 7352 12768 7404
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 16304 7327 16356 7336
rect 3608 7191 3660 7200
rect 3608 7157 3617 7191
rect 3617 7157 3651 7191
rect 3651 7157 3660 7191
rect 3608 7148 3660 7157
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 7104 7148 7156 7200
rect 8576 7191 8628 7200
rect 8576 7157 8585 7191
rect 8585 7157 8619 7191
rect 8619 7157 8628 7191
rect 8576 7148 8628 7157
rect 8852 7191 8904 7200
rect 8852 7157 8861 7191
rect 8861 7157 8895 7191
rect 8895 7157 8904 7191
rect 10968 7259 11020 7268
rect 10968 7225 10977 7259
rect 10977 7225 11011 7259
rect 11011 7225 11020 7259
rect 10968 7216 11020 7225
rect 12256 7216 12308 7268
rect 14372 7259 14424 7268
rect 14372 7225 14381 7259
rect 14381 7225 14415 7259
rect 14415 7225 14424 7259
rect 14372 7216 14424 7225
rect 15292 7216 15344 7268
rect 15568 7216 15620 7268
rect 16304 7293 16313 7327
rect 16313 7293 16347 7327
rect 16347 7293 16356 7327
rect 16304 7284 16356 7293
rect 8852 7148 8904 7157
rect 9864 7148 9916 7200
rect 13360 7191 13412 7200
rect 13360 7157 13369 7191
rect 13369 7157 13403 7191
rect 13403 7157 13412 7191
rect 13360 7148 13412 7157
rect 15844 7191 15896 7200
rect 15844 7157 15853 7191
rect 15853 7157 15887 7191
rect 15887 7157 15896 7191
rect 15844 7148 15896 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 2504 6944 2556 6996
rect 3240 6944 3292 6996
rect 5356 6944 5408 6996
rect 8300 6944 8352 6996
rect 8668 6944 8720 6996
rect 10876 6987 10928 6996
rect 10876 6953 10885 6987
rect 10885 6953 10919 6987
rect 10919 6953 10928 6987
rect 10876 6944 10928 6953
rect 11980 6987 12032 6996
rect 11980 6953 11989 6987
rect 11989 6953 12023 6987
rect 12023 6953 12032 6987
rect 11980 6944 12032 6953
rect 12716 6944 12768 6996
rect 15476 6944 15528 6996
rect 17500 6987 17552 6996
rect 17500 6953 17509 6987
rect 17509 6953 17543 6987
rect 17543 6953 17552 6987
rect 17500 6944 17552 6953
rect 24860 6944 24912 6996
rect 2596 6919 2648 6928
rect 2596 6885 2605 6919
rect 2605 6885 2639 6919
rect 2639 6885 2648 6919
rect 2596 6876 2648 6885
rect 2872 6876 2924 6928
rect 4804 6876 4856 6928
rect 6184 6876 6236 6928
rect 6276 6876 6328 6928
rect 9864 6919 9916 6928
rect 9864 6885 9873 6919
rect 9873 6885 9907 6919
rect 9907 6885 9916 6919
rect 9864 6876 9916 6885
rect 11520 6876 11572 6928
rect 13360 6876 13412 6928
rect 14556 6876 14608 6928
rect 14832 6876 14884 6928
rect 9128 6851 9180 6860
rect 9128 6817 9137 6851
rect 9137 6817 9171 6851
rect 9171 6817 9180 6851
rect 9128 6808 9180 6817
rect 11888 6808 11940 6860
rect 2964 6740 3016 6792
rect 3516 6740 3568 6792
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 9588 6740 9640 6792
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 16856 6851 16908 6860
rect 16856 6817 16865 6851
rect 16865 6817 16899 6851
rect 16899 6817 16908 6851
rect 16856 6808 16908 6817
rect 27620 6876 27672 6928
rect 17316 6808 17368 6860
rect 24676 6851 24728 6860
rect 24676 6817 24678 6851
rect 24678 6817 24728 6851
rect 24676 6808 24728 6817
rect 7288 6715 7340 6724
rect 7288 6681 7297 6715
rect 7297 6681 7331 6715
rect 7331 6681 7340 6715
rect 7288 6672 7340 6681
rect 8668 6672 8720 6724
rect 15292 6672 15344 6724
rect 2044 6604 2096 6656
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 7748 6604 7800 6613
rect 12348 6647 12400 6656
rect 12348 6613 12357 6647
rect 12357 6613 12391 6647
rect 12391 6613 12400 6647
rect 12348 6604 12400 6613
rect 12716 6604 12768 6656
rect 15752 6604 15804 6656
rect 16304 6647 16356 6656
rect 16304 6613 16313 6647
rect 16313 6613 16347 6647
rect 16347 6613 16356 6647
rect 16304 6604 16356 6613
rect 17224 6604 17276 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2964 6443 3016 6452
rect 2964 6409 2973 6443
rect 2973 6409 3007 6443
rect 3007 6409 3016 6443
rect 2964 6400 3016 6409
rect 4712 6400 4764 6452
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 9220 6400 9272 6452
rect 10140 6400 10192 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 12348 6400 12400 6452
rect 13360 6400 13412 6452
rect 4896 6332 4948 6384
rect 6184 6332 6236 6384
rect 2228 6264 2280 6316
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 4804 6307 4856 6316
rect 4804 6273 4813 6307
rect 4813 6273 4847 6307
rect 4847 6273 4856 6307
rect 4804 6264 4856 6273
rect 5540 6264 5592 6316
rect 6736 6264 6788 6316
rect 2320 6196 2372 6248
rect 3608 6128 3660 6180
rect 4804 6128 4856 6180
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 2596 6060 2648 6112
rect 3148 6060 3200 6112
rect 4068 6060 4120 6112
rect 5908 6128 5960 6180
rect 9772 6264 9824 6316
rect 13728 6264 13780 6316
rect 14372 6400 14424 6452
rect 14648 6400 14700 6452
rect 16856 6400 16908 6452
rect 24676 6443 24728 6452
rect 24676 6409 24685 6443
rect 24685 6409 24719 6443
rect 24719 6409 24728 6443
rect 24676 6400 24728 6409
rect 17224 6375 17276 6384
rect 17224 6341 17233 6375
rect 17233 6341 17267 6375
rect 17267 6341 17276 6375
rect 17224 6332 17276 6341
rect 18696 6264 18748 6316
rect 8852 6128 8904 6180
rect 15200 6239 15252 6248
rect 15200 6205 15209 6239
rect 15209 6205 15243 6239
rect 15243 6205 15252 6239
rect 15200 6196 15252 6205
rect 15660 6196 15712 6248
rect 16304 6239 16356 6248
rect 16304 6205 16313 6239
rect 16313 6205 16347 6239
rect 16347 6205 16356 6239
rect 16304 6196 16356 6205
rect 10048 6171 10100 6180
rect 10048 6137 10057 6171
rect 10057 6137 10091 6171
rect 10091 6137 10100 6171
rect 10048 6128 10100 6137
rect 10140 6171 10192 6180
rect 10140 6137 10149 6171
rect 10149 6137 10183 6171
rect 10183 6137 10192 6171
rect 10140 6128 10192 6137
rect 12164 6128 12216 6180
rect 12716 6171 12768 6180
rect 12716 6137 12725 6171
rect 12725 6137 12759 6171
rect 12759 6137 12768 6171
rect 12716 6128 12768 6137
rect 6184 6060 6236 6112
rect 6368 6060 6420 6112
rect 7104 6103 7156 6112
rect 7104 6069 7113 6103
rect 7113 6069 7147 6103
rect 7147 6069 7156 6103
rect 7104 6060 7156 6069
rect 9128 6103 9180 6112
rect 9128 6069 9137 6103
rect 9137 6069 9171 6103
rect 9171 6069 9180 6103
rect 9128 6060 9180 6069
rect 9496 6103 9548 6112
rect 9496 6069 9505 6103
rect 9505 6069 9539 6103
rect 9539 6069 9548 6103
rect 9496 6060 9548 6069
rect 12348 6060 12400 6112
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 19248 6060 19300 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1860 5856 1912 5908
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 2228 5856 2280 5908
rect 3608 5856 3660 5908
rect 5540 5856 5592 5908
rect 6276 5856 6328 5908
rect 6736 5856 6788 5908
rect 7748 5856 7800 5908
rect 1216 5720 1268 5772
rect 3056 5763 3108 5772
rect 3056 5729 3065 5763
rect 3065 5729 3099 5763
rect 3099 5729 3108 5763
rect 5908 5788 5960 5840
rect 6184 5788 6236 5840
rect 9128 5856 9180 5908
rect 9864 5899 9916 5908
rect 9864 5865 9873 5899
rect 9873 5865 9907 5899
rect 9907 5865 9916 5899
rect 9864 5856 9916 5865
rect 13728 5899 13780 5908
rect 13728 5865 13737 5899
rect 13737 5865 13771 5899
rect 13771 5865 13780 5899
rect 13728 5856 13780 5865
rect 14832 5856 14884 5908
rect 15568 5899 15620 5908
rect 15568 5865 15577 5899
rect 15577 5865 15611 5899
rect 15611 5865 15620 5899
rect 15568 5856 15620 5865
rect 16304 5899 16356 5908
rect 16304 5865 16313 5899
rect 16313 5865 16347 5899
rect 16347 5865 16356 5899
rect 16304 5856 16356 5865
rect 17316 5899 17368 5908
rect 17316 5865 17325 5899
rect 17325 5865 17359 5899
rect 17359 5865 17368 5899
rect 17316 5856 17368 5865
rect 9772 5788 9824 5840
rect 12716 5831 12768 5840
rect 12716 5797 12725 5831
rect 12725 5797 12759 5831
rect 12759 5797 12768 5831
rect 12716 5788 12768 5797
rect 12808 5831 12860 5840
rect 12808 5797 12817 5831
rect 12817 5797 12851 5831
rect 12851 5797 12860 5831
rect 12808 5788 12860 5797
rect 4712 5763 4764 5772
rect 3056 5720 3108 5729
rect 4712 5729 4721 5763
rect 4721 5729 4755 5763
rect 4755 5729 4764 5763
rect 4712 5720 4764 5729
rect 7196 5720 7248 5772
rect 9036 5763 9088 5772
rect 9036 5729 9045 5763
rect 9045 5729 9079 5763
rect 9079 5729 9088 5763
rect 9036 5720 9088 5729
rect 11244 5763 11296 5772
rect 11244 5729 11253 5763
rect 11253 5729 11287 5763
rect 11287 5729 11296 5763
rect 11244 5720 11296 5729
rect 11336 5720 11388 5772
rect 14556 5720 14608 5772
rect 15660 5763 15712 5772
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 6000 5652 6052 5704
rect 7840 5652 7892 5704
rect 8760 5652 8812 5704
rect 9772 5652 9824 5704
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 12072 5652 12124 5704
rect 13452 5652 13504 5704
rect 15568 5652 15620 5704
rect 15752 5584 15804 5636
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 10784 5559 10836 5568
rect 10784 5525 10793 5559
rect 10793 5525 10827 5559
rect 10827 5525 10836 5559
rect 10784 5516 10836 5525
rect 12440 5559 12492 5568
rect 12440 5525 12449 5559
rect 12449 5525 12483 5559
rect 12483 5525 12492 5559
rect 12440 5516 12492 5525
rect 12532 5516 12584 5568
rect 14464 5516 14516 5568
rect 22836 5516 22888 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2964 5355 3016 5364
rect 2964 5321 2973 5355
rect 2973 5321 3007 5355
rect 3007 5321 3016 5355
rect 2964 5312 3016 5321
rect 6368 5312 6420 5364
rect 9036 5312 9088 5364
rect 10784 5312 10836 5364
rect 12256 5355 12308 5364
rect 12256 5321 12265 5355
rect 12265 5321 12299 5355
rect 12299 5321 12308 5355
rect 12256 5312 12308 5321
rect 12624 5312 12676 5364
rect 12716 5312 12768 5364
rect 15292 5312 15344 5364
rect 15660 5312 15712 5364
rect 20904 5355 20956 5364
rect 20904 5321 20913 5355
rect 20913 5321 20947 5355
rect 20947 5321 20956 5355
rect 20904 5312 20956 5321
rect 8300 5244 8352 5296
rect 9128 5244 9180 5296
rect 1768 5176 1820 5228
rect 3148 5219 3200 5228
rect 3148 5185 3157 5219
rect 3157 5185 3191 5219
rect 3191 5185 3200 5219
rect 3148 5176 3200 5185
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 7656 5176 7708 5228
rect 9220 5176 9272 5228
rect 1952 5108 2004 5160
rect 2964 5108 3016 5160
rect 3608 5151 3660 5160
rect 3608 5117 3617 5151
rect 3617 5117 3651 5151
rect 3651 5117 3660 5151
rect 3608 5108 3660 5117
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 8944 5108 8996 5160
rect 3056 5040 3108 5092
rect 8300 5040 8352 5092
rect 11336 5108 11388 5160
rect 12440 5219 12492 5228
rect 12440 5185 12449 5219
rect 12449 5185 12483 5219
rect 12483 5185 12492 5219
rect 12440 5176 12492 5185
rect 13360 5244 13412 5296
rect 12900 5176 12952 5228
rect 15476 5176 15528 5228
rect 3608 4972 3660 5024
rect 4712 4972 4764 5024
rect 5356 4972 5408 5024
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 6828 4972 6880 5024
rect 10692 4972 10744 5024
rect 11244 4972 11296 5024
rect 15384 5108 15436 5160
rect 21548 5244 21600 5296
rect 17868 5108 17920 5160
rect 19248 5108 19300 5160
rect 12624 5040 12676 5092
rect 12900 5040 12952 5092
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 14280 5015 14332 5024
rect 14280 4981 14289 5015
rect 14289 4981 14323 5015
rect 14323 4981 14332 5015
rect 14280 4972 14332 4981
rect 18420 4972 18472 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1216 4768 1268 4820
rect 4436 4768 4488 4820
rect 4988 4811 5040 4820
rect 4988 4777 4997 4811
rect 4997 4777 5031 4811
rect 5031 4777 5040 4811
rect 4988 4768 5040 4777
rect 6000 4811 6052 4820
rect 6000 4777 6009 4811
rect 6009 4777 6043 4811
rect 6043 4777 6052 4811
rect 6000 4768 6052 4777
rect 1952 4743 2004 4752
rect 1952 4709 1961 4743
rect 1961 4709 1995 4743
rect 1995 4709 2004 4743
rect 1952 4700 2004 4709
rect 2412 4743 2464 4752
rect 2412 4709 2421 4743
rect 2421 4709 2455 4743
rect 2455 4709 2464 4743
rect 2412 4700 2464 4709
rect 2964 4700 3016 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 5448 4700 5500 4752
rect 8024 4768 8076 4820
rect 9036 4811 9088 4820
rect 9036 4777 9045 4811
rect 9045 4777 9079 4811
rect 9079 4777 9088 4811
rect 9036 4768 9088 4777
rect 9772 4768 9824 4820
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 12808 4768 12860 4820
rect 14556 4811 14608 4820
rect 14556 4777 14565 4811
rect 14565 4777 14599 4811
rect 14599 4777 14608 4811
rect 14556 4768 14608 4777
rect 14740 4768 14792 4820
rect 6184 4700 6236 4752
rect 8668 4700 8720 4752
rect 10508 4743 10560 4752
rect 10508 4709 10517 4743
rect 10517 4709 10551 4743
rect 10551 4709 10560 4743
rect 10508 4700 10560 4709
rect 12256 4700 12308 4752
rect 13360 4700 13412 4752
rect 15844 4700 15896 4752
rect 112 4564 164 4616
rect 2780 4607 2832 4616
rect 2780 4573 2789 4607
rect 2789 4573 2823 4607
rect 2823 4573 2832 4607
rect 2780 4564 2832 4573
rect 3148 4496 3200 4548
rect 5356 4675 5408 4684
rect 5356 4641 5365 4675
rect 5365 4641 5399 4675
rect 5399 4641 5408 4675
rect 5356 4632 5408 4641
rect 6828 4675 6880 4684
rect 6828 4641 6842 4675
rect 6842 4641 6880 4675
rect 6828 4632 6880 4641
rect 8024 4632 8076 4684
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 11888 4632 11940 4684
rect 12532 4632 12584 4684
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 15384 4632 15436 4684
rect 17224 4632 17276 4684
rect 18420 4632 18472 4684
rect 8760 4607 8812 4616
rect 8760 4573 8769 4607
rect 8769 4573 8803 4607
rect 8803 4573 8812 4607
rect 8760 4564 8812 4573
rect 9588 4564 9640 4616
rect 10876 4564 10928 4616
rect 11244 4564 11296 4616
rect 12992 4564 13044 4616
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 14372 4564 14424 4616
rect 10048 4496 10100 4548
rect 13636 4496 13688 4548
rect 15292 4496 15344 4548
rect 2320 4428 2372 4480
rect 3056 4428 3108 4480
rect 4344 4428 4396 4480
rect 4620 4471 4672 4480
rect 4620 4437 4629 4471
rect 4629 4437 4663 4471
rect 4663 4437 4672 4471
rect 4620 4428 4672 4437
rect 6368 4428 6420 4480
rect 6460 4428 6512 4480
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 7012 4428 7064 4480
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 16396 4471 16448 4480
rect 16396 4437 16405 4471
rect 16405 4437 16439 4471
rect 16439 4437 16448 4471
rect 16396 4428 16448 4437
rect 18880 4471 18932 4480
rect 18880 4437 18889 4471
rect 18889 4437 18923 4471
rect 18923 4437 18932 4471
rect 18880 4428 18932 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1584 4224 1636 4276
rect 3240 4224 3292 4276
rect 3792 4224 3844 4276
rect 4068 4267 4120 4276
rect 4068 4233 4077 4267
rect 4077 4233 4111 4267
rect 4111 4233 4120 4267
rect 4068 4224 4120 4233
rect 6368 4267 6420 4276
rect 2320 4156 2372 4208
rect 4252 4156 4304 4208
rect 4620 4156 4672 4208
rect 4896 4199 4948 4208
rect 4896 4165 4905 4199
rect 4905 4165 4939 4199
rect 4939 4165 4948 4199
rect 6368 4233 6377 4267
rect 6377 4233 6411 4267
rect 6411 4233 6420 4267
rect 6368 4224 6420 4233
rect 6460 4224 6512 4276
rect 10508 4224 10560 4276
rect 17040 4224 17092 4276
rect 18420 4224 18472 4276
rect 4896 4156 4948 4165
rect 5448 4156 5500 4208
rect 1492 4063 1544 4072
rect 1492 4029 1501 4063
rect 1501 4029 1535 4063
rect 1535 4029 1544 4063
rect 1492 4020 1544 4029
rect 2964 4063 3016 4072
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 3148 4020 3200 4072
rect 3516 4020 3568 4072
rect 4068 4020 4120 4072
rect 2320 3884 2372 3936
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 4344 4020 4396 4072
rect 6920 4088 6972 4140
rect 10692 4156 10744 4208
rect 10876 4156 10928 4208
rect 11888 4199 11940 4208
rect 11888 4165 11897 4199
rect 11897 4165 11931 4199
rect 11931 4165 11940 4199
rect 11888 4156 11940 4165
rect 12256 4199 12308 4208
rect 12256 4165 12265 4199
rect 12265 4165 12299 4199
rect 12299 4165 12308 4199
rect 12256 4156 12308 4165
rect 14648 4156 14700 4208
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 11796 4088 11848 4140
rect 12808 4131 12860 4140
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 12992 4088 13044 4140
rect 16396 4088 16448 4140
rect 4620 3995 4672 4004
rect 4620 3961 4629 3995
rect 4629 3961 4663 3995
rect 4663 3961 4672 3995
rect 4620 3952 4672 3961
rect 6828 3952 6880 4004
rect 2780 3884 2832 3893
rect 4344 3884 4396 3936
rect 5080 3884 5132 3936
rect 5356 3884 5408 3936
rect 6460 3884 6512 3936
rect 8484 4020 8536 4072
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 11244 4020 11296 4029
rect 12624 4063 12676 4072
rect 12624 4029 12633 4063
rect 12633 4029 12667 4063
rect 12667 4029 12676 4063
rect 12624 4020 12676 4029
rect 8852 3995 8904 4004
rect 8852 3961 8861 3995
rect 8861 3961 8895 3995
rect 8895 3961 8904 3995
rect 8852 3952 8904 3961
rect 9864 3995 9916 4004
rect 9864 3961 9873 3995
rect 9873 3961 9907 3995
rect 9907 3961 9916 3995
rect 9864 3952 9916 3961
rect 11520 3952 11572 4004
rect 13360 3952 13412 4004
rect 8944 3884 8996 3936
rect 10048 3884 10100 3936
rect 12348 3884 12400 3936
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 14648 3995 14700 4004
rect 14648 3961 14657 3995
rect 14657 3961 14691 3995
rect 14691 3961 14700 3995
rect 14648 3952 14700 3961
rect 15752 3952 15804 4004
rect 16304 3995 16356 4004
rect 16304 3961 16313 3995
rect 16313 3961 16347 3995
rect 16347 3961 16356 3995
rect 16304 3952 16356 3961
rect 16396 3952 16448 4004
rect 17592 3952 17644 4004
rect 15844 3884 15896 3936
rect 17224 3927 17276 3936
rect 17224 3893 17233 3927
rect 17233 3893 17267 3927
rect 17267 3893 17276 3927
rect 17224 3884 17276 3893
rect 17408 3884 17460 3936
rect 17500 3884 17552 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1400 3680 1452 3732
rect 3516 3723 3568 3732
rect 3516 3689 3525 3723
rect 3525 3689 3559 3723
rect 3559 3689 3568 3723
rect 3516 3680 3568 3689
rect 3700 3680 3752 3732
rect 4620 3680 4672 3732
rect 6184 3680 6236 3732
rect 6460 3723 6512 3732
rect 6460 3689 6469 3723
rect 6469 3689 6503 3723
rect 6503 3689 6512 3723
rect 6460 3680 6512 3689
rect 8024 3723 8076 3732
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 8760 3680 8812 3732
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 9864 3680 9916 3732
rect 12808 3723 12860 3732
rect 12808 3689 12817 3723
rect 12817 3689 12851 3723
rect 12851 3689 12860 3723
rect 12808 3680 12860 3689
rect 13360 3723 13412 3732
rect 13360 3689 13369 3723
rect 13369 3689 13403 3723
rect 13403 3689 13412 3723
rect 13360 3680 13412 3689
rect 4988 3612 5040 3664
rect 5172 3612 5224 3664
rect 7196 3655 7248 3664
rect 7196 3621 7205 3655
rect 7205 3621 7239 3655
rect 7239 3621 7248 3655
rect 7196 3612 7248 3621
rect 7840 3612 7892 3664
rect 10048 3655 10100 3664
rect 10048 3621 10051 3655
rect 10051 3621 10085 3655
rect 10085 3621 10100 3655
rect 10048 3612 10100 3621
rect 11520 3655 11572 3664
rect 11520 3621 11529 3655
rect 11529 3621 11563 3655
rect 11563 3621 11572 3655
rect 11520 3612 11572 3621
rect 11612 3655 11664 3664
rect 11612 3621 11621 3655
rect 11621 3621 11655 3655
rect 11655 3621 11664 3655
rect 11612 3612 11664 3621
rect 12992 3612 13044 3664
rect 15752 3680 15804 3732
rect 15660 3612 15712 3664
rect 1308 3544 1360 3596
rect 1584 3544 1636 3596
rect 2228 3587 2280 3596
rect 2228 3553 2237 3587
rect 2237 3553 2271 3587
rect 2271 3553 2280 3587
rect 2228 3544 2280 3553
rect 3056 3587 3108 3596
rect 3056 3553 3065 3587
rect 3065 3553 3099 3587
rect 3099 3553 3108 3587
rect 3056 3544 3108 3553
rect 4528 3544 4580 3596
rect 4712 3544 4764 3596
rect 6552 3544 6604 3596
rect 8576 3587 8628 3596
rect 8576 3553 8585 3587
rect 8585 3553 8619 3587
rect 8619 3553 8628 3587
rect 8576 3544 8628 3553
rect 16304 3612 16356 3664
rect 17316 3544 17368 3596
rect 19064 3587 19116 3596
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 4896 3476 4948 3528
rect 5264 3519 5316 3528
rect 5264 3485 5273 3519
rect 5273 3485 5307 3519
rect 5307 3485 5316 3519
rect 5264 3476 5316 3485
rect 6644 3476 6696 3528
rect 7104 3519 7156 3528
rect 7104 3485 7113 3519
rect 7113 3485 7147 3519
rect 7147 3485 7156 3519
rect 7104 3476 7156 3485
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 8852 3476 8904 3528
rect 4344 3408 4396 3460
rect 11244 3408 11296 3460
rect 12992 3519 13044 3528
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 14280 3476 14332 3528
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 15476 3476 15528 3528
rect 14832 3408 14884 3460
rect 4436 3340 4488 3392
rect 7196 3340 7248 3392
rect 8484 3340 8536 3392
rect 15752 3340 15804 3392
rect 16488 3408 16540 3460
rect 20260 3408 20312 3460
rect 17960 3340 18012 3392
rect 18052 3340 18104 3392
rect 19524 3340 19576 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1308 3136 1360 3188
rect 2964 3179 3016 3188
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 5172 3136 5224 3188
rect 6276 3136 6328 3188
rect 6552 3179 6604 3188
rect 6552 3145 6561 3179
rect 6561 3145 6595 3179
rect 6595 3145 6604 3179
rect 6552 3136 6604 3145
rect 7012 3136 7064 3188
rect 7840 3179 7892 3188
rect 7840 3145 7849 3179
rect 7849 3145 7883 3179
rect 7883 3145 7892 3179
rect 7840 3136 7892 3145
rect 8852 3179 8904 3188
rect 8852 3145 8861 3179
rect 8861 3145 8895 3179
rect 8895 3145 8904 3179
rect 8852 3136 8904 3145
rect 8944 3136 8996 3188
rect 11060 3179 11112 3188
rect 4344 3068 4396 3120
rect 4528 3111 4580 3120
rect 4528 3077 4537 3111
rect 4537 3077 4571 3111
rect 4571 3077 4580 3111
rect 4528 3068 4580 3077
rect 6000 3068 6052 3120
rect 7104 3068 7156 3120
rect 2136 3000 2188 3052
rect 5264 3000 5316 3052
rect 6368 3000 6420 3052
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 848 2932 900 2984
rect 1492 2975 1544 2984
rect 1492 2941 1501 2975
rect 1501 2941 1535 2975
rect 1535 2941 1544 2975
rect 1492 2932 1544 2941
rect 2412 2932 2464 2984
rect 3884 2975 3936 2984
rect 1860 2864 1912 2916
rect 3884 2941 3893 2975
rect 3893 2941 3927 2975
rect 3927 2941 3936 2975
rect 4988 2975 5040 2984
rect 3884 2932 3936 2941
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 5080 2864 5132 2916
rect 5172 2864 5224 2916
rect 4988 2796 5040 2848
rect 6736 2864 6788 2916
rect 7012 2907 7064 2916
rect 7012 2873 7021 2907
rect 7021 2873 7055 2907
rect 7055 2873 7064 2907
rect 7564 2907 7616 2916
rect 7012 2864 7064 2873
rect 7564 2873 7573 2907
rect 7573 2873 7607 2907
rect 7607 2873 7616 2907
rect 7564 2864 7616 2873
rect 11060 3145 11069 3179
rect 11069 3145 11103 3179
rect 11103 3145 11112 3179
rect 11060 3136 11112 3145
rect 12992 3136 13044 3188
rect 13360 3136 13412 3188
rect 13544 3136 13596 3188
rect 15384 3136 15436 3188
rect 15660 3179 15712 3188
rect 15660 3145 15669 3179
rect 15669 3145 15703 3179
rect 15703 3145 15712 3179
rect 15660 3136 15712 3145
rect 16580 3136 16632 3188
rect 17316 3179 17368 3188
rect 17316 3145 17325 3179
rect 17325 3145 17359 3179
rect 17359 3145 17368 3179
rect 17316 3136 17368 3145
rect 17408 3136 17460 3188
rect 11612 3068 11664 3120
rect 12716 3068 12768 3120
rect 17960 3068 18012 3120
rect 19064 3111 19116 3120
rect 11060 2932 11112 2984
rect 14740 3000 14792 3052
rect 16488 3000 16540 3052
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 17040 3000 17092 3052
rect 19064 3077 19073 3111
rect 19073 3077 19107 3111
rect 19107 3077 19116 3111
rect 19064 3068 19116 3077
rect 9956 2864 10008 2916
rect 13452 2864 13504 2916
rect 7196 2796 7248 2848
rect 10692 2796 10744 2848
rect 11612 2796 11664 2848
rect 15936 2796 15988 2848
rect 16488 2907 16540 2916
rect 16488 2873 16497 2907
rect 16497 2873 16531 2907
rect 16531 2873 16540 2907
rect 16488 2864 16540 2873
rect 23848 2864 23900 2916
rect 20168 2796 20220 2848
rect 20904 2796 20956 2848
rect 25964 2796 26016 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 3424 2592 3476 2644
rect 3884 2592 3936 2644
rect 4528 2635 4580 2644
rect 4528 2601 4537 2635
rect 4537 2601 4571 2635
rect 4571 2601 4580 2635
rect 4528 2592 4580 2601
rect 5356 2592 5408 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 6644 2635 6696 2644
rect 6644 2601 6653 2635
rect 6653 2601 6687 2635
rect 6687 2601 6696 2635
rect 6644 2592 6696 2601
rect 4988 2524 5040 2576
rect 7564 2592 7616 2644
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 9956 2635 10008 2644
rect 9956 2601 9965 2635
rect 9965 2601 9999 2635
rect 9999 2601 10008 2635
rect 9956 2592 10008 2601
rect 12348 2635 12400 2644
rect 12348 2601 12357 2635
rect 12357 2601 12391 2635
rect 12391 2601 12400 2635
rect 12348 2592 12400 2601
rect 13360 2635 13412 2644
rect 13360 2601 13369 2635
rect 13369 2601 13403 2635
rect 13403 2601 13412 2635
rect 13360 2592 13412 2601
rect 15936 2635 15988 2644
rect 15936 2601 15945 2635
rect 15945 2601 15979 2635
rect 15979 2601 15988 2635
rect 15936 2592 15988 2601
rect 16212 2592 16264 2644
rect 4804 2456 4856 2508
rect 7104 2567 7156 2576
rect 7104 2533 7113 2567
rect 7113 2533 7147 2567
rect 7147 2533 7156 2567
rect 7104 2524 7156 2533
rect 11520 2524 11572 2576
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 15476 2524 15528 2576
rect 16580 2524 16632 2576
rect 14832 2456 14884 2508
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 5356 2388 5408 2397
rect 7288 2320 7340 2372
rect 2412 2252 2464 2304
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 9220 2320 9272 2372
rect 11612 2320 11664 2372
rect 8576 2252 8628 2304
rect 15568 2456 15620 2508
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 20168 2592 20220 2644
rect 20260 2592 20312 2644
rect 19524 2456 19576 2508
rect 24860 2524 24912 2576
rect 18696 2388 18748 2440
rect 17500 2252 17552 2304
rect 19708 2252 19760 2304
rect 21456 2252 21508 2304
rect 23204 2252 23256 2304
rect 27068 2252 27120 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 4344 76 4396 128
rect 8392 76 8444 128
rect 18880 76 18932 128
rect 20628 76 20680 128
<< metal2 >>
rect 938 27520 994 28000
rect 2870 27520 2926 28000
rect 4894 27554 4950 28000
rect 4816 27526 4950 27554
rect 952 23662 980 27520
rect 2884 24274 2912 27520
rect 3146 24984 3202 24993
rect 3146 24919 3202 24928
rect 2872 24268 2924 24274
rect 2872 24210 2924 24216
rect 2884 23866 2912 24210
rect 3160 23866 3188 24919
rect 3608 24064 3660 24070
rect 3608 24006 3660 24012
rect 2872 23860 2924 23866
rect 2872 23802 2924 23808
rect 3148 23860 3200 23866
rect 3148 23802 3200 23808
rect 3424 23792 3476 23798
rect 3424 23734 3476 23740
rect 940 23656 992 23662
rect 940 23598 992 23604
rect 1308 23520 1360 23526
rect 1308 23462 1360 23468
rect 1582 23488 1638 23497
rect 1214 20088 1270 20097
rect 1214 20023 1270 20032
rect 1228 19310 1256 20023
rect 1216 19304 1268 19310
rect 1216 19246 1268 19252
rect 1320 15502 1348 23462
rect 1582 23423 1638 23432
rect 1596 22778 1624 23423
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 2044 22432 2096 22438
rect 2044 22374 2096 22380
rect 1582 21720 1638 21729
rect 1582 21655 1638 21664
rect 1596 20602 1624 21655
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 1400 19168 1452 19174
rect 1400 19110 1452 19116
rect 1412 15609 1440 19110
rect 1780 18970 1808 20334
rect 2056 18970 2084 22374
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 2964 18828 3016 18834
rect 2964 18770 3016 18776
rect 1688 17542 1716 18770
rect 2412 18624 2464 18630
rect 2412 18566 2464 18572
rect 2424 18222 2452 18566
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1492 17060 1544 17066
rect 1492 17002 1544 17008
rect 1398 15600 1454 15609
rect 1398 15535 1454 15544
rect 1308 15496 1360 15502
rect 1308 15438 1360 15444
rect 1504 9586 1532 17002
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1688 15706 1716 16594
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1780 16250 1808 16526
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 1780 15910 1808 16186
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1582 15192 1638 15201
rect 1582 15127 1638 15136
rect 1596 14482 1624 15127
rect 1688 14890 1716 15642
rect 1860 15632 1912 15638
rect 1860 15574 1912 15580
rect 1676 14884 1728 14890
rect 1676 14826 1728 14832
rect 1872 14822 1900 15574
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1596 14074 1624 14418
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1688 11558 1716 12242
rect 1780 11830 1808 14214
rect 1872 12850 1900 14758
rect 1964 13326 1992 18022
rect 2424 17746 2452 18158
rect 2976 18086 3004 18770
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2148 17134 2176 17682
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 2240 14618 2268 14826
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 2056 13734 2084 14214
rect 2240 14074 2268 14554
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2332 13938 2360 17614
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 15978 2728 17478
rect 2976 17241 3004 18022
rect 2962 17232 3018 17241
rect 2962 17167 3018 17176
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2884 16454 2912 17070
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3146 16824 3202 16833
rect 3146 16759 3202 16768
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2700 15094 2728 15914
rect 2688 15088 2740 15094
rect 2688 15030 2740 15036
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 2056 13462 2084 13670
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1952 12640 2004 12646
rect 2056 12628 2084 13398
rect 2516 13258 2544 14350
rect 2792 13734 2820 14486
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2504 13252 2556 13258
rect 2504 13194 2556 13200
rect 2004 12600 2084 12628
rect 1952 12582 2004 12588
rect 1768 11824 1820 11830
rect 1768 11766 1820 11772
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11014 1716 11494
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1688 10810 1716 10950
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1584 9444 1636 9450
rect 1584 9386 1636 9392
rect 1596 8838 1624 9386
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1214 8528 1270 8537
rect 1214 8463 1270 8472
rect 110 7440 166 7449
rect 110 7375 166 7384
rect 124 7342 152 7375
rect 112 7336 164 7342
rect 112 7278 164 7284
rect 1228 5778 1256 8463
rect 1216 5772 1268 5778
rect 1216 5714 1268 5720
rect 1228 4826 1256 5714
rect 1398 5264 1454 5273
rect 1398 5199 1454 5208
rect 1216 4820 1268 4826
rect 1216 4762 1268 4768
rect 1412 4690 1440 5199
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 112 4616 164 4622
rect 112 4558 164 4564
rect 124 4185 152 4558
rect 110 4176 166 4185
rect 110 4111 166 4120
rect 1412 3738 1440 4626
rect 1596 4282 1624 8774
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 6118 1716 7686
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1780 5234 1808 10542
rect 1964 10470 1992 12582
rect 2608 12442 2636 13262
rect 2792 13190 2820 13670
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2792 12782 2820 13126
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2056 11286 2084 12038
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2044 11280 2096 11286
rect 2044 11222 2096 11228
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 9908 1992 10406
rect 2056 10266 2084 11222
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2148 10130 2176 10406
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2044 9920 2096 9926
rect 1964 9880 2044 9908
rect 2044 9862 2096 9868
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1872 7750 1900 8910
rect 1964 8498 1992 9046
rect 2056 8838 2084 9862
rect 2148 8906 2176 10066
rect 2332 9450 2360 11494
rect 2516 11286 2544 11562
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2516 10674 2544 11222
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2884 10266 2912 16390
rect 3160 16250 3188 16759
rect 3148 16244 3200 16250
rect 3148 16186 3200 16192
rect 3160 16046 3188 16186
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2976 15026 3004 15302
rect 3068 15094 3096 15846
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3160 15162 3188 15438
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3056 15088 3108 15094
rect 3056 15030 3108 15036
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 2976 14414 3004 14962
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 3068 11257 3096 12718
rect 3252 12238 3280 16934
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3252 11898 3280 12174
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3160 11354 3188 11494
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3054 11248 3110 11257
rect 3054 11183 3110 11192
rect 2872 10260 2924 10266
rect 2924 10220 3004 10248
rect 2872 10202 2924 10208
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2608 9722 2636 9862
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2700 9674 2728 9998
rect 2700 9646 2820 9674
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1964 7954 1992 8298
rect 2056 8090 2084 8774
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 5914 1900 7686
rect 2056 7206 2084 8026
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2056 6662 2084 7142
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1964 5166 1992 5850
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1964 4758 1992 5102
rect 1952 4752 2004 4758
rect 1872 4712 1952 4740
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 1308 3596 1360 3602
rect 1308 3538 1360 3544
rect 1504 3584 1532 4014
rect 1584 3596 1636 3602
rect 1504 3556 1584 3584
rect 1320 3194 1348 3538
rect 1308 3188 1360 3194
rect 1308 3130 1360 3136
rect 1504 2990 1532 3556
rect 1584 3538 1636 3544
rect 848 2984 900 2990
rect 848 2926 900 2932
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 570 82 626 480
rect 860 82 888 2926
rect 1872 2922 1900 4712
rect 1952 4694 2004 4700
rect 2056 4154 2084 6598
rect 1964 4126 2084 4154
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 570 54 888 82
rect 1674 82 1730 480
rect 1964 82 1992 4126
rect 2148 3058 2176 8842
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2240 6322 2268 8570
rect 2318 7848 2374 7857
rect 2318 7783 2374 7792
rect 2332 7002 2360 7783
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2240 5914 2268 6258
rect 2332 6254 2360 6938
rect 2424 6882 2452 9318
rect 2792 8974 2820 9646
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2516 8566 2544 8910
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 2516 7002 2544 8502
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2700 8294 2728 8366
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2700 8090 2728 8230
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2596 6928 2648 6934
rect 2424 6854 2544 6882
rect 2596 6870 2648 6876
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2240 3602 2268 5510
rect 2424 4758 2452 5646
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4214 2360 4422
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 2516 4154 2544 6854
rect 2608 6118 2636 6870
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2792 4622 2820 8910
rect 2976 7290 3004 10220
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 8838 3280 9318
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3068 7410 3096 8026
rect 3436 7546 3464 23734
rect 3620 15162 3648 24006
rect 4816 23866 4844 27526
rect 4894 27520 4950 27526
rect 6918 27554 6974 28000
rect 6918 27526 7052 27554
rect 6918 27520 6974 27526
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 7024 23866 7052 27526
rect 7748 27532 7800 27538
rect 8850 27532 8906 28000
rect 8850 27520 8852 27532
rect 7748 27474 7800 27480
rect 8904 27520 8906 27532
rect 10874 27520 10930 28000
rect 12898 27554 12954 28000
rect 12544 27526 12954 27554
rect 8852 27474 8904 27480
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 4816 23662 4844 23802
rect 4804 23656 4856 23662
rect 4804 23598 4856 23604
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 3974 18456 4030 18465
rect 3974 18391 4030 18400
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 3712 16998 3740 17682
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3712 16794 3740 16934
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3620 15026 3648 15098
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 10146 3556 13126
rect 3804 12918 3832 18090
rect 3988 17134 4016 18391
rect 4080 17882 4108 23462
rect 7484 23322 7512 23598
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 7760 17882 7788 27474
rect 8864 27443 8892 27474
rect 8298 26616 8354 26625
rect 8298 26551 8354 26560
rect 8312 23730 8340 26551
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10888 23866 10916 27520
rect 12544 24274 12572 27526
rect 12898 27520 12954 27526
rect 14922 27520 14978 28000
rect 16854 27520 16910 28000
rect 18878 27520 18934 28000
rect 20902 27520 20958 28000
rect 22834 27520 22890 28000
rect 24858 27520 24914 28000
rect 26882 27520 26938 28000
rect 14936 25650 14964 27520
rect 14844 25622 14964 25650
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 11992 23866 12020 24210
rect 12716 24132 12768 24138
rect 12716 24074 12768 24080
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 11980 23860 12032 23866
rect 11980 23802 12032 23808
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 8484 22976 8536 22982
rect 8484 22918 8536 22924
rect 8496 22438 8524 22918
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 8484 22432 8536 22438
rect 8484 22374 8536 22380
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 4632 17338 4660 17682
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 4620 17332 4672 17338
rect 4540 17292 4620 17320
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3896 15366 3924 16390
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3804 11762 3832 12854
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3620 10266 3648 10610
rect 3712 10538 3740 10950
rect 3700 10532 3752 10538
rect 3700 10474 3752 10480
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3528 10118 3648 10146
rect 3620 9602 3648 10118
rect 3712 9722 3740 10474
rect 3896 10198 3924 15302
rect 3988 13814 4016 16594
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 4356 15910 4384 16390
rect 4436 15972 4488 15978
rect 4436 15914 4488 15920
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4448 15162 4476 15914
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4448 14890 4476 15098
rect 4436 14884 4488 14890
rect 4436 14826 4488 14832
rect 4540 14414 4568 17292
rect 4620 17274 4672 17280
rect 7392 17270 7420 17682
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 6184 17060 6236 17066
rect 6184 17002 6236 17008
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 5000 16250 5028 16594
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5092 16046 5120 16390
rect 5080 16040 5132 16046
rect 5132 16000 5212 16028
rect 5080 15982 5132 15988
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4632 14550 4660 15302
rect 5000 15162 5028 15506
rect 4988 15156 5040 15162
rect 4908 15116 4988 15144
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4080 14074 4108 14350
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4540 14006 4568 14350
rect 4632 14074 4660 14486
rect 4724 14278 4752 14962
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4724 13938 4752 14214
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 3988 13786 4108 13814
rect 4908 13802 4936 15116
rect 4988 15098 5040 15104
rect 4080 12306 4108 13786
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4908 13530 4936 13738
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 3988 11218 4016 11727
rect 4080 11694 4108 12242
rect 4172 12102 4200 12718
rect 4356 12442 4384 13262
rect 4632 12714 4660 13466
rect 5080 13456 5132 13462
rect 5184 13444 5212 16000
rect 5460 15910 5488 16526
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5132 13416 5212 13444
rect 5080 13398 5132 13404
rect 5184 12986 5212 13416
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 5184 12442 5212 12922
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4080 11354 4108 11630
rect 4172 11558 4200 12038
rect 5092 11694 5120 12242
rect 5276 12102 5304 15846
rect 5460 12238 5488 15846
rect 6196 15502 6224 17002
rect 7392 16794 7420 17206
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7576 16726 7604 16934
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6288 16114 6316 16594
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6656 16250 6684 16526
rect 7576 16250 7604 16662
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 7668 15978 7696 17070
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7484 15638 7512 15914
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6196 15162 6224 15438
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6840 15094 6868 15574
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 7484 15026 7512 15574
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7668 14618 7696 15914
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7760 14890 7788 15302
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6380 13326 6408 14214
rect 7024 13734 7052 14554
rect 7760 14074 7788 14826
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3988 10810 4016 11154
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3516 9580 3568 9586
rect 3620 9574 3740 9602
rect 3516 9522 3568 9528
rect 3528 9178 3556 9522
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 2872 7268 2924 7274
rect 2976 7262 3096 7290
rect 2872 7210 2924 7216
rect 2884 6934 2912 7210
rect 2872 6928 2924 6934
rect 2872 6870 2924 6876
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2976 6458 3004 6734
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 3068 6168 3096 7262
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3252 6322 3280 6938
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3528 6322 3556 6734
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3528 6225 3556 6258
rect 2976 6140 3096 6168
rect 3514 6216 3570 6225
rect 3620 6186 3648 7142
rect 3514 6151 3570 6160
rect 3608 6180 3660 6186
rect 2976 5370 3004 6140
rect 3608 6122 3660 6128
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2976 5166 3004 5306
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 3068 5098 3096 5714
rect 3160 5234 3188 6054
rect 3620 5914 3648 6122
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3620 5166 3648 5850
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3056 5092 3108 5098
rect 3056 5034 3108 5040
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2332 3942 2360 4150
rect 2424 4126 2544 4154
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2332 1465 2360 3878
rect 2424 2990 2452 4126
rect 2792 3942 2820 4558
rect 2976 4078 3004 4694
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2792 3097 2820 3878
rect 2976 3194 3004 4014
rect 3068 3602 3096 4422
rect 3160 4078 3188 4490
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3252 3913 3280 4218
rect 3422 4176 3478 4185
rect 3422 4111 3478 4120
rect 3238 3904 3294 3913
rect 3238 3839 3294 3848
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2778 3088 2834 3097
rect 2778 3023 2834 3032
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2424 2310 2452 2926
rect 3436 2650 3464 4111
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3528 3738 3556 4014
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 2318 1456 2374 1465
rect 2318 1391 2374 1400
rect 1674 54 1992 82
rect 2424 82 2452 2246
rect 2778 82 2834 480
rect 2424 54 2834 82
rect 3620 82 3648 4966
rect 3712 3738 3740 9574
rect 3896 8294 3924 10134
rect 4264 9722 4292 10134
rect 4816 10062 4844 10610
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4448 9722 4476 9998
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4448 9178 4476 9658
rect 4816 9625 4844 9998
rect 4802 9616 4858 9625
rect 4802 9551 4858 9560
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 4842 3924 8230
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3804 4814 3924 4842
rect 3804 4282 3832 4814
rect 4080 4282 4108 6054
rect 4448 4826 4476 8774
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4250 4312 4306 4321
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 4068 4276 4120 4282
rect 4250 4247 4306 4256
rect 4068 4218 4120 4224
rect 4080 4078 4108 4218
rect 4264 4214 4292 4247
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4356 4078 4384 4422
rect 4540 4154 4568 9114
rect 4908 9110 4936 11630
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5092 10198 5120 10474
rect 5276 10470 5304 11154
rect 5368 11014 5396 11494
rect 5920 11286 5948 11494
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4908 8634 4936 9046
rect 5276 9042 5304 10406
rect 5368 9926 5396 10950
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5276 8634 5304 8978
rect 5368 8974 5396 9862
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5460 8566 5488 10406
rect 5736 10266 5764 10542
rect 6012 10266 6040 12786
rect 6196 12345 6224 13262
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6182 12336 6238 12345
rect 6092 12300 6144 12306
rect 6182 12271 6238 12280
rect 6092 12242 6144 12248
rect 6104 11558 6132 12242
rect 6184 12164 6236 12170
rect 6288 12152 6316 12922
rect 6656 12646 6684 13670
rect 6734 13424 6790 13433
rect 6734 13359 6790 13368
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6236 12124 6316 12152
rect 6184 12106 6236 12112
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6196 11218 6224 12106
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6276 11552 6328 11558
rect 6472 11540 6500 12038
rect 6564 11898 6592 12174
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6328 11512 6500 11540
rect 6276 11494 6328 11500
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6196 10470 6224 11154
rect 6288 10742 6316 11494
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6288 9994 6316 10678
rect 6472 10674 6500 10950
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6656 10470 6684 12582
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6472 9586 6500 10134
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6472 9178 6500 9386
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6656 9110 6684 10406
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5460 8430 5488 8502
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4632 7954 4660 8298
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 8090 5120 8230
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4724 6458 4752 7822
rect 5368 7274 5396 7890
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5368 7002 5396 7210
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4894 6896 4950 6905
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4724 6168 4752 6394
rect 4816 6322 4844 6870
rect 4894 6831 4950 6840
rect 4908 6798 4936 6831
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6390 4936 6734
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4804 6180 4856 6186
rect 4724 6140 4804 6168
rect 4804 6122 4856 6128
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4724 5030 4752 5714
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 4214 4660 4422
rect 4448 4126 4568 4154
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 4356 3466 4384 3878
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4448 3398 4476 4126
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4632 3738 4660 3946
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4724 3602 4752 4966
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4894 4312 4950 4321
rect 4894 4247 4950 4256
rect 4908 4214 4936 4247
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 5000 3670 5028 4762
rect 5368 4690 5396 4966
rect 5460 4758 5488 8366
rect 5828 7954 5856 8366
rect 6196 8294 6224 9046
rect 6748 8430 6776 13359
rect 7116 13190 7144 13874
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7116 12646 7144 13126
rect 7392 12782 7420 13262
rect 7760 12986 7788 13330
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7392 12374 7420 12718
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7208 11354 7236 11698
rect 7300 11558 7328 12106
rect 7852 11830 7880 22374
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 7932 16516 7984 16522
rect 7932 16458 7984 16464
rect 7944 16114 7972 16458
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 8220 15706 8248 16526
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8036 14074 8064 14350
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8036 13530 8064 14010
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 7024 10198 7052 11086
rect 7300 10538 7328 11494
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7484 10606 7512 11222
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7668 10266 7696 10610
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7852 10198 7880 11562
rect 8036 11286 8064 11766
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 7840 10192 7892 10198
rect 7840 10134 7892 10140
rect 7024 9586 7052 10134
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 8036 9382 8064 10406
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 6840 9178 6868 9318
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5828 7857 5856 7890
rect 5814 7848 5870 7857
rect 5814 7783 5870 7792
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5552 6322 5580 7346
rect 6196 6934 6224 8230
rect 7484 8090 7512 8910
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 6550 7984 6606 7993
rect 6550 7919 6552 7928
rect 6604 7919 6606 7928
rect 6552 7890 6604 7896
rect 6564 7206 6592 7890
rect 8036 7750 8064 9318
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7116 7206 7144 7686
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6196 6390 6224 6870
rect 6288 6458 6316 6870
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6184 6384 6236 6390
rect 6184 6326 6236 6332
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5552 5166 5580 5850
rect 5920 5846 5948 6122
rect 6196 6118 6224 6326
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5846 6224 6054
rect 6288 5914 6316 6394
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 5908 5840 5960 5846
rect 5722 5808 5778 5817
rect 5908 5782 5960 5788
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 5722 5743 5778 5752
rect 5736 5710 5764 5743
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 6012 4826 6040 5646
rect 6196 5012 6224 5782
rect 6380 5370 6408 6054
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6276 5024 6328 5030
rect 6196 4984 6276 5012
rect 6276 4966 6328 4972
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5368 3942 5396 4626
rect 5460 4214 5488 4694
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 6196 4146 6224 4694
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4540 3126 4568 3538
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3896 2650 3924 2926
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3882 82 3938 480
rect 4356 134 4384 3062
rect 4526 2952 4582 2961
rect 4526 2887 4582 2896
rect 4540 2650 4568 2887
rect 4908 2825 4936 3470
rect 5000 2990 5028 3606
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5092 2922 5120 3878
rect 6196 3738 6224 4082
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5184 3194 5212 3606
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5184 2922 5212 3130
rect 5276 3058 5304 3470
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6288 3194 6316 4966
rect 6380 4486 6408 5306
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6472 4282 6500 4422
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6380 4162 6408 4218
rect 6564 4162 6592 7142
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6748 6322 6776 6734
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6748 5914 6776 6258
rect 7116 6118 7144 7142
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 5234 6960 5510
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4690 6868 4966
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6748 4162 6776 4422
rect 6380 4134 6776 4162
rect 6840 4010 6868 4626
rect 6932 4146 6960 5170
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6460 3936 6512 3942
rect 6458 3904 6460 3913
rect 6512 3904 6514 3913
rect 6458 3839 6514 3848
rect 6472 3738 6500 3839
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 7024 3641 7052 4422
rect 7102 3768 7158 3777
rect 7102 3703 7158 3712
rect 7010 3632 7066 3641
rect 6552 3596 6604 3602
rect 7010 3567 7066 3576
rect 6552 3538 6604 3544
rect 6564 3194 6592 3538
rect 7116 3534 7144 3703
rect 7208 3670 7236 5714
rect 7300 5234 7328 6666
rect 7760 6662 7788 7278
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 5914 7788 6598
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 4988 2848 5040 2854
rect 4894 2816 4950 2825
rect 4988 2790 5040 2796
rect 4894 2751 4950 2760
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 5000 2582 5028 2790
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4816 2310 4844 2450
rect 5368 2446 5396 2586
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 3620 54 3938 82
rect 4344 128 4396 134
rect 4344 70 4396 76
rect 4816 82 4844 2246
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 4986 82 5042 480
rect 4816 54 5042 82
rect 6012 82 6040 3062
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6380 2650 6408 2994
rect 6656 2650 6684 3470
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7024 2922 7052 3130
rect 7116 3126 7144 3470
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 6736 2916 6788 2922
rect 7012 2916 7064 2922
rect 6788 2876 6960 2904
rect 6736 2858 6788 2864
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6932 2564 6960 2876
rect 7012 2858 7064 2864
rect 7208 2854 7236 3334
rect 7576 2922 7604 3470
rect 7668 3097 7696 5170
rect 7852 4486 7880 5646
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8036 4690 8064 4762
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 4185 7880 4422
rect 7838 4176 7894 4185
rect 7838 4111 7894 4120
rect 8036 3738 8064 4626
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7852 3194 7880 3606
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7654 3088 7710 3097
rect 7654 3023 7710 3032
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7104 2576 7156 2582
rect 6932 2536 7104 2564
rect 7104 2518 7156 2524
rect 7208 1873 7236 2790
rect 7576 2650 7604 2858
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7194 1864 7250 1873
rect 7194 1799 7250 1808
rect 6090 82 6146 480
rect 6012 54 6146 82
rect 570 0 626 54
rect 1674 0 1730 54
rect 2778 0 2834 54
rect 3882 0 3938 54
rect 4986 0 5042 54
rect 6090 0 6146 54
rect 7194 82 7250 480
rect 7300 82 7328 2314
rect 8220 2009 8248 14758
rect 8864 13814 8892 23462
rect 10152 18426 10180 23598
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 9588 17808 9640 17814
rect 9588 17750 9640 17756
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9140 17338 9168 17546
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9600 16998 9628 17750
rect 10152 17678 10180 18158
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10152 17202 10180 17614
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11164 17202 11192 17546
rect 11242 17232 11298 17241
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 11152 17196 11204 17202
rect 11242 17167 11298 17176
rect 11152 17138 11204 17144
rect 9784 17066 9812 17138
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 9600 16794 9628 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 10704 16726 10732 16934
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9048 16182 9076 16526
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 9508 15910 9536 16662
rect 10704 16114 10732 16662
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 9784 15978 9812 16050
rect 10690 16008 10746 16017
rect 9772 15972 9824 15978
rect 10690 15943 10746 15952
rect 9772 15914 9824 15920
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9508 15638 9536 15846
rect 9496 15632 9548 15638
rect 9496 15574 9548 15580
rect 9784 15570 9812 15914
rect 10704 15910 10732 15943
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9784 14618 9812 15506
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10796 14890 10824 15438
rect 11164 15026 11192 15846
rect 11256 15094 11284 17167
rect 11336 17060 11388 17066
rect 11336 17002 11388 17008
rect 11348 16658 11376 17002
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11348 16250 11376 16594
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 13938 8984 14214
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8772 13786 8892 13814
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8312 11558 8340 12038
rect 8588 11898 8616 12174
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8588 11354 8616 11834
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8588 10674 8616 11290
rect 8576 10668 8628 10674
rect 8496 10628 8576 10656
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8312 10130 8340 10542
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8312 9178 8340 10066
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8404 9382 8432 9590
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8312 7818 8340 8502
rect 8404 7993 8432 9318
rect 8496 8634 8524 10628
rect 8576 10610 8628 10616
rect 8576 10532 8628 10538
rect 8680 10520 8708 12242
rect 8628 10492 8708 10520
rect 8576 10474 8628 10480
rect 8680 10266 8708 10492
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8588 8838 8616 9522
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8588 8294 8616 8774
rect 8680 8430 8708 10202
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8390 7984 8446 7993
rect 8390 7919 8446 7928
rect 8588 7886 8616 8230
rect 8680 8022 8708 8366
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8312 7002 8340 7754
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8312 5302 8340 6938
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8312 4690 8340 5034
rect 8496 4690 8524 7686
rect 8588 7206 8616 7822
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8588 6361 8616 7142
rect 8680 7002 8708 7958
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8680 6730 8708 6938
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8574 6352 8630 6361
rect 8574 6287 8630 6296
rect 8680 4758 8708 6666
rect 8772 5710 8800 13786
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8956 12782 8984 13262
rect 9508 13190 9536 14350
rect 9784 14074 9812 14554
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9784 13530 9812 13738
rect 9876 13734 9904 14554
rect 11256 14346 11284 15030
rect 11348 14618 11376 16186
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10796 13530 10824 13874
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9140 12850 9168 13126
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 12374 8984 12718
rect 9692 12714 9720 13330
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12850 11192 13126
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 9692 12306 9720 12650
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10980 12442 11008 12718
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 9692 11898 9720 12242
rect 10152 11898 10180 12242
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8864 10470 8892 10678
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 9654 8892 10406
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 9048 9450 9076 11018
rect 9416 9926 9444 11086
rect 9784 11014 9812 11494
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9784 10742 9812 10950
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9416 9518 9444 9862
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 9048 9178 9076 9386
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8864 6186 8892 7142
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8496 4078 8524 4626
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8496 3738 8524 4014
rect 8772 3738 8800 4558
rect 8864 4128 8892 6122
rect 9048 5778 9076 9114
rect 9784 8566 9812 10678
rect 10060 10674 10088 11086
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10152 10130 10180 11834
rect 10612 11762 10640 12174
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10980 11354 11008 12378
rect 11336 12300 11388 12306
rect 11256 12260 11336 12288
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10980 10606 11008 11290
rect 11164 11286 11192 11494
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 9876 9722 9904 10066
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 10152 9586 10180 10066
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 9586 10364 9998
rect 10704 9926 10732 10542
rect 11164 10470 11192 11222
rect 11256 11014 11284 12260
rect 11336 12242 11388 12248
rect 11440 11234 11468 21898
rect 11624 21894 11652 23122
rect 12268 22574 12296 23258
rect 12360 22642 12388 24006
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12256 22568 12308 22574
rect 12452 22522 12480 23462
rect 12636 23338 12664 24006
rect 12728 23594 12756 24074
rect 13464 23866 13492 24210
rect 14844 23866 14872 25622
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 16868 24410 16896 27520
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 15844 24268 15896 24274
rect 15844 24210 15896 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15856 23866 15884 24210
rect 18892 23866 18920 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 16488 23860 16540 23866
rect 16488 23802 16540 23808
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12716 23588 12768 23594
rect 12716 23530 12768 23536
rect 12256 22510 12308 22516
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 11888 20800 11940 20806
rect 11888 20742 11940 20748
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11624 15162 11652 15506
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11624 14550 11652 15098
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11532 13433 11560 14350
rect 11624 14074 11652 14486
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11518 13424 11574 13433
rect 11518 13359 11574 13368
rect 11716 12646 11744 13466
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11532 11626 11560 12582
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11808 11676 11836 12174
rect 11900 11898 11928 20742
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11888 11688 11940 11694
rect 11808 11648 11888 11676
rect 11888 11630 11940 11636
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11440 11206 11560 11234
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11256 10810 11284 10950
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11440 10674 11468 11086
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10704 9722 10732 9862
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 6866 9168 7278
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9140 6769 9168 6802
rect 9126 6760 9182 6769
rect 9126 6695 9182 6704
rect 9232 6458 9260 7210
rect 9876 7206 9904 7890
rect 10060 7410 10088 9318
rect 10152 9178 10180 9522
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 9178 10732 9522
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 8634 10180 8774
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10520 7546 10548 7822
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10888 7410 10916 8910
rect 10980 8430 11008 9590
rect 11164 9450 11192 10406
rect 11440 10266 11468 10610
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11532 10198 11560 11206
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11242 9208 11298 9217
rect 11532 9178 11560 10134
rect 11624 9450 11652 10134
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11612 9444 11664 9450
rect 11612 9386 11664 9392
rect 11242 9143 11298 9152
rect 11520 9172 11572 9178
rect 11256 9110 11284 9143
rect 11520 9114 11572 9120
rect 11244 9104 11296 9110
rect 11244 9046 11296 9052
rect 11256 8634 11284 9046
rect 11808 8906 11836 9998
rect 11900 9722 11928 11630
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11900 9042 11928 9658
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6934 9904 7142
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10888 7002 10916 7346
rect 10980 7274 11008 7482
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9218 6352 9274 6361
rect 9218 6287 9274 6296
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9140 5914 9168 6054
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9036 5772 9088 5778
rect 8956 5732 9036 5760
rect 8956 5166 8984 5732
rect 9036 5714 9088 5720
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 9048 4826 9076 5306
rect 9140 5302 9168 5850
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9232 5234 9260 6287
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5681 9536 6054
rect 9494 5672 9550 5681
rect 9494 5607 9550 5616
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9600 4622 9628 6734
rect 9784 6322 9812 6734
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9784 5846 9812 6258
rect 9876 5914 9904 6870
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10152 6186 10180 6394
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9784 4826 9812 5646
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9784 4146 9812 4762
rect 10060 4554 10088 6122
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 5370 10824 5510
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 10520 4282 10548 4694
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10704 4214 10732 4966
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 4214 10916 4558
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 9772 4140 9824 4146
rect 8864 4100 8984 4128
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8496 2514 8524 3334
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8588 2310 8616 3538
rect 8864 3534 8892 3946
rect 8956 3942 8984 4100
rect 9772 4082 9824 4088
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8864 3194 8892 3470
rect 8956 3194 8984 3878
rect 9876 3738 9904 3946
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9416 3058 9444 3674
rect 10060 3670 10088 3878
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 11072 3194 11100 8230
rect 11164 8090 11192 8366
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11532 7410 11560 8502
rect 11808 8430 11836 8842
rect 11992 8634 12020 8910
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11532 6934 11560 7346
rect 11520 6928 11572 6934
rect 11520 6870 11572 6876
rect 11900 6866 11928 7686
rect 11992 7002 12020 7890
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11900 6458 11928 6802
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11256 5030 11284 5714
rect 11348 5166 11376 5714
rect 12084 5710 12112 21830
rect 12268 21298 12296 22510
rect 12360 22494 12480 22522
rect 12544 23310 12664 23338
rect 12360 21486 12388 22494
rect 12440 22160 12492 22166
rect 12440 22102 12492 22108
rect 12452 21554 12480 22102
rect 12544 22030 12572 23310
rect 12624 23248 12676 23254
rect 12624 23190 12676 23196
rect 12636 23089 12664 23190
rect 12622 23080 12678 23089
rect 12622 23015 12678 23024
rect 12820 22030 12848 23666
rect 14922 23624 14978 23633
rect 14922 23559 14924 23568
rect 14976 23559 14978 23568
rect 15568 23588 15620 23594
rect 14924 23530 14976 23536
rect 15568 23530 15620 23536
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13096 22778 13124 23054
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 13096 22545 13124 22714
rect 13082 22536 13138 22545
rect 13280 22506 13308 23054
rect 14752 22778 14780 23462
rect 14936 23322 14964 23530
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15396 22778 15424 23054
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15488 22574 15516 23190
rect 15580 23118 15608 23530
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 13082 22471 13138 22480
rect 13268 22500 13320 22506
rect 13268 22442 13320 22448
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12544 21690 12572 21966
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12268 21270 12388 21298
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12176 13394 12204 14758
rect 12268 14278 12296 14826
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12268 14074 12296 14214
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12360 13814 12388 21270
rect 12544 20806 12572 21422
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12268 13786 12388 13814
rect 12268 13530 12296 13786
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12176 12782 12204 13330
rect 12544 12850 12572 14758
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 13004 14074 13032 14418
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12164 12776 12216 12782
rect 12216 12736 12296 12764
rect 12164 12718 12216 12724
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12176 11898 12204 12174
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12268 9722 12296 12736
rect 12544 12442 12572 12786
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12912 12306 12940 12650
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 13004 12170 13032 14010
rect 13096 13938 13124 14554
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13188 12442 13216 13670
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12820 11354 12848 11766
rect 13188 11558 13216 12378
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12544 10062 12572 10474
rect 12636 10198 12664 10474
rect 12728 10470 12756 11018
rect 13096 11014 13124 11290
rect 13280 11286 13308 22442
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 14200 14074 14228 22374
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15580 20058 15608 23054
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13372 13530 13400 13806
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13556 12714 13584 13330
rect 14292 12850 14320 19994
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 14292 12442 14320 12786
rect 14384 12714 14412 13126
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14384 12306 14412 12650
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13924 11626 13952 12174
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14108 11762 14136 12038
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13912 11620 13964 11626
rect 13912 11562 13964 11568
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 13096 10130 13124 10950
rect 13188 10538 13216 11018
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13188 10130 13216 10474
rect 13280 10266 13308 11222
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 13096 9722 13124 10066
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12268 9518 12296 9658
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12268 7478 12296 8026
rect 12544 7954 12572 9318
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12268 7274 12296 7414
rect 12728 7410 12756 9114
rect 13004 9042 13032 9454
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 12912 8294 12940 8978
rect 13004 8838 13032 8978
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13004 8634 13032 8774
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13188 8498 13216 8978
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11348 4826 11376 5102
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11256 4078 11284 4558
rect 11808 4146 11836 5646
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11900 4214 11928 4626
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11256 3466 11284 4014
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11532 3670 11560 3946
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 11072 2990 11100 3130
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9494 2816 9550 2825
rect 9494 2751 9550 2760
rect 9508 2650 9536 2751
rect 9968 2650 9996 2858
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8206 2000 8262 2009
rect 8206 1935 8262 1944
rect 7194 54 7328 82
rect 8390 128 8446 480
rect 8390 76 8392 128
rect 8444 76 8446 128
rect 7194 0 7250 54
rect 8390 0 8446 76
rect 9232 82 9260 2314
rect 9494 82 9550 480
rect 9232 54 9550 82
rect 9494 0 9550 54
rect 10598 82 10654 480
rect 10704 82 10732 2790
rect 11532 2582 11560 3606
rect 11624 3126 11652 3606
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 11624 2854 11652 3062
rect 12176 2961 12204 6122
rect 12268 5370 12296 7210
rect 12728 7002 12756 7346
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12360 6458 12388 6598
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12360 6118 12388 6394
rect 12728 6186 12756 6598
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12452 5234 12480 5510
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12268 4214 12296 4694
rect 12544 4690 12572 5510
rect 12728 5370 12756 5782
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12636 5098 12664 5306
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12820 5080 12848 5782
rect 12912 5234 12940 8230
rect 13464 7750 13492 8298
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 6934 13400 7142
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13372 6458 13400 6870
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12900 5092 12952 5098
rect 12820 5052 12900 5080
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12636 4078 12664 5034
rect 12820 4826 12848 5052
rect 12900 5034 12952 5040
rect 13372 5030 13400 5238
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 13372 4758 13400 4966
rect 13360 4752 13412 4758
rect 13360 4694 13412 4700
rect 13464 4622 13492 5646
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13004 4146 13032 4558
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12162 2952 12218 2961
rect 12162 2887 12218 2896
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 12360 2650 12388 3878
rect 12820 3738 12848 4082
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 13004 3670 13032 4082
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13372 3738 13400 3946
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 3194 13032 3470
rect 13372 3194 13400 3674
rect 13556 3194 13584 11562
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13832 10742 13860 10950
rect 14476 10810 14504 14418
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14568 11830 14596 12786
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15764 12306 15792 12650
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15764 11898 15792 12242
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 14280 10736 14332 10742
rect 14280 10678 14332 10684
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 9042 13676 10406
rect 13740 10266 13768 10474
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13832 9654 13860 10678
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 14016 10266 14044 10474
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14096 9920 14148 9926
rect 14292 9908 14320 10678
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14384 10470 14412 10610
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 14148 9880 14320 9908
rect 14464 9920 14516 9926
rect 14096 9862 14148 9868
rect 14464 9862 14516 9868
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 14016 9217 14044 9386
rect 14002 9208 14058 9217
rect 14002 9143 14058 9152
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 14108 8537 14136 9862
rect 14094 8528 14150 8537
rect 13728 8492 13780 8498
rect 14094 8463 14150 8472
rect 13728 8434 13780 8440
rect 13740 6798 13768 8434
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 8090 13860 8230
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13924 7546 13952 7822
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 6322 13768 6734
rect 14384 6458 14412 7210
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13740 5914 13768 6258
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 14476 5574 14504 9862
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 10066
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 14832 9648 14884 9654
rect 14832 9590 14884 9596
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14660 8634 14688 9522
rect 14844 8838 14872 9590
rect 15396 9042 15424 10202
rect 15580 10062 15608 10406
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14660 8430 14688 8570
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14568 6934 14596 7346
rect 14556 6928 14608 6934
rect 14556 6870 14608 6876
rect 14568 5778 14596 6870
rect 14660 6458 14688 8366
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14752 6905 14780 8230
rect 14844 7750 14872 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15488 8430 15516 9046
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 15844 8900 15896 8906
rect 15844 8842 15896 8848
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15658 8528 15714 8537
rect 15658 8463 15714 8472
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14844 6934 14872 7686
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 7274 15332 7890
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 14832 6928 14884 6934
rect 14738 6896 14794 6905
rect 14832 6870 14884 6876
rect 14738 6831 14794 6840
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14844 5914 14872 6870
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15198 6352 15254 6361
rect 15304 6338 15332 6666
rect 15254 6310 15332 6338
rect 15198 6287 15254 6296
rect 15212 6254 15240 6287
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 15396 5817 15424 8026
rect 15488 7954 15516 8366
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15488 7002 15516 7890
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15580 5914 15608 7210
rect 15672 6644 15700 8463
rect 15764 7857 15792 8774
rect 15856 8294 15884 8842
rect 16224 8634 16252 8910
rect 16500 8634 16528 23802
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 16868 23089 16896 23598
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 16854 23080 16910 23089
rect 16854 23015 16910 23024
rect 20088 22778 20116 23462
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 20640 22545 20668 24006
rect 20916 23866 20944 27520
rect 22848 23866 22876 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23866 24716 24210
rect 20904 23860 20956 23866
rect 20904 23802 20956 23808
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24872 23798 24900 27520
rect 25226 25120 25282 25129
rect 25226 25055 25282 25064
rect 25240 23866 25268 25055
rect 26896 24274 26924 27520
rect 26884 24268 26936 24274
rect 26884 24210 26936 24216
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 24860 23792 24912 23798
rect 24860 23734 24912 23740
rect 25240 23662 25268 23802
rect 25228 23656 25280 23662
rect 24582 23624 24638 23633
rect 25228 23598 25280 23604
rect 24582 23559 24638 23568
rect 24596 23526 24624 23559
rect 22744 23520 22796 23526
rect 22744 23462 22796 23468
rect 24584 23520 24636 23526
rect 24584 23462 24636 23468
rect 20626 22536 20682 22545
rect 20626 22471 20682 22480
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18616 12753 18644 12854
rect 18602 12744 18658 12753
rect 18602 12679 18658 12688
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 17038 9616 17094 9625
rect 17038 9551 17094 9560
rect 17052 9518 17080 9551
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16868 8294 16896 8978
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 15856 7993 15884 8230
rect 15842 7984 15898 7993
rect 15842 7919 15898 7928
rect 15750 7848 15806 7857
rect 15750 7783 15806 7792
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 6769 15884 7142
rect 15842 6760 15898 6769
rect 15842 6695 15898 6704
rect 16316 6662 16344 7278
rect 16868 6866 16896 8230
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17512 7002 17540 7890
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 15752 6656 15804 6662
rect 15672 6616 15752 6644
rect 15752 6598 15804 6604
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15568 5908 15620 5914
rect 15488 5868 15568 5896
rect 15382 5808 15438 5817
rect 14556 5772 14608 5778
rect 15382 5743 15438 5752
rect 14556 5714 14608 5720
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 10598 54 10732 82
rect 11624 82 11652 2314
rect 11702 82 11758 480
rect 11624 54 11758 82
rect 12728 82 12756 3062
rect 13372 2904 13400 3130
rect 13452 2916 13504 2922
rect 13372 2876 13452 2904
rect 13372 2650 13400 2876
rect 13452 2858 13504 2864
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 12806 82 12862 480
rect 12728 54 12862 82
rect 13648 82 13676 4490
rect 14292 3534 14320 4966
rect 14568 4826 14596 5714
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14384 3942 14412 4558
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14660 4010 14688 4150
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3641 14412 3878
rect 14660 3641 14688 3946
rect 14370 3632 14426 3641
rect 14370 3567 14426 3576
rect 14646 3632 14702 3641
rect 14646 3567 14702 3576
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14752 3058 14780 4762
rect 15304 4690 15332 5306
rect 15488 5234 15516 5868
rect 15568 5850 15620 5856
rect 15672 5778 15700 6190
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15396 4690 15424 5102
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14844 2514 14872 3402
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 13910 82 13966 480
rect 13648 54 13966 82
rect 10598 0 10654 54
rect 11702 0 11758 54
rect 12806 0 12862 54
rect 13910 0 13966 54
rect 15106 82 15162 480
rect 15304 82 15332 4490
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15396 3194 15424 3470
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15488 2582 15516 3470
rect 15476 2576 15528 2582
rect 15476 2518 15528 2524
rect 15580 2514 15608 5646
rect 15672 5370 15700 5714
rect 15764 5642 15792 6598
rect 16316 6254 16344 6598
rect 16868 6458 16896 6802
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 17236 6390 17264 6598
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15856 5681 15884 6054
rect 16316 5914 16344 6190
rect 17328 5914 17356 6802
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 15842 5672 15898 5681
rect 15752 5636 15804 5642
rect 15842 5607 15898 5616
rect 15752 5578 15804 5584
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 15844 4752 15896 4758
rect 15844 4694 15896 4700
rect 15752 4004 15804 4010
rect 15752 3946 15804 3952
rect 15764 3738 15792 3946
rect 15856 3942 15884 4694
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 16408 4146 16436 4422
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 15672 3194 15700 3606
rect 15764 3398 15792 3674
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15856 1601 15884 3878
rect 16316 3670 16344 3946
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 15948 2650 15976 2790
rect 15936 2644 15988 2650
rect 16212 2644 16264 2650
rect 15988 2604 16212 2632
rect 15936 2586 15988 2592
rect 16212 2586 16264 2592
rect 15842 1592 15898 1601
rect 15842 1527 15898 1536
rect 15106 54 15332 82
rect 16210 82 16266 480
rect 16408 82 16436 3946
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16500 3058 16528 3402
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16488 2916 16540 2922
rect 16592 2904 16620 3130
rect 17052 3058 17080 4218
rect 17236 3942 17264 4626
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17328 3194 17356 3538
rect 17420 3194 17448 3878
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16540 2876 16620 2904
rect 16488 2858 16540 2864
rect 16592 2582 16620 2876
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16684 2446 16712 2994
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 17512 2310 17540 3878
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 16210 54 16436 82
rect 17314 82 17370 480
rect 17604 82 17632 3946
rect 17880 3097 17908 5102
rect 18064 3398 18092 9318
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 22112 8362 22140 19110
rect 22756 16017 22784 23462
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 25134 20496 25190 20505
rect 25134 20431 25190 20440
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 25148 19514 25176 20431
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25148 19310 25176 19450
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 22742 16008 22798 16017
rect 22742 15943 22798 15952
rect 25134 15872 25190 15881
rect 25134 15807 25190 15816
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 25148 15162 25176 15807
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25148 14958 25176 15098
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 23848 14544 23900 14550
rect 23848 14486 23900 14492
rect 23860 13734 23888 14486
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24688 13814 24716 13874
rect 24688 13786 24808 13814
rect 24872 13802 24900 14350
rect 25148 14346 25176 14758
rect 25136 14340 25188 14346
rect 25136 14282 25188 14288
rect 25148 14074 25176 14282
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 23860 13394 23888 13670
rect 24044 13530 24072 13670
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23860 12850 23888 13330
rect 24780 13172 24808 13786
rect 24860 13796 24912 13802
rect 24860 13738 24912 13744
rect 24872 13433 24900 13738
rect 24858 13424 24914 13433
rect 24858 13359 24914 13368
rect 24860 13184 24912 13190
rect 24780 13144 24860 13172
rect 24860 13126 24912 13132
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23860 12753 23888 12786
rect 23846 12744 23902 12753
rect 23846 12679 23902 12688
rect 24214 12336 24270 12345
rect 24214 12271 24270 12280
rect 24228 11898 24256 12271
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 24872 7002 24900 13126
rect 27618 11656 27674 11665
rect 27618 11591 27674 11600
rect 27632 11558 27660 11591
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27618 7032 27674 7041
rect 24860 6996 24912 7002
rect 27618 6967 27674 6976
rect 24860 6938 24912 6944
rect 27632 6934 27660 6967
rect 27620 6928 27672 6934
rect 27620 6870 27672 6876
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6458 24716 6802
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18708 6225 18736 6258
rect 18694 6216 18750 6225
rect 18694 6151 18750 6160
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19260 5166 19288 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20916 5370 20944 5714
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 21548 5296 21600 5302
rect 21548 5238 21600 5244
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18432 4690 18460 4966
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 18420 4684 18472 4690
rect 18420 4626 18472 4632
rect 18432 4282 18460 4626
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 17972 3126 18000 3334
rect 17960 3120 18012 3126
rect 17866 3088 17922 3097
rect 17960 3062 18012 3068
rect 17866 3023 17922 3032
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 17314 54 17632 82
rect 18418 82 18474 480
rect 18708 82 18736 2382
rect 18892 134 18920 4422
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20902 3632 20958 3641
rect 19064 3596 19116 3602
rect 20902 3567 20958 3576
rect 19064 3538 19116 3544
rect 19076 3126 19104 3538
rect 20260 3460 20312 3466
rect 20260 3402 20312 3408
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 19536 2514 19564 3334
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20180 2650 20208 2790
rect 20272 2650 20300 3402
rect 20916 2854 20944 3567
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 19524 2508 19576 2514
rect 19524 2450 19576 2456
rect 19708 2304 19760 2310
rect 19708 2246 19760 2252
rect 21456 2304 21508 2310
rect 21456 2246 21508 2252
rect 18418 54 18736 82
rect 18880 128 18932 134
rect 18880 70 18932 76
rect 19522 82 19578 480
rect 19720 82 19748 2246
rect 21468 1873 21496 2246
rect 21454 1864 21510 1873
rect 21454 1799 21510 1808
rect 19522 54 19748 82
rect 20626 128 20682 480
rect 20626 76 20628 128
rect 20680 76 20682 128
rect 15106 0 15162 54
rect 16210 0 16266 54
rect 17314 0 17370 54
rect 18418 0 18474 54
rect 19522 0 19578 54
rect 20626 0 20682 76
rect 21560 82 21588 5238
rect 21822 82 21878 480
rect 21560 54 21878 82
rect 22848 82 22876 5510
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 23848 2916 23900 2922
rect 23848 2858 23900 2864
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 23216 2009 23244 2246
rect 23202 2000 23258 2009
rect 23202 1935 23258 1944
rect 22926 82 22982 480
rect 22848 54 22982 82
rect 23860 82 23888 2858
rect 25964 2848 26016 2854
rect 25964 2790 26016 2796
rect 24860 2576 24912 2582
rect 24860 2518 24912 2524
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24030 82 24086 480
rect 23860 54 24086 82
rect 24872 82 24900 2518
rect 25134 82 25190 480
rect 24872 54 25190 82
rect 25976 82 26004 2790
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 26238 82 26294 480
rect 25976 54 26294 82
rect 27080 82 27108 2246
rect 27342 82 27398 480
rect 27080 54 27398 82
rect 21822 0 21878 54
rect 22926 0 22982 54
rect 24030 0 24086 54
rect 25134 0 25190 54
rect 26238 0 26294 54
rect 27342 0 27398 54
<< via2 >>
rect 3146 24928 3202 24984
rect 1214 20032 1270 20088
rect 1582 23432 1638 23488
rect 1582 21664 1638 21720
rect 1398 15544 1454 15600
rect 1582 15136 1638 15192
rect 2962 17176 3018 17232
rect 3146 16768 3202 16824
rect 1214 8472 1270 8528
rect 110 7384 166 7440
rect 1398 5208 1454 5264
rect 110 4120 166 4176
rect 3054 11192 3110 11248
rect 2318 7792 2374 7848
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 3974 18400 4030 18456
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 8298 26560 8354 26616
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 3974 11736 4030 11792
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 3514 6160 3570 6216
rect 3422 4120 3478 4176
rect 3238 3848 3294 3904
rect 2778 3032 2834 3088
rect 2318 1400 2374 1456
rect 4802 9560 4858 9616
rect 4250 4256 4306 4312
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6182 12280 6238 12336
rect 6734 13368 6790 13424
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 4894 6840 4950 6896
rect 4894 4256 4950 4312
rect 5814 7792 5870 7848
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 6550 7948 6606 7984
rect 6550 7928 6552 7948
rect 6552 7928 6604 7948
rect 6604 7928 6606 7948
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5722 5752 5778 5808
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 4526 2896 4582 2952
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6458 3884 6460 3904
rect 6460 3884 6512 3904
rect 6512 3884 6514 3904
rect 6458 3848 6514 3884
rect 7102 3712 7158 3768
rect 7010 3576 7066 3632
rect 4894 2760 4950 2816
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7838 4120 7894 4176
rect 7654 3032 7710 3088
rect 7194 1808 7250 1864
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 11242 17176 11298 17232
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10690 15952 10746 16008
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 8390 7928 8446 7984
rect 8574 6296 8630 6352
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 11518 13368 11574 13424
rect 9126 6704 9182 6760
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 11242 9152 11298 9208
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 9218 6296 9274 6352
rect 9494 5616 9550 5672
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 12622 23024 12678 23080
rect 14922 23588 14978 23624
rect 14922 23568 14924 23588
rect 14924 23568 14976 23588
rect 14976 23568 14978 23588
rect 13082 22480 13138 22536
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 9494 2760 9550 2816
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 8206 1944 8262 2000
rect 12162 2896 12218 2952
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14002 9152 14058 9208
rect 14094 8472 14150 8528
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15658 8472 15714 8528
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14738 6840 14794 6896
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15198 6296 15254 6352
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 16854 23024 16910 23080
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 25226 25064 25282 25120
rect 24582 23568 24638 23624
rect 20626 22480 20682 22536
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 18602 12688 18658 12744
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 17038 9560 17094 9616
rect 15842 7928 15898 7984
rect 15750 7792 15806 7848
rect 15842 6704 15898 6760
rect 15382 5752 15438 5808
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14370 3576 14426 3632
rect 14646 3576 14702 3632
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15842 5616 15898 5672
rect 15842 1536 15898 1592
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 25134 20440 25190 20496
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 22742 15952 22798 16008
rect 25134 15816 25190 15872
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24858 13368 24914 13424
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 23846 12688 23902 12744
rect 24214 12280 24270 12336
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 27618 11600 27674 11656
rect 27618 6976 27674 7032
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 18694 6160 18750 6216
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 17866 3032 17922 3088
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20902 3576 20958 3632
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 21454 1808 21510 1864
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 23202 1944 23258 2000
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
<< metal3 >>
rect 0 27072 480 27192
rect 62 26618 122 27072
rect 8293 26618 8359 26621
rect 62 26616 8359 26618
rect 62 26560 8298 26616
rect 8354 26560 8359 26616
rect 62 26558 8359 26560
rect 8293 26555 8359 26558
rect 10277 25600 10597 25601
rect 0 25440 480 25560
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 27520 25576 28000 25696
rect 19610 25535 19930 25536
rect 62 24986 122 25440
rect 25221 25122 25287 25125
rect 27662 25122 27722 25576
rect 25221 25120 27722 25122
rect 25221 25064 25226 25120
rect 25282 25064 27722 25120
rect 25221 25062 27722 25064
rect 25221 25059 25287 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 3141 24986 3207 24989
rect 62 24984 3207 24986
rect 62 24928 3146 24984
rect 3202 24928 3207 24984
rect 62 24926 3207 24928
rect 3141 24923 3207 24926
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 5610 23968 5930 23969
rect 0 23808 480 23928
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 62 23490 122 23808
rect 14917 23626 14983 23629
rect 24577 23626 24643 23629
rect 14917 23624 24643 23626
rect 14917 23568 14922 23624
rect 14978 23568 24582 23624
rect 24638 23568 24643 23624
rect 14917 23566 24643 23568
rect 14917 23563 14983 23566
rect 24577 23563 24643 23566
rect 1577 23490 1643 23493
rect 62 23488 1643 23490
rect 62 23432 1582 23488
rect 1638 23432 1643 23488
rect 62 23430 1643 23432
rect 1577 23427 1643 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 12617 23082 12683 23085
rect 16849 23082 16915 23085
rect 12617 23080 16915 23082
rect 12617 23024 12622 23080
rect 12678 23024 16854 23080
rect 16910 23024 16915 23080
rect 12617 23022 16915 23024
rect 12617 23019 12683 23022
rect 16849 23019 16915 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 13077 22538 13143 22541
rect 20621 22538 20687 22541
rect 13077 22536 20687 22538
rect 13077 22480 13082 22536
rect 13138 22480 20626 22536
rect 20682 22480 20687 22536
rect 13077 22478 20687 22480
rect 13077 22475 13143 22478
rect 20621 22475 20687 22478
rect 10277 22336 10597 22337
rect 0 22176 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 62 21722 122 22176
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 1577 21722 1643 21725
rect 62 21720 1643 21722
rect 62 21664 1582 21720
rect 1638 21664 1643 21720
rect 62 21662 1643 21664
rect 1577 21659 1643 21662
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 27520 20952 28000 21072
rect 5610 20704 5930 20705
rect 0 20544 480 20664
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 62 20090 122 20544
rect 25129 20498 25195 20501
rect 27662 20498 27722 20952
rect 25129 20496 27722 20498
rect 25129 20440 25134 20496
rect 25190 20440 27722 20496
rect 25129 20438 27722 20440
rect 25129 20435 25195 20438
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1209 20090 1275 20093
rect 62 20088 1275 20090
rect 62 20032 1214 20088
rect 1270 20032 1275 20088
rect 62 20030 1275 20032
rect 1209 20027 1275 20030
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 10277 19072 10597 19073
rect 0 18912 480 19032
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 62 18458 122 18912
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 3969 18458 4035 18461
rect 62 18456 4035 18458
rect 62 18400 3974 18456
rect 4030 18400 4035 18456
rect 62 18398 4035 18400
rect 3969 18395 4035 18398
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 5610 17440 5930 17441
rect 0 17280 480 17400
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 62 16826 122 17280
rect 2957 17234 3023 17237
rect 11237 17234 11303 17237
rect 2957 17232 11303 17234
rect 2957 17176 2962 17232
rect 3018 17176 11242 17232
rect 11298 17176 11303 17232
rect 2957 17174 11303 17176
rect 2957 17171 3023 17174
rect 11237 17171 11303 17174
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 3141 16826 3207 16829
rect 62 16824 3207 16826
rect 62 16768 3146 16824
rect 3202 16768 3207 16824
rect 62 16766 3207 16768
rect 3141 16763 3207 16766
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 27520 16328 28000 16448
rect 24277 16287 24597 16288
rect 10685 16010 10751 16013
rect 22737 16010 22803 16013
rect 10685 16008 22803 16010
rect 10685 15952 10690 16008
rect 10746 15952 22742 16008
rect 22798 15952 22803 16008
rect 10685 15950 22803 15952
rect 10685 15947 10751 15950
rect 22737 15947 22803 15950
rect 25129 15874 25195 15877
rect 27662 15874 27722 16328
rect 25129 15872 27722 15874
rect 25129 15816 25134 15872
rect 25190 15816 27722 15872
rect 25129 15814 27722 15816
rect 25129 15811 25195 15814
rect 10277 15808 10597 15809
rect 0 15648 480 15768
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 62 15194 122 15648
rect 1393 15602 1459 15605
rect 1894 15602 1900 15604
rect 1393 15600 1900 15602
rect 1393 15544 1398 15600
rect 1454 15544 1900 15600
rect 1393 15542 1900 15544
rect 1393 15539 1459 15542
rect 1894 15540 1900 15542
rect 1964 15540 1970 15604
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 1577 15194 1643 15197
rect 62 15192 1643 15194
rect 62 15136 1582 15192
rect 1638 15136 1643 15192
rect 62 15134 1643 15136
rect 1577 15131 1643 15134
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13880 480 14000
rect 62 13426 122 13880
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 6729 13426 6795 13429
rect 62 13424 6795 13426
rect 62 13368 6734 13424
rect 6790 13368 6795 13424
rect 62 13366 6795 13368
rect 6729 13363 6795 13366
rect 11513 13426 11579 13429
rect 24853 13426 24919 13429
rect 11513 13424 24919 13426
rect 11513 13368 11518 13424
rect 11574 13368 24858 13424
rect 24914 13368 24919 13424
rect 11513 13366 24919 13368
rect 11513 13363 11579 13366
rect 24853 13363 24919 13366
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 18597 12746 18663 12749
rect 23841 12746 23907 12749
rect 18597 12744 23907 12746
rect 18597 12688 18602 12744
rect 18658 12688 23846 12744
rect 23902 12688 23907 12744
rect 18597 12686 23907 12688
rect 18597 12683 18663 12686
rect 23841 12683 23907 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 0 12248 480 12368
rect 6177 12338 6243 12341
rect 24209 12338 24275 12341
rect 6177 12336 24275 12338
rect 6177 12280 6182 12336
rect 6238 12280 24214 12336
rect 24270 12280 24275 12336
rect 6177 12278 24275 12280
rect 6177 12275 6243 12278
rect 24209 12275 24275 12278
rect 62 11794 122 12248
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 3969 11794 4035 11797
rect 62 11792 4035 11794
rect 62 11736 3974 11792
rect 4030 11736 4035 11792
rect 62 11734 4035 11736
rect 3969 11731 4035 11734
rect 27520 11656 28000 11688
rect 27520 11600 27618 11656
rect 27674 11600 28000 11656
rect 27520 11568 28000 11600
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3049 11250 3115 11253
rect 62 11248 3115 11250
rect 62 11192 3054 11248
rect 3110 11192 3115 11248
rect 62 11190 3115 11192
rect 62 10736 122 11190
rect 3049 11187 3115 11190
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10616 480 10736
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 4797 9618 4863 9621
rect 17033 9618 17099 9621
rect 4797 9616 17099 9618
rect 4797 9560 4802 9616
rect 4858 9560 17038 9616
rect 17094 9560 17099 9616
rect 4797 9558 17099 9560
rect 4797 9555 4863 9558
rect 17033 9555 17099 9558
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 11237 9210 11303 9213
rect 13997 9210 14063 9213
rect 11237 9208 14063 9210
rect 11237 9152 11242 9208
rect 11298 9152 14002 9208
rect 14058 9152 14063 9208
rect 11237 9150 14063 9152
rect 11237 9147 11303 9150
rect 13997 9147 14063 9150
rect 0 8984 480 9104
rect 62 8530 122 8984
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 1209 8530 1275 8533
rect 14089 8530 14155 8533
rect 15653 8530 15719 8533
rect 62 8528 1275 8530
rect 62 8472 1214 8528
rect 1270 8472 1275 8528
rect 62 8470 1275 8472
rect 13962 8528 15719 8530
rect 13962 8472 14094 8528
rect 14150 8472 15658 8528
rect 15714 8472 15719 8528
rect 13962 8470 15719 8472
rect 1209 8467 1275 8470
rect 14089 8467 14155 8470
rect 15653 8467 15719 8470
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 6545 7986 6611 7989
rect 8385 7986 8451 7989
rect 15837 7986 15903 7989
rect 6545 7984 15903 7986
rect 6545 7928 6550 7984
rect 6606 7928 8390 7984
rect 8446 7928 15842 7984
rect 15898 7928 15903 7984
rect 6545 7926 15903 7928
rect 6545 7923 6611 7926
rect 8385 7923 8451 7926
rect 15837 7923 15903 7926
rect 2313 7850 2379 7853
rect 5809 7850 5875 7853
rect 15745 7850 15811 7853
rect 2313 7848 15811 7850
rect 2313 7792 2318 7848
rect 2374 7792 5814 7848
rect 5870 7792 15750 7848
rect 15806 7792 15811 7848
rect 2313 7790 15811 7792
rect 2313 7787 2379 7790
rect 5809 7787 5875 7790
rect 15745 7787 15811 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 0 7440 480 7472
rect 0 7384 110 7440
rect 166 7384 480 7440
rect 0 7352 480 7384
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 27520 7032 28000 7064
rect 27520 6976 27618 7032
rect 27674 6976 28000 7032
rect 27520 6944 28000 6976
rect 4889 6898 4955 6901
rect 14733 6898 14799 6901
rect 4889 6896 14799 6898
rect 4889 6840 4894 6896
rect 4950 6840 14738 6896
rect 14794 6840 14799 6896
rect 4889 6838 14799 6840
rect 4889 6835 4955 6838
rect 14733 6835 14799 6838
rect 9121 6762 9187 6765
rect 15837 6762 15903 6765
rect 9121 6760 15903 6762
rect 9121 6704 9126 6760
rect 9182 6704 15842 6760
rect 15898 6704 15903 6760
rect 9121 6702 15903 6704
rect 9121 6699 9187 6702
rect 15837 6699 15903 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 8569 6354 8635 6357
rect 9213 6354 9279 6357
rect 15193 6354 15259 6357
rect 8569 6352 15259 6354
rect 8569 6296 8574 6352
rect 8630 6296 9218 6352
rect 9274 6296 15198 6352
rect 15254 6296 15259 6352
rect 8569 6294 15259 6296
rect 8569 6291 8635 6294
rect 9213 6291 9279 6294
rect 15193 6291 15259 6294
rect 3509 6218 3575 6221
rect 18689 6218 18755 6221
rect 3509 6216 18755 6218
rect 3509 6160 3514 6216
rect 3570 6160 18694 6216
rect 18750 6160 18755 6216
rect 3509 6158 18755 6160
rect 3509 6155 3575 6158
rect 18689 6155 18755 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 0 5720 480 5840
rect 5717 5810 5783 5813
rect 15377 5810 15443 5813
rect 5717 5808 15443 5810
rect 5717 5752 5722 5808
rect 5778 5752 15382 5808
rect 15438 5752 15443 5808
rect 5717 5750 15443 5752
rect 5717 5747 5783 5750
rect 15377 5747 15443 5750
rect 62 5266 122 5720
rect 9489 5674 9555 5677
rect 15837 5674 15903 5677
rect 9489 5672 15903 5674
rect 9489 5616 9494 5672
rect 9550 5616 15842 5672
rect 15898 5616 15903 5672
rect 9489 5614 15903 5616
rect 9489 5611 9555 5614
rect 15837 5611 15903 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 1393 5266 1459 5269
rect 62 5264 1459 5266
rect 62 5208 1398 5264
rect 1454 5208 1459 5264
rect 62 5206 1459 5208
rect 1393 5203 1459 5206
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 4245 4314 4311 4317
rect 4889 4314 4955 4317
rect 4245 4312 4955 4314
rect 4245 4256 4250 4312
rect 4306 4256 4894 4312
rect 4950 4256 4955 4312
rect 4245 4254 4955 4256
rect 4245 4251 4311 4254
rect 4889 4251 4955 4254
rect 0 4176 480 4208
rect 0 4120 110 4176
rect 166 4120 480 4176
rect 0 4088 480 4120
rect 3417 4178 3483 4181
rect 7833 4178 7899 4181
rect 3417 4176 7899 4178
rect 3417 4120 3422 4176
rect 3478 4120 7838 4176
rect 7894 4120 7899 4176
rect 3417 4118 7899 4120
rect 3417 4115 3483 4118
rect 7833 4115 7899 4118
rect 3233 3906 3299 3909
rect 6453 3906 6519 3909
rect 3233 3904 6519 3906
rect 3233 3848 3238 3904
rect 3294 3848 6458 3904
rect 6514 3848 6519 3904
rect 3233 3846 6519 3848
rect 3233 3843 3299 3846
rect 6453 3843 6519 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 1894 3708 1900 3772
rect 1964 3770 1970 3772
rect 7097 3770 7163 3773
rect 1964 3768 7163 3770
rect 1964 3712 7102 3768
rect 7158 3712 7163 3768
rect 1964 3710 7163 3712
rect 1964 3708 1970 3710
rect 7097 3707 7163 3710
rect 7005 3634 7071 3637
rect 14365 3634 14431 3637
rect 7005 3632 14431 3634
rect 7005 3576 7010 3632
rect 7066 3576 14370 3632
rect 14426 3576 14431 3632
rect 7005 3574 14431 3576
rect 7005 3571 7071 3574
rect 14365 3571 14431 3574
rect 14641 3634 14707 3637
rect 20897 3634 20963 3637
rect 14641 3632 20963 3634
rect 14641 3576 14646 3632
rect 14702 3576 20902 3632
rect 20958 3576 20963 3632
rect 14641 3574 20963 3576
rect 14641 3571 14707 3574
rect 20897 3571 20963 3574
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 2773 3090 2839 3093
rect 62 3088 2839 3090
rect 62 3032 2778 3088
rect 2834 3032 2839 3088
rect 62 3030 2839 3032
rect 62 2576 122 3030
rect 2773 3027 2839 3030
rect 7649 3090 7715 3093
rect 17861 3090 17927 3093
rect 7649 3088 17927 3090
rect 7649 3032 7654 3088
rect 7710 3032 17866 3088
rect 17922 3032 17927 3088
rect 7649 3030 17927 3032
rect 7649 3027 7715 3030
rect 17861 3027 17927 3030
rect 4521 2954 4587 2957
rect 12157 2954 12223 2957
rect 4521 2952 12223 2954
rect 4521 2896 4526 2952
rect 4582 2896 12162 2952
rect 12218 2896 12223 2952
rect 4521 2894 12223 2896
rect 4521 2891 4587 2894
rect 12157 2891 12223 2894
rect 4889 2818 4955 2821
rect 9489 2818 9555 2821
rect 4889 2816 9555 2818
rect 4889 2760 4894 2816
rect 4950 2760 9494 2816
rect 9550 2760 9555 2816
rect 4889 2758 9555 2760
rect 4889 2755 4955 2758
rect 9489 2755 9555 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 0 2456 480 2576
rect 27520 2320 28000 2440
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 8201 2002 8267 2005
rect 23197 2002 23263 2005
rect 8201 2000 23263 2002
rect 8201 1944 8206 2000
rect 8262 1944 23202 2000
rect 23258 1944 23263 2000
rect 8201 1942 23263 1944
rect 8201 1939 8267 1942
rect 23197 1939 23263 1942
rect 7189 1866 7255 1869
rect 21449 1866 21515 1869
rect 7189 1864 21515 1866
rect 7189 1808 7194 1864
rect 7250 1808 21454 1864
rect 21510 1808 21515 1864
rect 7189 1806 21515 1808
rect 7189 1803 7255 1806
rect 21449 1803 21515 1806
rect 15837 1594 15903 1597
rect 27662 1594 27722 2320
rect 15837 1592 27722 1594
rect 15837 1536 15842 1592
rect 15898 1536 27722 1592
rect 15837 1534 27722 1536
rect 15837 1531 15903 1534
rect 2313 1458 2379 1461
rect 62 1456 2379 1458
rect 62 1400 2318 1456
rect 2374 1400 2379 1456
rect 62 1398 2379 1400
rect 62 944 122 1398
rect 2313 1395 2379 1398
rect 0 824 480 944
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 1900 15540 1964 15604
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 1900 3708 1964 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 1899 15604 1965 15605
rect 1899 15540 1900 15604
rect 1964 15540 1965 15604
rect 1899 15539 1965 15540
rect 1902 3773 1962 15539
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 1899 3772 1965 3773
rect 1899 3708 1900 3772
rect 1964 3708 1965 3772
rect 1899 3707 1965 3708
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_fill_1  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_13
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_nand2_4  _126_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1472 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_17
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__D
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_21
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _125_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _086_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_82
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _204_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 406 592
use scs8hd_conb_1  _187_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9936 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 1050 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_109
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_101 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_117 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_121
timestamp 1586364061
transform 1 0 12236 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_135
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 1050 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_144
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_148
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_156
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_160
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_172
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_176 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _102_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _213_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_204
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_215
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_219 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_231
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_243
timestamp 1586364061
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24288 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_251
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_255
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_259
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_271
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 590 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_35
timestamp 1586364061
transform 1 0 4324 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_40
timestamp 1586364061
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_73
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_77
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_121
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_140
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_4  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_4  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_8  _092_
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_180
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_197
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_nand2_4  _148_
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_or4_4  _123_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__C
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_33
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_47
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 314 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_56
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_60
timestamp 1586364061
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_65
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_69
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_85
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_89
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_102
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_106
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_113
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_155
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_182
timestamp 1586364061
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_187
timestamp 1586364061
transform 1 0 18308 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_191
timestamp 1586364061
transform 1 0 18676 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_198
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_202
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_226
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _173_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 406 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_6  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 590 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__C
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_109
timestamp 1586364061
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 11316 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_139
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_148
timestamp 1586364061
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_175
timestamp 1586364061
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _211_
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_187
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_195
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_207
timestamp 1586364061
transform 1 0 20148 0 -1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _111_
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_18
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_35
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _107_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_or4_4  _133_
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_78
timestamp 1586364061
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_91
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 774 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_134
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_151
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 314 592
use scs8hd_inv_8  _091_
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_172
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_180
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_187
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_203
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_217
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_241
timestamp 1586364061
transform 1 0 23276 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_14
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_18
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _085_
timestamp 1586364061
transform 1 0 4140 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_42
timestamp 1586364061
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_48
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_52
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_69
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_69
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_65
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use scs8hd_or2_4  _121_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 682 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_73
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__D
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 866 592
use scs8hd_conb_1  _194_
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_100
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_104
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_109
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_3  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_134
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_155
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_168
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_173
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_174
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__C
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__D
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_192
timestamp 1586364061
transform 1 0 18768 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_200
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_219
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_212
timestamp 1586364061
transform 1 0 20608 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_231
timestamp 1586364061
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_224
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_243
timestamp 1586364061
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_255
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_253
timestamp 1586364061
transform 1 0 24380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_267
timestamp 1586364061
transform 1 0 25668 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_38
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_52
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _193_
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_73
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_77
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_8  _114_
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_115
timestamp 1586364061
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_128
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_132
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__D
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _155_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _158_
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_4  FILLER_8_167
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_180
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_192
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_212
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_258
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_270
timestamp 1586364061
transform 1 0 25944 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_14
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_28
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 866 592
use scs8hd_decap_6  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use scs8hd_inv_8  _106_
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_78
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_151
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_18
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_26
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _108_
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_38
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_48
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_52
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_8  _105_
timestamp 1586364061
transform 1 0 9752 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_138
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_142
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_150
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_175
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_187
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_199
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_inv_8  _112_
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__C
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_65
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 314 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_83
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use scs8hd_or4_4  _167_
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__167__D
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_100
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_111
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_131
timestamp 1586364061
transform 1 0 13156 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_141
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_158
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_162
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_169
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_177
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_16
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_20
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_24
timestamp 1586364061
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_28
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_35
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 590 592
use scs8hd_nor3_4  _177_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 1234 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_75
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_79
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__D
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_98
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_121
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 774 592
use scs8hd_conb_1  _192_
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_151
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_or4_4  _164_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_175
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_187
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_11
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_or4_4  _152_
timestamp 1586364061
transform 1 0 2300 0 -1 10336
box -38 -48 866 592
use scs8hd_or2_4  _122_
timestamp 1586364061
transform 1 0 1472 0 1 9248
box -38 -48 682 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_26
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_38
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _120_
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_48
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_58
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_8  _119_
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 866 592
use scs8hd_or4_4  _127_
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_82
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__C
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__D
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_86
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_115
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_111
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _099_
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_8  _087_
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_149
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_150
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_157
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_169
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_181
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_193
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 1050 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__D
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_20
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_24
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _103_
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__C
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_52
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_56
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 314 592
use scs8hd_or4_4  _136_
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__C
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_90
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _170_
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 774 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_172
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_180
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_16
timestamp 1586364061
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_20
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_28
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_35
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_39
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 222 592
use scs8hd_nor3_4  _176_
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 1234 592
use scs8hd_decap_3  FILLER_16_43
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_76
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 590 592
use scs8hd_or4_4  _145_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__D
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_16_123
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_127
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_140
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_24
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_nor3_4  _175_
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_28
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_45
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_49
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_83
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_90
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_129
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_133
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_146
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 774 592
use scs8hd_conb_1  _195_
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_157
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_253
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_262
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_17_274
timestamp 1586364061
transform 1 0 26312 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_inv_8  _104_
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_14
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_18
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_26
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 314 592
use scs8hd_nor3_4  _174_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__142__D
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 130 592
use scs8hd_or4_4  _142_
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__C
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_71
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_146
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_8  _093_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_187
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_8  _110_
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_17
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_28
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_47
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 590 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_79
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 590 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_95
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 774 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_139
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_163
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _116_
timestamp 1586364061
transform 1 0 23736 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_249
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_245
timestamp 1586364061
transform 1 0 23644 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24748 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_261
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_255
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_273
timestamp 1586364061
transform 1 0 26220 0 1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 1050 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_29
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_33
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_46
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_50
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_54
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_81
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_128
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_259
timestamp 1586364061
transform 1 0 24932 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_263
timestamp 1586364061
transform 1 0 25300 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_21_275
timestamp 1586364061
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_48
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_22_60
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_72
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_86
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_258
timestamp 1586364061
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_270
timestamp 1586364061
transform 1 0 25944 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_9
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_19
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_29
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_42
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_46
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 590 592
use scs8hd_inv_8  _096_
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  FILLER_23_94
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_156
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_168
timestamp 1586364061
transform 1 0 16560 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_253
timestamp 1586364061
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_262
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_23_274
timestamp 1586364061
transform 1 0 26312 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_16
timestamp 1586364061
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_20
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_8  _117_
timestamp 1586364061
transform 1 0 4324 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_28
timestamp 1586364061
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_4  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_69
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 8188 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_73
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_8  _098_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_8  _115_
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_143
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_16
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_20
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 406 592
use scs8hd_inv_8  _118_
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__D
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_45
timestamp 1586364061
transform 1 0 5244 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_49
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_81
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_88
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _180_
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_105
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_116
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 590 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_inv_8  _109_
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_10
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_16
timestamp 1586364061
transform 1 0 2576 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_20
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_21
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_25
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_32
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_28
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 1142 592
use scs8hd_or4_4  _161_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_45
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_53
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_27_52
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 774 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_59
timestamp 1586364061
transform 1 0 6532 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_76
timestamp 1586364061
transform 1 0 8096 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_76
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_80
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_84
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_88
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _097_
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_105
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_120
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_143
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_151
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_17
timestamp 1586364061
transform 1 0 2668 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_29
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_35
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_47
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_59
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_67
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_12  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_114
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_126
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_138
timestamp 1586364061
transform 1 0 13800 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_28_150
timestamp 1586364061
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _163_
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_17
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_21
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_33
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_45
timestamp 1586364061
transform 1 0 5244 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_94
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_103
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_29_115
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1472 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_6
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_10
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_22
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_34
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_46
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_58
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_258
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_262
timestamp 1586364061
transform 1 0 25208 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_31_274
timestamp 1586364061
transform 1 0 26312 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_35
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_47
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_137
timestamp 1586364061
transform 1 0 13708 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 590 592
use scs8hd_inv_8  _088_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_144
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12328 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_115
timestamp 1586364061
transform 1 0 11684 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_121
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_131
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_143
timestamp 1586364061
transform 1 0 14260 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_151
timestamp 1586364061
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_23
timestamp 1586364061
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_35
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_47
timestamp 1586364061
transform 1 0 5428 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_80
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_83
timestamp 1586364061
transform 1 0 8740 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 774 592
use scs8hd_inv_8  _100_
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_132
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_136
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_140
timestamp 1586364061
transform 1 0 13984 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_154
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_158
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_162
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_174
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_182
timestamp 1586364061
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_116
timestamp 1586364061
transform 1 0 11776 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_133
timestamp 1586364061
transform 1 0 13340 0 -1 23392
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_151
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_175
timestamp 1586364061
transform 1 0 17204 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_187
timestamp 1586364061
transform 1 0 18308 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_199
timestamp 1586364061
transform 1 0 19412 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_211
timestamp 1586364061
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 2944 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2760 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_24
timestamp 1586364061
transform 1 0 3312 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_21
timestamp 1586364061
transform 1 0 3036 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_28
timestamp 1586364061
transform 1 0 3680 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_37
timestamp 1586364061
transform 1 0 4508 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_41
timestamp 1586364061
transform 1 0 4876 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_40_29
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_39_70
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_78
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_84
timestamp 1586364061
transform 1 0 8832 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_88
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_96
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_100
timestamp 1586364061
transform 1 0 10304 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_112
timestamp 1586364061
transform 1 0 11408 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_120
timestamp 1586364061
transform 1 0 12144 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_119
timestamp 1586364061
transform 1 0 12052 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_136
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_131
timestamp 1586364061
transform 1 0 13156 0 -1 24480
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_144
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_143
timestamp 1586364061
transform 1 0 14260 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_151
timestamp 1586364061
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_2  _212_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_162
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_158
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_170
timestamp 1586364061
transform 1 0 16744 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_182
timestamp 1586364061
transform 1 0 17848 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18952 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_197
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_201
timestamp 1586364061
transform 1 0 19596 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_194
timestamp 1586364061
transform 1 0 18952 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_206
timestamp 1586364061
transform 1 0 20056 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_213
timestamp 1586364061
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_218
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_222
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_234
timestamp 1586364061
transform 1 0 22632 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_242
timestamp 1586364061
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_248
timestamp 1586364061
transform 1 0 23920 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_252
timestamp 1586364061
transform 1 0 24288 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_258
timestamp 1586364061
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_270
timestamp 1586364061
transform 1 0 25944 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal3 s 27520 2320 28000 2440 6 address[0]
port 0 nsew default input
rlabel metal2 s 2778 0 2834 480 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 824 480 944 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 2456 480 2576 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 4088 480 4208 6 address[4]
port 4 nsew default input
rlabel metal2 s 3882 0 3938 480 6 address[5]
port 5 nsew default input
rlabel metal3 s 27520 6944 28000 7064 6 bottom_left_grid_pin_11_
port 6 nsew default input
rlabel metal2 s 2870 27520 2926 28000 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal3 s 0 10616 480 10736 6 bottom_left_grid_pin_15_
port 8 nsew default input
rlabel metal3 s 0 5720 480 5840 6 bottom_left_grid_pin_1_
port 9 nsew default input
rlabel metal3 s 0 7352 480 7472 6 bottom_left_grid_pin_3_
port 10 nsew default input
rlabel metal2 s 938 27520 994 28000 6 bottom_left_grid_pin_5_
port 11 nsew default input
rlabel metal3 s 0 8984 480 9104 6 bottom_left_grid_pin_7_
port 12 nsew default input
rlabel metal2 s 4986 0 5042 480 6 bottom_left_grid_pin_9_
port 13 nsew default input
rlabel metal3 s 0 12248 480 12368 6 bottom_right_grid_pin_11_
port 14 nsew default input
rlabel metal3 s 27520 11568 28000 11688 6 chanx_right_in[0]
port 15 nsew default input
rlabel metal3 s 27520 16328 28000 16448 6 chanx_right_in[1]
port 16 nsew default input
rlabel metal3 s 27520 20952 28000 21072 6 chanx_right_in[2]
port 17 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_right_in[3]
port 18 nsew default input
rlabel metal2 s 6090 0 6146 480 6 chanx_right_in[4]
port 19 nsew default input
rlabel metal2 s 4894 27520 4950 28000 6 chanx_right_in[5]
port 20 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chanx_right_in[6]
port 21 nsew default input
rlabel metal3 s 0 15648 480 15768 6 chanx_right_in[7]
port 22 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chanx_right_in[8]
port 23 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chanx_right_out[0]
port 24 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 chanx_right_out[1]
port 25 nsew default tristate
rlabel metal2 s 11702 0 11758 480 6 chanx_right_out[2]
port 26 nsew default tristate
rlabel metal2 s 6918 27520 6974 28000 6 chanx_right_out[3]
port 27 nsew default tristate
rlabel metal2 s 12806 0 12862 480 6 chanx_right_out[4]
port 28 nsew default tristate
rlabel metal2 s 8850 27520 8906 28000 6 chanx_right_out[5]
port 29 nsew default tristate
rlabel metal2 s 10874 27520 10930 28000 6 chanx_right_out[6]
port 30 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 chanx_right_out[7]
port 31 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 chanx_right_out[8]
port 32 nsew default tristate
rlabel metal2 s 12898 27520 12954 28000 6 chany_bottom_in[0]
port 33 nsew default input
rlabel metal3 s 0 17280 480 17400 6 chany_bottom_in[1]
port 34 nsew default input
rlabel metal3 s 0 18912 480 19032 6 chany_bottom_in[2]
port 35 nsew default input
rlabel metal3 s 27520 25576 28000 25696 6 chany_bottom_in[3]
port 36 nsew default input
rlabel metal2 s 16210 0 16266 480 6 chany_bottom_in[4]
port 37 nsew default input
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_in[5]
port 38 nsew default input
rlabel metal2 s 14922 27520 14978 28000 6 chany_bottom_in[6]
port 39 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chany_bottom_in[7]
port 40 nsew default input
rlabel metal2 s 18418 0 18474 480 6 chany_bottom_in[8]
port 41 nsew default input
rlabel metal2 s 19522 0 19578 480 6 chany_bottom_out[0]
port 42 nsew default tristate
rlabel metal2 s 16854 27520 16910 28000 6 chany_bottom_out[1]
port 43 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_out[2]
port 44 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chany_bottom_out[3]
port 45 nsew default tristate
rlabel metal2 s 21822 0 21878 480 6 chany_bottom_out[4]
port 46 nsew default tristate
rlabel metal2 s 22926 0 22982 480 6 chany_bottom_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 23808 480 23928 6 chany_bottom_out[6]
port 48 nsew default tristate
rlabel metal3 s 0 25440 480 25560 6 chany_bottom_out[7]
port 49 nsew default tristate
rlabel metal2 s 18878 27520 18934 28000 6 chany_bottom_out[8]
port 50 nsew default tristate
rlabel metal2 s 1674 0 1730 480 6 data_in
port 51 nsew default input
rlabel metal2 s 570 0 626 480 6 enable
port 52 nsew default input
rlabel metal2 s 24030 0 24086 480 6 right_bottom_grid_pin_12_
port 53 nsew default input
rlabel metal2 s 27342 0 27398 480 6 right_top_grid_pin_11_
port 54 nsew default input
rlabel metal2 s 24858 27520 24914 28000 6 right_top_grid_pin_13_
port 55 nsew default input
rlabel metal2 s 26882 27520 26938 28000 6 right_top_grid_pin_15_
port 56 nsew default input
rlabel metal2 s 25134 0 25190 480 6 right_top_grid_pin_1_
port 57 nsew default input
rlabel metal2 s 20902 27520 20958 28000 6 right_top_grid_pin_3_
port 58 nsew default input
rlabel metal3 s 0 27072 480 27192 6 right_top_grid_pin_5_
port 59 nsew default input
rlabel metal2 s 26238 0 26294 480 6 right_top_grid_pin_7_
port 60 nsew default input
rlabel metal2 s 22834 27520 22890 28000 6 right_top_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
