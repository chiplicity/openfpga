magic
tech sky130A
magscale 1 2
timestamp 1608763783
<< checkpaint >>
rect -1260 -1260 21260 18260
<< locali >>
rect 6653 12699 6687 12937
rect 11621 12155 11655 12325
rect 7757 11679 7791 11781
rect 13185 11543 13219 11849
rect 15669 11611 15703 11849
rect 9965 10455 9999 10557
rect 11989 10047 12023 10217
rect 4997 9435 5031 9673
rect 2881 8823 2915 8993
rect 9505 8891 9539 9061
rect 12909 7939 12943 8041
rect 3709 7191 3743 7293
rect 13737 7259 13771 7361
rect 6653 5015 6687 5321
rect 2421 4539 2455 4641
rect 6561 4063 6595 4165
rect 12173 3927 12207 4097
rect 12817 3451 12851 3621
rect 9781 2295 9815 2465
rect 13461 2295 13495 2601
<< viali >>
rect 1593 14433 1627 14467
rect 1777 14365 1811 14399
rect 6285 14025 6319 14059
rect 18245 14025 18279 14059
rect 16681 13957 16715 13991
rect 1777 13889 1811 13923
rect 2605 13889 2639 13923
rect 10057 13889 10091 13923
rect 10609 13889 10643 13923
rect 17325 13889 17359 13923
rect 1593 13821 1627 13855
rect 2329 13821 2363 13855
rect 6101 13821 6135 13855
rect 9873 13821 9907 13855
rect 10425 13821 10459 13855
rect 16497 13821 16531 13855
rect 17049 13821 17083 13855
rect 18061 13821 18095 13855
rect 9413 13685 9447 13719
rect 9781 13685 9815 13719
rect 11437 13413 11471 13447
rect 1869 13345 1903 13379
rect 2605 13345 2639 13379
rect 10333 13345 10367 13379
rect 10425 13345 10459 13379
rect 11345 13345 11379 13379
rect 16957 13345 16991 13379
rect 17693 13345 17727 13379
rect 2053 13277 2087 13311
rect 10517 13277 10551 13311
rect 11529 13277 11563 13311
rect 17233 13277 17267 13311
rect 17969 13277 18003 13311
rect 2789 13209 2823 13243
rect 9965 13141 9999 13175
rect 10977 13141 11011 13175
rect 6653 12937 6687 12971
rect 11345 12937 11379 12971
rect 3065 12869 3099 12903
rect 1777 12801 1811 12835
rect 3617 12801 3651 12835
rect 1593 12733 1627 12767
rect 3525 12733 3559 12767
rect 7849 12869 7883 12903
rect 16681 12869 16715 12903
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 8401 12801 8435 12835
rect 9965 12801 9999 12835
rect 10977 12801 11011 12835
rect 11989 12801 12023 12835
rect 17233 12801 17267 12835
rect 11805 12733 11839 12767
rect 18061 12733 18095 12767
rect 3433 12665 3467 12699
rect 6653 12665 6687 12699
rect 6837 12597 6871 12631
rect 7205 12597 7239 12631
rect 8217 12597 8251 12631
rect 8309 12597 8343 12631
rect 9321 12597 9355 12631
rect 9689 12597 9723 12631
rect 9781 12597 9815 12631
rect 10333 12597 10367 12631
rect 10701 12597 10735 12631
rect 10793 12597 10827 12631
rect 11713 12597 11747 12631
rect 17049 12597 17083 12631
rect 17141 12597 17175 12631
rect 18245 12597 18279 12631
rect 1869 12393 1903 12427
rect 3249 12393 3283 12427
rect 7573 12393 7607 12427
rect 8953 12393 8987 12427
rect 9045 12393 9079 12427
rect 9689 12393 9723 12427
rect 10149 12393 10183 12427
rect 10701 12393 10735 12427
rect 11713 12393 11747 12427
rect 17325 12393 17359 12427
rect 17785 12393 17819 12427
rect 7941 12325 7975 12359
rect 11621 12325 11655 12359
rect 12081 12325 12115 12359
rect 2237 12257 2271 12291
rect 6184 12257 6218 12291
rect 10057 12257 10091 12291
rect 11069 12257 11103 12291
rect 11161 12257 11195 12291
rect 2329 12189 2363 12223
rect 2513 12189 2547 12223
rect 3341 12189 3375 12223
rect 3433 12189 3467 12223
rect 5917 12189 5951 12223
rect 8033 12189 8067 12223
rect 8125 12189 8159 12223
rect 9229 12189 9263 12223
rect 10333 12189 10367 12223
rect 11253 12189 11287 12223
rect 12173 12257 12207 12291
rect 13921 12257 13955 12291
rect 15577 12257 15611 12291
rect 16681 12257 16715 12291
rect 16773 12257 16807 12291
rect 17693 12257 17727 12291
rect 12265 12189 12299 12223
rect 14289 12189 14323 12223
rect 15761 12189 15795 12223
rect 16957 12189 16991 12223
rect 17877 12189 17911 12223
rect 2881 12121 2915 12155
rect 7297 12121 7331 12155
rect 11621 12121 11655 12155
rect 8585 12053 8619 12087
rect 16313 12053 16347 12087
rect 2145 11849 2179 11883
rect 3157 11849 3191 11883
rect 4629 11849 4663 11883
rect 8861 11849 8895 11883
rect 10701 11849 10735 11883
rect 13185 11849 13219 11883
rect 6837 11781 6871 11815
rect 7757 11781 7791 11815
rect 7849 11781 7883 11815
rect 2697 11713 2731 11747
rect 3709 11713 3743 11747
rect 5273 11713 5307 11747
rect 6193 11713 6227 11747
rect 6377 11713 6411 11747
rect 7481 11713 7515 11747
rect 8309 11713 8343 11747
rect 8493 11713 8527 11747
rect 9413 11713 9447 11747
rect 11161 11713 11195 11747
rect 11345 11713 11379 11747
rect 2513 11645 2547 11679
rect 5089 11645 5123 11679
rect 6101 11645 6135 11679
rect 7757 11645 7791 11679
rect 3525 11577 3559 11611
rect 7205 11577 7239 11611
rect 7297 11577 7331 11611
rect 9321 11577 9355 11611
rect 15669 11849 15703 11883
rect 13921 11713 13955 11747
rect 15117 11645 15151 11679
rect 15853 11713 15887 11747
rect 17509 11713 17543 11747
rect 18061 11645 18095 11679
rect 13737 11577 13771 11611
rect 15393 11577 15427 11611
rect 15669 11577 15703 11611
rect 16120 11577 16154 11611
rect 2605 11509 2639 11543
rect 3617 11509 3651 11543
rect 4997 11509 5031 11543
rect 5733 11509 5767 11543
rect 8217 11509 8251 11543
rect 9229 11509 9263 11543
rect 11069 11509 11103 11543
rect 13185 11509 13219 11543
rect 13369 11509 13403 11543
rect 13829 11509 13863 11543
rect 17233 11509 17267 11543
rect 18245 11509 18279 11543
rect 3525 11305 3559 11339
rect 7481 11305 7515 11339
rect 11069 11305 11103 11339
rect 11345 11305 11379 11339
rect 17233 11305 17267 11339
rect 6000 11237 6034 11271
rect 9956 11237 9990 11271
rect 12725 11237 12759 11271
rect 17601 11237 17635 11271
rect 2145 11169 2179 11203
rect 2412 11169 2446 11203
rect 4077 11169 4111 11203
rect 4344 11169 4378 11203
rect 5733 11169 5767 11203
rect 8208 11169 8242 11203
rect 12633 11169 12667 11203
rect 13544 11169 13578 11203
rect 15568 11169 15602 11203
rect 1685 11101 1719 11135
rect 7941 11101 7975 11135
rect 9689 11101 9723 11135
rect 12909 11101 12943 11135
rect 13277 11101 13311 11135
rect 15301 11101 15335 11135
rect 17693 11101 17727 11135
rect 17877 11101 17911 11135
rect 5457 11033 5491 11067
rect 7113 11033 7147 11067
rect 9321 11033 9355 11067
rect 14657 11033 14691 11067
rect 16681 11033 16715 11067
rect 12265 10965 12299 10999
rect 2145 10761 2179 10795
rect 3433 10761 3467 10795
rect 5457 10761 5491 10795
rect 6837 10761 6871 10795
rect 9873 10761 9907 10795
rect 11161 10761 11195 10795
rect 16957 10761 16991 10795
rect 7849 10693 7883 10727
rect 2789 10625 2823 10659
rect 4077 10625 4111 10659
rect 4997 10625 5031 10659
rect 6009 10625 6043 10659
rect 7389 10625 7423 10659
rect 8493 10625 8527 10659
rect 10609 10625 10643 10659
rect 10701 10625 10735 10659
rect 11621 10625 11655 10659
rect 11713 10625 11747 10659
rect 17417 10625 17451 10659
rect 17601 10625 17635 10659
rect 1593 10557 1627 10591
rect 2513 10557 2547 10591
rect 5917 10557 5951 10591
rect 7205 10557 7239 10591
rect 8033 10557 8067 10591
rect 9965 10557 9999 10591
rect 10517 10557 10551 10591
rect 12449 10557 12483 10591
rect 12716 10557 12750 10591
rect 14197 10557 14231 10591
rect 14749 10557 14783 10591
rect 16405 10557 16439 10591
rect 18061 10557 18095 10591
rect 3801 10489 3835 10523
rect 4905 10489 4939 10523
rect 5825 10489 5859 10523
rect 8760 10489 8794 10523
rect 15016 10489 15050 10523
rect 1777 10421 1811 10455
rect 2605 10421 2639 10455
rect 3893 10421 3927 10455
rect 4445 10421 4479 10455
rect 4813 10421 4847 10455
rect 7297 10421 7331 10455
rect 9965 10421 9999 10455
rect 10149 10421 10183 10455
rect 11529 10421 11563 10455
rect 13829 10421 13863 10455
rect 14381 10421 14415 10455
rect 16129 10421 16163 10455
rect 16589 10421 16623 10455
rect 17325 10421 17359 10455
rect 18245 10421 18279 10455
rect 2789 10217 2823 10251
rect 4445 10217 4479 10251
rect 10149 10217 10183 10251
rect 11989 10217 12023 10251
rect 13553 10217 13587 10251
rect 13921 10217 13955 10251
rect 14289 10217 14323 10251
rect 15301 10217 15335 10251
rect 16313 10217 16347 10251
rect 17785 10217 17819 10251
rect 1676 10149 1710 10183
rect 6644 10149 6678 10183
rect 8493 10149 8527 10183
rect 10057 10149 10091 10183
rect 11529 10149 11563 10183
rect 11621 10149 11655 10183
rect 1409 10081 1443 10115
rect 3065 10081 3099 10115
rect 4813 10081 4847 10115
rect 5641 10081 5675 10115
rect 6377 10081 6411 10115
rect 8401 10081 8435 10115
rect 10977 10081 11011 10115
rect 16681 10149 16715 10183
rect 12440 10081 12474 10115
rect 15117 10081 15151 10115
rect 15669 10081 15703 10115
rect 15761 10081 15795 10115
rect 16773 10081 16807 10115
rect 17693 10081 17727 10115
rect 4905 10013 4939 10047
rect 4997 10013 5031 10047
rect 8585 10013 8619 10047
rect 10241 10013 10275 10047
rect 11805 10013 11839 10047
rect 11989 10013 12023 10047
rect 12173 10013 12207 10047
rect 14381 10013 14415 10047
rect 14473 10013 14507 10047
rect 15853 10013 15887 10047
rect 16865 10013 16899 10047
rect 17877 10013 17911 10047
rect 5457 9945 5491 9979
rect 8033 9945 8067 9979
rect 10793 9945 10827 9979
rect 17325 9945 17359 9979
rect 3249 9877 3283 9911
rect 7757 9877 7791 9911
rect 9689 9877 9723 9911
rect 11161 9877 11195 9911
rect 14933 9877 14967 9911
rect 4997 9673 5031 9707
rect 6469 9673 6503 9707
rect 8861 9673 8895 9707
rect 4721 9537 4755 9571
rect 1409 9469 1443 9503
rect 1961 9469 1995 9503
rect 2228 9469 2262 9503
rect 3801 9469 3835 9503
rect 11069 9605 11103 9639
rect 11345 9605 11379 9639
rect 12633 9605 12667 9639
rect 14013 9605 14047 9639
rect 7481 9537 7515 9571
rect 11989 9537 12023 9571
rect 13553 9537 13587 9571
rect 14565 9537 14599 9571
rect 15577 9537 15611 9571
rect 5089 9469 5123 9503
rect 7205 9469 7239 9503
rect 9137 9469 9171 9503
rect 11253 9469 11287 9503
rect 11713 9469 11747 9503
rect 12449 9469 12483 9503
rect 15025 9469 15059 9503
rect 15844 9469 15878 9503
rect 17233 9469 17267 9503
rect 18061 9469 18095 9503
rect 4997 9401 5031 9435
rect 5356 9401 5390 9435
rect 7748 9401 7782 9435
rect 9382 9401 9416 9435
rect 14473 9401 14507 9435
rect 17509 9401 17543 9435
rect 1593 9333 1627 9367
rect 3341 9333 3375 9367
rect 3617 9333 3651 9367
rect 4077 9333 4111 9367
rect 4445 9333 4479 9367
rect 4537 9333 4571 9367
rect 7021 9333 7055 9367
rect 10517 9333 10551 9367
rect 11805 9333 11839 9367
rect 13001 9333 13035 9367
rect 13369 9333 13403 9367
rect 13461 9333 13495 9367
rect 14381 9333 14415 9367
rect 15209 9333 15243 9367
rect 16957 9333 16991 9367
rect 18245 9333 18279 9367
rect 5457 9129 5491 9163
rect 5733 9129 5767 9163
rect 7941 9129 7975 9163
rect 9689 9129 9723 9163
rect 10149 9129 10183 9163
rect 11437 9129 11471 9163
rect 12449 9129 12483 9163
rect 14841 9129 14875 9163
rect 15761 9129 15795 9163
rect 15853 9129 15887 9163
rect 1676 9061 1710 9095
rect 8401 9061 8435 9095
rect 9505 9061 9539 9095
rect 10057 9061 10091 9095
rect 10977 9061 11011 9095
rect 12909 9061 12943 9095
rect 1409 8993 1443 9027
rect 2881 8993 2915 9027
rect 3065 8993 3099 9027
rect 4344 8993 4378 9027
rect 6285 8993 6319 9027
rect 6552 8993 6586 9027
rect 8309 8993 8343 9027
rect 4077 8925 4111 8959
rect 8585 8925 8619 8959
rect 10701 8993 10735 9027
rect 11805 8993 11839 9027
rect 12817 8993 12851 9027
rect 13728 8993 13762 9027
rect 16405 8993 16439 9027
rect 16672 8993 16706 9027
rect 18061 8993 18095 9027
rect 10241 8925 10275 8959
rect 11897 8925 11931 8959
rect 12081 8925 12115 8959
rect 13093 8925 13127 8959
rect 13461 8925 13495 8959
rect 15945 8925 15979 8959
rect 3249 8857 3283 8891
rect 9505 8857 9539 8891
rect 2789 8789 2823 8823
rect 2881 8789 2915 8823
rect 7665 8789 7699 8823
rect 15393 8789 15427 8823
rect 17785 8789 17819 8823
rect 18245 8789 18279 8823
rect 3985 8585 4019 8619
rect 9229 8585 9263 8619
rect 1869 8517 1903 8551
rect 3709 8517 3743 8551
rect 4997 8517 5031 8551
rect 11437 8517 11471 8551
rect 11529 8517 11563 8551
rect 13553 8517 13587 8551
rect 18245 8517 18279 8551
rect 4537 8449 4571 8483
rect 5549 8449 5583 8483
rect 7573 8449 7607 8483
rect 9781 8449 9815 8483
rect 12081 8449 12115 8483
rect 13093 8449 13127 8483
rect 14105 8449 14139 8483
rect 14565 8449 14599 8483
rect 17233 8449 17267 8483
rect 1685 8381 1719 8415
rect 2329 8381 2363 8415
rect 6009 8381 6043 8415
rect 9597 8381 9631 8415
rect 10057 8381 10091 8415
rect 10324 8381 10358 8415
rect 11897 8381 11931 8415
rect 11989 8381 12023 8415
rect 12817 8381 12851 8415
rect 13921 8381 13955 8415
rect 15025 8381 15059 8415
rect 17049 8381 17083 8415
rect 17141 8381 17175 8415
rect 18061 8381 18095 8415
rect 2596 8313 2630 8347
rect 5457 8313 5491 8347
rect 7113 8313 7147 8347
rect 7840 8313 7874 8347
rect 9689 8313 9723 8347
rect 12909 8313 12943 8347
rect 14013 8313 14047 8347
rect 15292 8313 15326 8347
rect 4353 8245 4387 8279
rect 4445 8245 4479 8279
rect 5365 8245 5399 8279
rect 6193 8245 6227 8279
rect 8953 8245 8987 8279
rect 12449 8245 12483 8279
rect 16405 8245 16439 8279
rect 16681 8245 16715 8279
rect 2329 8041 2363 8075
rect 2973 8041 3007 8075
rect 3433 8041 3467 8075
rect 4077 8041 4111 8075
rect 8401 8041 8435 8075
rect 8769 8041 8803 8075
rect 10333 8041 10367 8075
rect 12725 8041 12759 8075
rect 12909 8041 12943 8075
rect 14381 8041 14415 8075
rect 17417 8041 17451 8075
rect 5356 7973 5390 8007
rect 8861 7973 8895 8007
rect 1409 7905 1443 7939
rect 3341 7905 3375 7939
rect 4445 7905 4479 7939
rect 5089 7905 5123 7939
rect 7012 7905 7046 7939
rect 9689 7905 9723 7939
rect 10701 7905 10735 7939
rect 11612 7905 11646 7939
rect 12909 7905 12943 7939
rect 13257 7905 13291 7939
rect 14657 7905 14691 7939
rect 15568 7905 15602 7939
rect 17325 7905 17359 7939
rect 17969 7905 18003 7939
rect 2421 7837 2455 7871
rect 2605 7837 2639 7871
rect 3525 7837 3559 7871
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 6745 7837 6779 7871
rect 8953 7837 8987 7871
rect 9873 7837 9907 7871
rect 10793 7837 10827 7871
rect 10977 7837 11011 7871
rect 11345 7837 11379 7871
rect 13008 7837 13042 7871
rect 15301 7837 15335 7871
rect 17509 7837 17543 7871
rect 1593 7769 1627 7803
rect 6469 7769 6503 7803
rect 1961 7701 1995 7735
rect 8125 7701 8159 7735
rect 14841 7701 14875 7735
rect 16681 7701 16715 7735
rect 16957 7701 16991 7735
rect 18153 7701 18187 7735
rect 2881 7497 2915 7531
rect 5917 7497 5951 7531
rect 10241 7497 10275 7531
rect 12633 7497 12667 7531
rect 12909 7497 12943 7531
rect 15301 7497 15335 7531
rect 1869 7429 1903 7463
rect 11345 7429 11379 7463
rect 1409 7361 1443 7395
rect 2513 7361 2547 7395
rect 3433 7361 3467 7395
rect 7389 7361 7423 7395
rect 11989 7361 12023 7395
rect 13461 7361 13495 7395
rect 13737 7361 13771 7395
rect 16589 7361 16623 7395
rect 3709 7293 3743 7327
rect 3893 7293 3927 7327
rect 4537 7293 4571 7327
rect 4804 7293 4838 7327
rect 6193 7293 6227 7327
rect 7849 7293 7883 7327
rect 8953 7293 8987 7327
rect 12817 7293 12851 7327
rect 13921 7293 13955 7327
rect 16497 7293 16531 7327
rect 17049 7293 17083 7327
rect 18061 7293 18095 7327
rect 7205 7225 7239 7259
rect 8125 7225 8159 7259
rect 11713 7225 11747 7259
rect 13277 7225 13311 7259
rect 13737 7225 13771 7259
rect 14188 7225 14222 7259
rect 17325 7225 17359 7259
rect 2237 7157 2271 7191
rect 2329 7157 2363 7191
rect 3249 7157 3283 7191
rect 3341 7157 3375 7191
rect 3709 7157 3743 7191
rect 4077 7157 4111 7191
rect 6377 7157 6411 7191
rect 6837 7157 6871 7191
rect 7297 7157 7331 7191
rect 10793 7157 10827 7191
rect 11805 7157 11839 7191
rect 13369 7157 13403 7191
rect 15577 7157 15611 7191
rect 16037 7157 16071 7191
rect 16405 7157 16439 7191
rect 18245 7157 18279 7191
rect 6285 6953 6319 6987
rect 7573 6953 7607 6987
rect 8953 6953 8987 6987
rect 10517 6953 10551 6987
rect 10885 6953 10919 6987
rect 13921 6953 13955 6987
rect 14289 6953 14323 6987
rect 14381 6953 14415 6987
rect 7941 6885 7975 6919
rect 1676 6817 1710 6851
rect 3065 6817 3099 6851
rect 3801 6817 3835 6851
rect 4077 6817 4111 6851
rect 4813 6817 4847 6851
rect 5172 6817 5206 6851
rect 6929 6817 6963 6851
rect 9689 6817 9723 6851
rect 10977 6817 11011 6851
rect 11785 6817 11819 6851
rect 13185 6817 13219 6851
rect 15752 6817 15786 6851
rect 17509 6817 17543 6851
rect 1409 6749 1443 6783
rect 4905 6749 4939 6783
rect 7021 6749 7055 6783
rect 7113 6749 7147 6783
rect 8033 6749 8067 6783
rect 8125 6749 8159 6783
rect 9045 6749 9079 6783
rect 9137 6749 9171 6783
rect 9873 6749 9907 6783
rect 11069 6749 11103 6783
rect 11529 6749 11563 6783
rect 13369 6749 13403 6783
rect 14473 6749 14507 6783
rect 15485 6749 15519 6783
rect 17601 6749 17635 6783
rect 17693 6749 17727 6783
rect 18153 6749 18187 6783
rect 2789 6681 2823 6715
rect 3249 6681 3283 6715
rect 8585 6681 8619 6715
rect 12909 6681 12943 6715
rect 3617 6613 3651 6647
rect 4261 6613 4295 6647
rect 4629 6613 4663 6647
rect 6561 6613 6595 6647
rect 16865 6613 16899 6647
rect 17141 6613 17175 6647
rect 1777 6409 1811 6443
rect 8217 6409 8251 6443
rect 14013 6409 14047 6443
rect 10057 6341 10091 6375
rect 13001 6341 13035 6375
rect 2421 6273 2455 6307
rect 2789 6273 2823 6307
rect 12449 6273 12483 6307
rect 13645 6273 13679 6307
rect 14565 6273 14599 6307
rect 15577 6273 15611 6307
rect 2145 6205 2179 6239
rect 3056 6205 3090 6239
rect 4445 6205 4479 6239
rect 6101 6205 6135 6239
rect 6837 6205 6871 6239
rect 8677 6205 8711 6239
rect 10149 6205 10183 6239
rect 10405 6205 10439 6239
rect 12265 6205 12299 6239
rect 16313 6205 16347 6239
rect 18061 6205 18095 6239
rect 4690 6137 4724 6171
rect 7104 6137 7138 6171
rect 8944 6137 8978 6171
rect 13369 6137 13403 6171
rect 15485 6137 15519 6171
rect 16580 6137 16614 6171
rect 2237 6069 2271 6103
rect 4169 6069 4203 6103
rect 5825 6069 5859 6103
rect 6285 6069 6319 6103
rect 11529 6069 11563 6103
rect 12081 6069 12115 6103
rect 13461 6069 13495 6103
rect 14381 6069 14415 6103
rect 14473 6069 14507 6103
rect 15025 6069 15059 6103
rect 15393 6069 15427 6103
rect 17693 6069 17727 6103
rect 18245 6069 18279 6103
rect 1869 5865 1903 5899
rect 2881 5865 2915 5899
rect 4077 5865 4111 5899
rect 4445 5865 4479 5899
rect 5457 5865 5491 5899
rect 6929 5865 6963 5899
rect 7941 5865 7975 5899
rect 9873 5865 9907 5899
rect 10333 5865 10367 5899
rect 14197 5865 14231 5899
rect 15853 5865 15887 5899
rect 17325 5865 17359 5899
rect 3341 5797 3375 5831
rect 8309 5797 8343 5831
rect 10057 5797 10091 5831
rect 13062 5797 13096 5831
rect 15761 5797 15795 5831
rect 2237 5729 2271 5763
rect 3249 5729 3283 5763
rect 4537 5729 4571 5763
rect 5549 5729 5583 5763
rect 6101 5729 6135 5763
rect 7297 5729 7331 5763
rect 9137 5729 9171 5763
rect 9689 5729 9723 5763
rect 10701 5729 10735 5763
rect 10793 5729 10827 5763
rect 11161 5729 11195 5763
rect 11428 5729 11462 5763
rect 12817 5729 12851 5763
rect 14473 5729 14507 5763
rect 16405 5729 16439 5763
rect 17969 5729 18003 5763
rect 2329 5661 2363 5695
rect 2513 5661 2547 5695
rect 3433 5661 3467 5695
rect 4629 5661 4663 5695
rect 5733 5661 5767 5695
rect 6285 5661 6319 5695
rect 7389 5661 7423 5695
rect 7481 5661 7515 5695
rect 8401 5661 8435 5695
rect 8585 5661 8619 5695
rect 9229 5661 9263 5695
rect 9321 5661 9355 5695
rect 10977 5661 11011 5695
rect 14657 5661 14691 5695
rect 16037 5661 16071 5695
rect 17417 5661 17451 5695
rect 17601 5661 17635 5695
rect 12541 5593 12575 5627
rect 5089 5525 5123 5559
rect 8769 5525 8803 5559
rect 15393 5525 15427 5559
rect 16589 5525 16623 5559
rect 16957 5525 16991 5559
rect 18153 5525 18187 5559
rect 3709 5321 3743 5355
rect 6653 5321 6687 5355
rect 6837 5321 6871 5355
rect 7849 5321 7883 5355
rect 11345 5321 11379 5355
rect 13553 5321 13587 5355
rect 4629 5185 4663 5219
rect 1685 5117 1719 5151
rect 2329 5117 2363 5151
rect 3985 5117 4019 5151
rect 4896 5117 4930 5151
rect 2574 5049 2608 5083
rect 10425 5253 10459 5287
rect 7481 5185 7515 5219
rect 8401 5185 8435 5219
rect 11989 5185 12023 5219
rect 12909 5185 12943 5219
rect 13093 5185 13127 5219
rect 14197 5185 14231 5219
rect 15117 5185 15151 5219
rect 17233 5185 17267 5219
rect 17325 5185 17359 5219
rect 8217 5117 8251 5151
rect 9045 5117 9079 5151
rect 13921 5117 13955 5151
rect 15384 5117 15418 5151
rect 17141 5117 17175 5151
rect 18061 5117 18095 5151
rect 9312 5049 9346 5083
rect 11713 5049 11747 5083
rect 12817 5049 12851 5083
rect 1869 4981 1903 5015
rect 4169 4981 4203 5015
rect 6009 4981 6043 5015
rect 6285 4981 6319 5015
rect 6653 4981 6687 5015
rect 7205 4981 7239 5015
rect 7297 4981 7331 5015
rect 8309 4981 8343 5015
rect 10885 4981 10919 5015
rect 11805 4981 11839 5015
rect 12449 4981 12483 5015
rect 14013 4981 14047 5015
rect 14565 4981 14599 5015
rect 16497 4981 16531 5015
rect 16773 4981 16807 5015
rect 18245 4981 18279 5015
rect 2605 4777 2639 4811
rect 4077 4777 4111 4811
rect 4445 4777 4479 4811
rect 5549 4777 5583 4811
rect 8493 4777 8527 4811
rect 12725 4777 12759 4811
rect 14933 4777 14967 4811
rect 15301 4777 15335 4811
rect 15761 4777 15795 4811
rect 17509 4777 17543 4811
rect 17601 4777 17635 4811
rect 9045 4709 9079 4743
rect 10048 4709 10082 4743
rect 15669 4709 15703 4743
rect 1501 4641 1535 4675
rect 2053 4641 2087 4675
rect 2421 4641 2455 4675
rect 2973 4641 3007 4675
rect 4537 4641 4571 4675
rect 5457 4641 5491 4675
rect 6469 4641 6503 4675
rect 7113 4641 7147 4675
rect 7380 4641 7414 4675
rect 8769 4641 8803 4675
rect 11621 4641 11655 4675
rect 13820 4641 13854 4675
rect 16313 4641 16347 4675
rect 3065 4573 3099 4607
rect 3249 4573 3283 4607
rect 4629 4573 4663 4607
rect 5733 4573 5767 4607
rect 6561 4573 6595 4607
rect 6745 4573 6779 4607
rect 9781 4573 9815 4607
rect 11897 4573 11931 4607
rect 12817 4573 12851 4607
rect 13001 4573 13035 4607
rect 13553 4573 13587 4607
rect 15945 4573 15979 4607
rect 16497 4573 16531 4607
rect 17693 4573 17727 4607
rect 2237 4505 2271 4539
rect 2421 4505 2455 4539
rect 5089 4505 5123 4539
rect 12357 4505 12391 4539
rect 1685 4437 1719 4471
rect 6101 4437 6135 4471
rect 11161 4437 11195 4471
rect 17141 4437 17175 4471
rect 8217 4233 8251 4267
rect 12541 4233 12575 4267
rect 6561 4165 6595 4199
rect 10333 4165 10367 4199
rect 14657 4165 14691 4199
rect 2145 4097 2179 4131
rect 3065 4097 3099 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 8493 4097 8527 4131
rect 10977 4097 11011 4131
rect 11897 4097 11931 4131
rect 12173 4097 12207 4131
rect 13001 4097 13035 4131
rect 13185 4097 13219 4131
rect 14289 4097 14323 4131
rect 15209 4097 15243 4131
rect 17509 4097 17543 4131
rect 1869 4029 1903 4063
rect 2881 4029 2915 4063
rect 3525 4029 3559 4063
rect 3792 4029 3826 4063
rect 6193 4029 6227 4063
rect 6561 4029 6595 4063
rect 6837 4029 6871 4063
rect 8749 4029 8783 4063
rect 11713 4029 11747 4063
rect 7082 3961 7116 3995
rect 10701 3961 10735 3995
rect 11805 3961 11839 3995
rect 12909 4029 12943 4063
rect 14013 4029 14047 4063
rect 14841 4029 14875 4063
rect 15476 4029 15510 4063
rect 18061 4029 18095 4063
rect 17417 3961 17451 3995
rect 1501 3893 1535 3927
rect 1961 3893 1995 3927
rect 2513 3893 2547 3927
rect 2973 3893 3007 3927
rect 4905 3893 4939 3927
rect 5181 3893 5215 3927
rect 5549 3893 5583 3927
rect 6377 3893 6411 3927
rect 9873 3893 9907 3927
rect 10793 3893 10827 3927
rect 11345 3893 11379 3927
rect 12173 3893 12207 3927
rect 13645 3893 13679 3927
rect 14105 3893 14139 3927
rect 16589 3893 16623 3927
rect 16957 3893 16991 3927
rect 17325 3893 17359 3927
rect 18245 3893 18279 3927
rect 2789 3689 2823 3723
rect 4629 3689 4663 3723
rect 6929 3689 6963 3723
rect 7297 3689 7331 3723
rect 7757 3689 7791 3723
rect 8677 3689 8711 3723
rect 8769 3689 8803 3723
rect 14289 3689 14323 3723
rect 16405 3689 16439 3723
rect 16497 3689 16531 3723
rect 17049 3689 17083 3723
rect 17417 3689 17451 3723
rect 18245 3689 18279 3723
rect 4721 3621 4755 3655
rect 5540 3621 5574 3655
rect 12817 3621 12851 3655
rect 13176 3621 13210 3655
rect 17509 3621 17543 3655
rect 1665 3553 1699 3587
rect 3249 3553 3283 3587
rect 7113 3553 7147 3587
rect 7665 3553 7699 3587
rect 9505 3553 9539 3587
rect 9689 3553 9723 3587
rect 10609 3553 10643 3587
rect 10701 3553 10735 3587
rect 11253 3553 11287 3587
rect 11509 3553 11543 3587
rect 1409 3485 1443 3519
rect 3433 3485 3467 3519
rect 4813 3485 4847 3519
rect 5273 3485 5307 3519
rect 7941 3485 7975 3519
rect 8953 3485 8987 3519
rect 10885 3485 10919 3519
rect 15301 3553 15335 3587
rect 18061 3553 18095 3587
rect 12909 3485 12943 3519
rect 15485 3485 15519 3519
rect 16589 3485 16623 3519
rect 17601 3485 17635 3519
rect 9873 3417 9907 3451
rect 10241 3417 10275 3451
rect 12633 3417 12667 3451
rect 12817 3417 12851 3451
rect 4261 3349 4295 3383
rect 6653 3349 6687 3383
rect 8309 3349 8343 3383
rect 9321 3349 9355 3383
rect 16037 3349 16071 3383
rect 8125 3145 8159 3179
rect 10609 3145 10643 3179
rect 12449 3145 12483 3179
rect 13737 3145 13771 3179
rect 2513 3009 2547 3043
rect 3341 3009 3375 3043
rect 3525 3009 3559 3043
rect 4537 3009 4571 3043
rect 5549 3009 5583 3043
rect 7665 3009 7699 3043
rect 8677 3009 8711 3043
rect 11437 3009 11471 3043
rect 13001 3009 13035 3043
rect 14381 3009 14415 3043
rect 15393 3009 15427 3043
rect 16313 3009 16347 3043
rect 17233 3009 17267 3043
rect 17325 3009 17359 3043
rect 4353 2941 4387 2975
rect 6009 2941 6043 2975
rect 8585 2941 8619 2975
rect 9229 2941 9263 2975
rect 11253 2941 11287 2975
rect 12909 2941 12943 2975
rect 14197 2941 14231 2975
rect 16129 2941 16163 2975
rect 16221 2941 16255 2975
rect 2237 2873 2271 2907
rect 3249 2873 3283 2907
rect 6285 2873 6319 2907
rect 7481 2873 7515 2907
rect 9496 2873 9530 2907
rect 12817 2873 12851 2907
rect 14105 2873 14139 2907
rect 15117 2873 15151 2907
rect 17141 2873 17175 2907
rect 1869 2805 1903 2839
rect 2329 2805 2363 2839
rect 2881 2805 2915 2839
rect 3893 2805 3927 2839
rect 4261 2805 4295 2839
rect 4997 2805 5031 2839
rect 5365 2805 5399 2839
rect 5457 2805 5491 2839
rect 7113 2805 7147 2839
rect 7573 2805 7607 2839
rect 8493 2805 8527 2839
rect 10885 2805 10919 2839
rect 11345 2805 11379 2839
rect 14749 2805 14783 2839
rect 15209 2805 15243 2839
rect 15761 2805 15795 2839
rect 16773 2805 16807 2839
rect 2973 2601 3007 2635
rect 3341 2601 3375 2635
rect 4537 2601 4571 2635
rect 4997 2601 5031 2635
rect 5825 2601 5859 2635
rect 7389 2601 7423 2635
rect 8677 2601 8711 2635
rect 9873 2601 9907 2635
rect 10333 2601 10367 2635
rect 11253 2601 11287 2635
rect 11345 2601 11379 2635
rect 13001 2601 13035 2635
rect 13461 2601 13495 2635
rect 13645 2601 13679 2635
rect 14013 2601 14047 2635
rect 15669 2601 15703 2635
rect 16681 2601 16715 2635
rect 17141 2601 17175 2635
rect 3433 2533 3467 2567
rect 4905 2533 4939 2567
rect 8217 2533 8251 2567
rect 9137 2533 9171 2567
rect 1409 2465 1443 2499
rect 1961 2465 1995 2499
rect 6193 2465 6227 2499
rect 7297 2465 7331 2499
rect 7941 2465 7975 2499
rect 9045 2465 9079 2499
rect 9781 2465 9815 2499
rect 10241 2465 10275 2499
rect 2145 2397 2179 2431
rect 3525 2397 3559 2431
rect 5181 2397 5215 2431
rect 6285 2397 6319 2431
rect 6377 2397 6411 2431
rect 7481 2397 7515 2431
rect 9321 2397 9355 2431
rect 10517 2397 10551 2431
rect 11437 2397 11471 2431
rect 13093 2397 13127 2431
rect 13277 2397 13311 2431
rect 12633 2329 12667 2363
rect 14933 2533 14967 2567
rect 16037 2533 16071 2567
rect 16129 2533 16163 2567
rect 17049 2533 17083 2567
rect 14657 2465 14691 2499
rect 14105 2397 14139 2431
rect 14197 2397 14231 2431
rect 16313 2397 16347 2431
rect 17233 2397 17267 2431
rect 1593 2261 1627 2295
rect 6929 2261 6963 2295
rect 9781 2261 9815 2295
rect 10885 2261 10919 2295
rect 13461 2261 13495 2295
<< metal1 >>
rect 4062 15240 4068 15292
rect 4120 15280 4126 15292
rect 10502 15280 10508 15292
rect 4120 15252 10508 15280
rect 4120 15240 4126 15252
rect 10502 15240 10508 15252
rect 10560 15240 10566 15292
rect 3970 15172 3976 15224
rect 4028 15212 4034 15224
rect 15010 15212 15016 15224
rect 4028 15184 15016 15212
rect 4028 15172 4034 15184
rect 15010 15172 15016 15184
rect 15068 15172 15074 15224
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 1578 14560 1584 14612
rect 1636 14560 1642 14612
rect 1596 14532 1624 14560
rect 16942 14532 16948 14544
rect 1596 14504 16948 14532
rect 16942 14492 16948 14504
rect 17000 14492 17006 14544
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 2958 14464 2964 14476
rect 1627 14436 2964 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 2958 14424 2964 14436
rect 3016 14464 3022 14476
rect 7742 14464 7748 14476
rect 3016 14436 7748 14464
rect 3016 14424 3022 14436
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 1762 14396 1768 14408
rect 1723 14368 1768 14396
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 5902 14016 5908 14068
rect 5960 14056 5966 14068
rect 6273 14059 6331 14065
rect 6273 14056 6285 14059
rect 5960 14028 6285 14056
rect 5960 14016 5966 14028
rect 6273 14025 6285 14028
rect 6319 14025 6331 14059
rect 6273 14019 6331 14025
rect 7576 14028 10732 14056
rect 1946 13948 1952 14000
rect 2004 13988 2010 14000
rect 7576 13988 7604 14028
rect 2004 13960 7604 13988
rect 2004 13948 2010 13960
rect 9766 13948 9772 14000
rect 9824 13988 9830 14000
rect 9824 13960 10640 13988
rect 9824 13948 9830 13960
rect 1670 13880 1676 13932
rect 1728 13920 1734 13932
rect 1765 13923 1823 13929
rect 1765 13920 1777 13923
rect 1728 13892 1777 13920
rect 1728 13880 1734 13892
rect 1765 13889 1777 13892
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2774 13920 2780 13932
rect 2639 13892 2780 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 10045 13923 10103 13929
rect 10045 13889 10057 13923
rect 10091 13920 10103 13923
rect 10226 13920 10232 13932
rect 10091 13892 10232 13920
rect 10091 13889 10103 13892
rect 10045 13883 10103 13889
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 10612 13929 10640 13960
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 2866 13852 2872 13864
rect 2363 13824 2872 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 6086 13852 6092 13864
rect 6047 13824 6092 13852
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 9861 13855 9919 13861
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 10413 13855 10471 13861
rect 9907 13824 10272 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 3234 13744 3240 13796
rect 3292 13784 3298 13796
rect 10244 13784 10272 13824
rect 10413 13821 10425 13855
rect 10459 13852 10471 13855
rect 10502 13852 10508 13864
rect 10459 13824 10508 13852
rect 10459 13821 10471 13824
rect 10413 13815 10471 13821
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 10704 13852 10732 14028
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 18233 14059 18291 14065
rect 18233 14056 18245 14059
rect 16448 14028 18245 14056
rect 16448 14016 16454 14028
rect 18233 14025 18245 14028
rect 18279 14025 18291 14059
rect 18233 14019 18291 14025
rect 13906 13948 13912 14000
rect 13964 13988 13970 14000
rect 16669 13991 16727 13997
rect 13964 13960 16620 13988
rect 13964 13948 13970 13960
rect 16485 13855 16543 13861
rect 16485 13852 16497 13855
rect 10704 13824 16497 13852
rect 16485 13821 16497 13824
rect 16531 13821 16543 13855
rect 16592 13852 16620 13960
rect 16669 13957 16681 13991
rect 16715 13988 16727 13991
rect 17586 13988 17592 14000
rect 16715 13960 17592 13988
rect 16715 13957 16727 13960
rect 16669 13951 16727 13957
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 17313 13923 17371 13929
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 17862 13920 17868 13932
rect 17359 13892 17868 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 17862 13880 17868 13892
rect 17920 13880 17926 13932
rect 17037 13855 17095 13861
rect 17037 13852 17049 13855
rect 16592 13824 17049 13852
rect 16485 13815 16543 13821
rect 17037 13821 17049 13824
rect 17083 13821 17095 13855
rect 17037 13815 17095 13821
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 11514 13784 11520 13796
rect 3292 13756 9904 13784
rect 10244 13756 11520 13784
rect 3292 13744 3298 13756
rect 9401 13719 9459 13725
rect 9401 13685 9413 13719
rect 9447 13716 9459 13719
rect 9490 13716 9496 13728
rect 9447 13688 9496 13716
rect 9447 13685 9459 13688
rect 9401 13679 9459 13685
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 9766 13716 9772 13728
rect 9727 13688 9772 13716
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 9876 13716 9904 13756
rect 11514 13744 11520 13756
rect 11572 13744 11578 13796
rect 16206 13716 16212 13728
rect 9876 13688 16212 13716
rect 16206 13676 16212 13688
rect 16264 13716 16270 13728
rect 18064 13716 18092 13815
rect 16264 13688 18092 13716
rect 16264 13676 16270 13688
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 1486 13472 1492 13524
rect 1544 13512 1550 13524
rect 15562 13512 15568 13524
rect 1544 13484 15568 13512
rect 1544 13472 1550 13484
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 2866 13444 2872 13456
rect 1872 13416 2872 13444
rect 1872 13385 1900 13416
rect 2866 13404 2872 13416
rect 2924 13404 2930 13456
rect 11425 13447 11483 13453
rect 11425 13413 11437 13447
rect 11471 13444 11483 13447
rect 12434 13444 12440 13456
rect 11471 13416 12440 13444
rect 11471 13413 11483 13416
rect 11425 13407 11483 13413
rect 12434 13404 12440 13416
rect 12492 13404 12498 13456
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13345 1915 13379
rect 1857 13339 1915 13345
rect 2593 13379 2651 13385
rect 2593 13345 2605 13379
rect 2639 13376 2651 13379
rect 2774 13376 2780 13388
rect 2639 13348 2780 13376
rect 2639 13345 2651 13348
rect 2593 13339 2651 13345
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 10318 13376 10324 13388
rect 10279 13348 10324 13376
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 11238 13376 11244 13388
rect 10459 13348 11244 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 11238 13336 11244 13348
rect 11296 13336 11302 13388
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 12618 13376 12624 13388
rect 11379 13348 12624 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 16942 13376 16948 13388
rect 16903 13348 16948 13376
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 17681 13379 17739 13385
rect 17681 13345 17693 13379
rect 17727 13345 17739 13379
rect 17681 13339 17739 13345
rect 2038 13308 2044 13320
rect 1999 13280 2044 13308
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 10502 13308 10508 13320
rect 10463 13280 10508 13308
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 10778 13268 10784 13320
rect 10836 13308 10842 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 10836 13280 11529 13308
rect 10836 13268 10842 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 17218 13308 17224 13320
rect 17179 13280 17224 13308
rect 11517 13271 11575 13277
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 2774 13200 2780 13252
rect 2832 13240 2838 13252
rect 2832 13212 2877 13240
rect 2832 13200 2838 13212
rect 7098 13200 7104 13252
rect 7156 13240 7162 13252
rect 10410 13240 10416 13252
rect 7156 13212 10416 13240
rect 7156 13200 7162 13212
rect 10410 13200 10416 13212
rect 10468 13200 10474 13252
rect 10594 13200 10600 13252
rect 10652 13240 10658 13252
rect 17696 13240 17724 13339
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18506 13308 18512 13320
rect 18003 13280 18512 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 10652 13212 17724 13240
rect 10652 13200 10658 13212
rect 3786 13132 3792 13184
rect 3844 13172 3850 13184
rect 8846 13172 8852 13184
rect 3844 13144 8852 13172
rect 3844 13132 3850 13144
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 9953 13175 10011 13181
rect 9953 13172 9965 13175
rect 8996 13144 9965 13172
rect 8996 13132 9002 13144
rect 9953 13141 9965 13144
rect 9999 13141 10011 13175
rect 9953 13135 10011 13141
rect 10965 13175 11023 13181
rect 10965 13141 10977 13175
rect 11011 13172 11023 13175
rect 11606 13172 11612 13184
rect 11011 13144 11612 13172
rect 11011 13141 11023 13144
rect 10965 13135 11023 13141
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 8386 12968 8392 12980
rect 6687 12940 8392 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 10318 12928 10324 12980
rect 10376 12968 10382 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 10376 12940 11345 12968
rect 10376 12928 10382 12940
rect 11333 12937 11345 12940
rect 11379 12937 11391 12971
rect 17770 12968 17776 12980
rect 11333 12931 11391 12937
rect 13648 12940 17776 12968
rect 3053 12903 3111 12909
rect 3053 12869 3065 12903
rect 3099 12900 3111 12903
rect 7837 12903 7895 12909
rect 3099 12872 7788 12900
rect 3099 12869 3111 12872
rect 3053 12863 3111 12869
rect 1762 12832 1768 12844
rect 1723 12804 1768 12832
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 3326 12792 3332 12844
rect 3384 12832 3390 12844
rect 3605 12835 3663 12841
rect 3605 12832 3617 12835
rect 3384 12804 3617 12832
rect 3384 12792 3390 12804
rect 3605 12801 3617 12804
rect 3651 12801 3663 12835
rect 3605 12795 3663 12801
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 7248 12804 7297 12832
rect 7248 12792 7254 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 7285 12795 7343 12801
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7760 12832 7788 12872
rect 7837 12869 7849 12903
rect 7883 12900 7895 12903
rect 8754 12900 8760 12912
rect 7883 12872 8760 12900
rect 7883 12869 7895 12872
rect 7837 12863 7895 12869
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 8846 12860 8852 12912
rect 8904 12900 8910 12912
rect 13262 12900 13268 12912
rect 8904 12872 13268 12900
rect 8904 12860 8910 12872
rect 13262 12860 13268 12872
rect 13320 12860 13326 12912
rect 7760 12804 8064 12832
rect 1486 12724 1492 12776
rect 1544 12764 1550 12776
rect 1581 12767 1639 12773
rect 1581 12764 1593 12767
rect 1544 12736 1593 12764
rect 1544 12724 1550 12736
rect 1581 12733 1593 12736
rect 1627 12733 1639 12767
rect 1581 12727 1639 12733
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12764 3571 12767
rect 7926 12764 7932 12776
rect 3559 12736 7932 12764
rect 3559 12733 3571 12736
rect 3513 12727 3571 12733
rect 7926 12724 7932 12736
rect 7984 12724 7990 12776
rect 8036 12764 8064 12804
rect 8110 12792 8116 12844
rect 8168 12832 8174 12844
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 8168 12804 8401 12832
rect 8168 12792 8174 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10594 12832 10600 12844
rect 9999 12804 10600 12832
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 10594 12792 10600 12804
rect 10652 12792 10658 12844
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10928 12804 10977 12832
rect 10928 12792 10934 12804
rect 10965 12801 10977 12804
rect 11011 12832 11023 12835
rect 11977 12835 12035 12841
rect 11977 12832 11989 12835
rect 11011 12804 11989 12832
rect 11011 12801 11023 12804
rect 10965 12795 11023 12801
rect 11977 12801 11989 12804
rect 12023 12832 12035 12835
rect 12250 12832 12256 12844
rect 12023 12804 12256 12832
rect 12023 12801 12035 12804
rect 11977 12795 12035 12801
rect 12250 12792 12256 12804
rect 12308 12792 12314 12844
rect 8478 12764 8484 12776
rect 8036 12736 8484 12764
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 11422 12724 11428 12776
rect 11480 12764 11486 12776
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11480 12736 11805 12764
rect 11480 12724 11486 12736
rect 11793 12733 11805 12736
rect 11839 12764 11851 12767
rect 13648 12764 13676 12940
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 14918 12860 14924 12912
rect 14976 12900 14982 12912
rect 16669 12903 16727 12909
rect 16669 12900 16681 12903
rect 14976 12872 16681 12900
rect 14976 12860 14982 12872
rect 16669 12869 16681 12872
rect 16715 12869 16727 12903
rect 16669 12863 16727 12869
rect 16942 12792 16948 12844
rect 17000 12832 17006 12844
rect 17221 12835 17279 12841
rect 17221 12832 17233 12835
rect 17000 12804 17233 12832
rect 17000 12792 17006 12804
rect 17221 12801 17233 12804
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 11839 12736 13676 12764
rect 11839 12733 11851 12736
rect 11793 12727 11851 12733
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 14332 12736 18061 12764
rect 14332 12724 14338 12736
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 3421 12699 3479 12705
rect 3421 12665 3433 12699
rect 3467 12696 3479 12699
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 3467 12668 6653 12696
rect 3467 12665 3479 12668
rect 3421 12659 3479 12665
rect 6641 12665 6653 12668
rect 6687 12665 6699 12699
rect 7098 12696 7104 12708
rect 6641 12659 6699 12665
rect 6840 12668 7104 12696
rect 6840 12637 6868 12668
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 11054 12656 11060 12708
rect 11112 12696 11118 12708
rect 15746 12696 15752 12708
rect 11112 12668 15752 12696
rect 11112 12656 11118 12668
rect 15746 12656 15752 12668
rect 15804 12656 15810 12708
rect 6825 12631 6883 12637
rect 6825 12597 6837 12631
rect 6871 12597 6883 12631
rect 6825 12591 6883 12597
rect 7193 12631 7251 12637
rect 7193 12597 7205 12631
rect 7239 12628 7251 12631
rect 7834 12628 7840 12640
rect 7239 12600 7840 12628
rect 7239 12597 7251 12600
rect 7193 12591 7251 12597
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 8202 12628 8208 12640
rect 8163 12600 8208 12628
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 8297 12631 8355 12637
rect 8297 12597 8309 12631
rect 8343 12628 8355 12631
rect 9030 12628 9036 12640
rect 8343 12600 9036 12628
rect 8343 12597 8355 12600
rect 8297 12591 8355 12597
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 9306 12628 9312 12640
rect 9267 12600 9312 12628
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 9674 12628 9680 12640
rect 9635 12600 9680 12628
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 9769 12631 9827 12637
rect 9769 12597 9781 12631
rect 9815 12628 9827 12631
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 9815 12600 10333 12628
rect 9815 12597 9827 12600
rect 9769 12591 9827 12597
rect 10321 12597 10333 12600
rect 10367 12597 10379 12631
rect 10686 12628 10692 12640
rect 10647 12600 10692 12628
rect 10321 12591 10379 12597
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 10781 12631 10839 12637
rect 10781 12597 10793 12631
rect 10827 12628 10839 12631
rect 11146 12628 11152 12640
rect 10827 12600 11152 12628
rect 10827 12597 10839 12600
rect 10781 12591 10839 12597
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 11698 12628 11704 12640
rect 11659 12600 11704 12628
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 15194 12628 15200 12640
rect 12584 12600 15200 12628
rect 12584 12588 12590 12600
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 17034 12628 17040 12640
rect 16995 12600 17040 12628
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 17126 12588 17132 12640
rect 17184 12628 17190 12640
rect 18230 12628 18236 12640
rect 17184 12600 17229 12628
rect 18191 12600 18236 12628
rect 17184 12588 17190 12600
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 1857 12427 1915 12433
rect 1857 12393 1869 12427
rect 1903 12424 1915 12427
rect 3237 12427 3295 12433
rect 3237 12424 3249 12427
rect 1903 12396 3249 12424
rect 1903 12393 1915 12396
rect 1857 12387 1915 12393
rect 3237 12393 3249 12396
rect 3283 12393 3295 12427
rect 3237 12387 3295 12393
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 7340 12396 7573 12424
rect 7340 12384 7346 12396
rect 7561 12393 7573 12396
rect 7607 12393 7619 12427
rect 8938 12424 8944 12436
rect 8899 12396 8944 12424
rect 7561 12387 7619 12393
rect 8938 12384 8944 12396
rect 8996 12384 9002 12436
rect 9033 12427 9091 12433
rect 9033 12393 9045 12427
rect 9079 12424 9091 12427
rect 9306 12424 9312 12436
rect 9079 12396 9312 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10137 12427 10195 12433
rect 10137 12393 10149 12427
rect 10183 12424 10195 12427
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 10183 12396 10701 12424
rect 10183 12393 10195 12396
rect 10137 12387 10195 12393
rect 10689 12393 10701 12396
rect 10735 12393 10747 12427
rect 10689 12387 10747 12393
rect 11238 12384 11244 12436
rect 11296 12424 11302 12436
rect 11701 12427 11759 12433
rect 11701 12424 11713 12427
rect 11296 12396 11713 12424
rect 11296 12384 11302 12396
rect 11701 12393 11713 12396
rect 11747 12393 11759 12427
rect 11701 12387 11759 12393
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 17313 12427 17371 12433
rect 17313 12424 17325 12427
rect 17092 12396 17325 12424
rect 17092 12384 17098 12396
rect 17313 12393 17325 12396
rect 17359 12393 17371 12427
rect 17770 12424 17776 12436
rect 17731 12396 17776 12424
rect 17313 12387 17371 12393
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 7929 12359 7987 12365
rect 7929 12356 7941 12359
rect 4120 12328 7941 12356
rect 4120 12316 4126 12328
rect 7929 12325 7941 12328
rect 7975 12356 7987 12359
rect 11609 12359 11667 12365
rect 11609 12356 11621 12359
rect 7975 12328 11621 12356
rect 7975 12325 7987 12328
rect 7929 12319 7987 12325
rect 11609 12325 11621 12328
rect 11655 12356 11667 12359
rect 12069 12359 12127 12365
rect 12069 12356 12081 12359
rect 11655 12328 12081 12356
rect 11655 12325 11667 12328
rect 11609 12319 11667 12325
rect 12069 12325 12081 12328
rect 12115 12325 12127 12359
rect 12069 12319 12127 12325
rect 2222 12288 2228 12300
rect 2183 12260 2228 12288
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 6172 12291 6230 12297
rect 6172 12257 6184 12291
rect 6218 12288 6230 12291
rect 8570 12288 8576 12300
rect 6218 12260 8576 12288
rect 6218 12257 6230 12260
rect 6172 12251 6230 12257
rect 2130 12180 2136 12232
rect 2188 12220 2194 12232
rect 2317 12223 2375 12229
rect 2317 12220 2329 12223
rect 2188 12192 2329 12220
rect 2188 12180 2194 12192
rect 2317 12189 2329 12192
rect 2363 12189 2375 12223
rect 2317 12183 2375 12189
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12220 2559 12223
rect 2682 12220 2688 12232
rect 2547 12192 2688 12220
rect 2547 12189 2559 12192
rect 2501 12183 2559 12189
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 3142 12180 3148 12232
rect 3200 12220 3206 12232
rect 3329 12223 3387 12229
rect 3329 12220 3341 12223
rect 3200 12192 3341 12220
rect 3200 12180 3206 12192
rect 3329 12189 3341 12192
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 3476 12192 3521 12220
rect 3476 12180 3482 12192
rect 5810 12180 5816 12232
rect 5868 12220 5874 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5868 12192 5917 12220
rect 5868 12180 5874 12192
rect 5905 12189 5917 12192
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 8128 12229 8156 12260
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 9180 12260 10057 12288
rect 9180 12248 9186 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 11054 12288 11060 12300
rect 11015 12260 11060 12288
rect 10045 12251 10103 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12288 11207 12291
rect 11974 12288 11980 12300
rect 11195 12260 11980 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 12158 12288 12164 12300
rect 12119 12260 12164 12288
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 13906 12288 13912 12300
rect 13867 12260 13912 12288
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 15562 12288 15568 12300
rect 15523 12260 15568 12288
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 16666 12288 16672 12300
rect 16627 12260 16672 12288
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 16761 12291 16819 12297
rect 16761 12257 16773 12291
rect 16807 12288 16819 12291
rect 17310 12288 17316 12300
rect 16807 12260 17316 12288
rect 16807 12257 16819 12260
rect 16761 12251 16819 12257
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 17494 12248 17500 12300
rect 17552 12288 17558 12300
rect 17681 12291 17739 12297
rect 17681 12288 17693 12291
rect 17552 12260 17693 12288
rect 17552 12248 17558 12260
rect 17681 12257 17693 12260
rect 17727 12257 17739 12291
rect 17681 12251 17739 12257
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 7892 12192 8033 12220
rect 7892 12180 7898 12192
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8938 12220 8944 12232
rect 8113 12183 8171 12189
rect 8404 12192 8944 12220
rect 2869 12155 2927 12161
rect 2869 12121 2881 12155
rect 2915 12152 2927 12155
rect 5626 12152 5632 12164
rect 2915 12124 5632 12152
rect 2915 12121 2927 12124
rect 2869 12115 2927 12121
rect 5626 12112 5632 12124
rect 5684 12112 5690 12164
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7285 12155 7343 12161
rect 7285 12152 7297 12155
rect 6972 12124 7297 12152
rect 6972 12112 6978 12124
rect 7285 12121 7297 12124
rect 7331 12152 7343 12155
rect 7374 12152 7380 12164
rect 7331 12124 7380 12152
rect 7331 12121 7343 12124
rect 7285 12115 7343 12121
rect 7374 12112 7380 12124
rect 7432 12112 7438 12164
rect 8036 12152 8064 12183
rect 8404 12152 8432 12192
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12220 9275 12223
rect 9398 12220 9404 12232
rect 9263 12192 9404 12220
rect 9263 12189 9275 12192
rect 9217 12183 9275 12189
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 10318 12220 10324 12232
rect 10231 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12220 10382 12232
rect 10870 12220 10876 12232
rect 10376 12192 10876 12220
rect 10376 12180 10382 12192
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 11238 12220 11244 12232
rect 11199 12192 11244 12220
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 12250 12180 12256 12232
rect 12308 12220 12314 12232
rect 14277 12223 14335 12229
rect 12308 12192 12353 12220
rect 12308 12180 12314 12192
rect 14277 12189 14289 12223
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 11609 12155 11667 12161
rect 8036 12124 8432 12152
rect 8496 12124 10916 12152
rect 4614 12044 4620 12096
rect 4672 12084 4678 12096
rect 8496 12084 8524 12124
rect 10888 12096 10916 12124
rect 11609 12121 11621 12155
rect 11655 12152 11667 12155
rect 14182 12152 14188 12164
rect 11655 12124 14188 12152
rect 11655 12121 11667 12124
rect 11609 12115 11667 12121
rect 14182 12112 14188 12124
rect 14240 12112 14246 12164
rect 4672 12056 8524 12084
rect 8573 12087 8631 12093
rect 4672 12044 4678 12056
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 10410 12084 10416 12096
rect 8619 12056 10416 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 10410 12044 10416 12056
rect 10468 12044 10474 12096
rect 10870 12044 10876 12096
rect 10928 12044 10934 12096
rect 11882 12044 11888 12096
rect 11940 12084 11946 12096
rect 14292 12084 14320 12183
rect 15378 12180 15384 12232
rect 15436 12220 15442 12232
rect 15749 12223 15807 12229
rect 15749 12220 15761 12223
rect 15436 12192 15761 12220
rect 15436 12180 15442 12192
rect 15749 12189 15761 12192
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 16945 12223 17003 12229
rect 16945 12189 16957 12223
rect 16991 12220 17003 12223
rect 17034 12220 17040 12232
rect 16991 12192 17040 12220
rect 16991 12189 17003 12192
rect 16945 12183 17003 12189
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 17862 12180 17868 12232
rect 17920 12220 17926 12232
rect 17920 12192 17965 12220
rect 17920 12180 17926 12192
rect 15562 12112 15568 12164
rect 15620 12152 15626 12164
rect 17678 12152 17684 12164
rect 15620 12124 17684 12152
rect 15620 12112 15626 12124
rect 17678 12112 17684 12124
rect 17736 12112 17742 12164
rect 16298 12084 16304 12096
rect 11940 12056 14320 12084
rect 16259 12056 16304 12084
rect 11940 12044 11946 12056
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 2130 11880 2136 11892
rect 2091 11852 2136 11880
rect 2130 11840 2136 11852
rect 2188 11840 2194 11892
rect 3142 11880 3148 11892
rect 3103 11852 3148 11880
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 4614 11880 4620 11892
rect 4575 11852 4620 11880
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 8846 11880 8852 11892
rect 6196 11852 8708 11880
rect 8807 11852 8852 11880
rect 3234 11812 3240 11824
rect 2516 11784 3240 11812
rect 2516 11685 2544 11784
rect 3234 11772 3240 11784
rect 3292 11772 3298 11824
rect 3602 11772 3608 11824
rect 3660 11812 3666 11824
rect 5994 11812 6000 11824
rect 3660 11784 6000 11812
rect 3660 11772 3666 11784
rect 5994 11772 6000 11784
rect 6052 11772 6058 11824
rect 2685 11747 2743 11753
rect 2685 11744 2697 11747
rect 2608 11716 2697 11744
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11645 2559 11679
rect 2501 11639 2559 11645
rect 2406 11568 2412 11620
rect 2464 11608 2470 11620
rect 2608 11608 2636 11716
rect 2685 11713 2697 11716
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11713 3755 11747
rect 5258 11744 5264 11756
rect 5219 11716 5264 11744
rect 3697 11707 3755 11713
rect 3712 11676 3740 11707
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 6196 11753 6224 11852
rect 6825 11815 6883 11821
rect 6825 11781 6837 11815
rect 6871 11812 6883 11815
rect 7650 11812 7656 11824
rect 6871 11784 7656 11812
rect 6871 11781 6883 11784
rect 6825 11775 6883 11781
rect 7650 11772 7656 11784
rect 7708 11772 7714 11824
rect 7745 11815 7803 11821
rect 7745 11781 7757 11815
rect 7791 11812 7803 11815
rect 7837 11815 7895 11821
rect 7837 11812 7849 11815
rect 7791 11784 7849 11812
rect 7791 11781 7803 11784
rect 7745 11775 7803 11781
rect 7837 11781 7849 11784
rect 7883 11781 7895 11815
rect 8680 11812 8708 11852
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 8938 11840 8944 11892
rect 8996 11880 9002 11892
rect 10686 11880 10692 11892
rect 8996 11852 10456 11880
rect 10647 11852 10692 11880
rect 8996 11840 9002 11852
rect 9674 11812 9680 11824
rect 8680 11784 9680 11812
rect 7837 11775 7895 11781
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11713 6239 11747
rect 6362 11744 6368 11756
rect 6275 11716 6368 11744
rect 6181 11707 6239 11713
rect 6362 11704 6368 11716
rect 6420 11744 6426 11756
rect 6914 11744 6920 11756
rect 6420 11716 6920 11744
rect 6420 11704 6426 11716
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 7466 11744 7472 11756
rect 7427 11716 7472 11744
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 8018 11704 8024 11756
rect 8076 11744 8082 11756
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 8076 11716 8309 11744
rect 8076 11704 8082 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11744 8539 11747
rect 8570 11744 8576 11756
rect 8527 11716 8576 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 5074 11676 5080 11688
rect 2700 11648 3740 11676
rect 5035 11648 5080 11676
rect 2700 11620 2728 11648
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 6089 11679 6147 11685
rect 6089 11645 6101 11679
rect 6135 11676 6147 11679
rect 6270 11676 6276 11688
rect 6135 11648 6276 11676
rect 6135 11645 6147 11648
rect 6089 11639 6147 11645
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 7374 11636 7380 11688
rect 7432 11676 7438 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 7432 11648 7757 11676
rect 7432 11636 7438 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8496 11676 8524 11707
rect 8570 11704 8576 11716
rect 8628 11744 8634 11756
rect 9401 11747 9459 11753
rect 9401 11744 9413 11747
rect 8628 11716 9413 11744
rect 8628 11704 8634 11716
rect 9401 11713 9413 11716
rect 9447 11713 9459 11747
rect 10428 11744 10456 11852
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 13173 11883 13231 11889
rect 13173 11849 13185 11883
rect 13219 11880 13231 11883
rect 13906 11880 13912 11892
rect 13219 11852 13912 11880
rect 13219 11849 13231 11852
rect 13173 11843 13231 11849
rect 13906 11840 13912 11852
rect 13964 11880 13970 11892
rect 15194 11880 15200 11892
rect 13964 11852 15200 11880
rect 13964 11840 13970 11852
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 15657 11883 15715 11889
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 19426 11880 19432 11892
rect 15703 11852 19432 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 12066 11812 12072 11824
rect 11164 11784 12072 11812
rect 11164 11753 11192 11784
rect 12066 11772 12072 11784
rect 12124 11812 12130 11824
rect 14458 11812 14464 11824
rect 12124 11784 14464 11812
rect 12124 11772 12130 11784
rect 14458 11772 14464 11784
rect 14516 11772 14522 11824
rect 15562 11812 15568 11824
rect 14660 11784 15568 11812
rect 11149 11747 11207 11753
rect 10428 11716 11100 11744
rect 9401 11707 9459 11713
rect 8260 11648 8524 11676
rect 8260 11636 8266 11648
rect 8662 11636 8668 11688
rect 8720 11676 8726 11688
rect 10962 11676 10968 11688
rect 8720 11648 10968 11676
rect 8720 11636 8726 11648
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11072 11676 11100 11716
rect 11149 11713 11161 11747
rect 11195 11713 11207 11747
rect 11330 11744 11336 11756
rect 11291 11716 11336 11744
rect 11149 11707 11207 11713
rect 11330 11704 11336 11716
rect 11388 11704 11394 11756
rect 13170 11704 13176 11756
rect 13228 11744 13234 11756
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 13228 11716 13921 11744
rect 13228 11704 13234 11716
rect 13909 11713 13921 11716
rect 13955 11713 13967 11747
rect 13909 11707 13967 11713
rect 14660 11676 14688 11784
rect 15562 11772 15568 11784
rect 15620 11772 15626 11824
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15841 11747 15899 11753
rect 15841 11744 15853 11747
rect 14792 11716 15853 11744
rect 14792 11704 14798 11716
rect 15841 11713 15853 11716
rect 15887 11713 15899 11747
rect 17494 11744 17500 11756
rect 17455 11716 17500 11744
rect 15841 11707 15899 11713
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 11072 11648 14688 11676
rect 15010 11636 15016 11688
rect 15068 11676 15074 11688
rect 15105 11679 15163 11685
rect 15105 11676 15117 11679
rect 15068 11648 15117 11676
rect 15068 11636 15074 11648
rect 15105 11645 15117 11648
rect 15151 11676 15163 11679
rect 15151 11648 16804 11676
rect 15151 11645 15163 11648
rect 15105 11639 15163 11645
rect 16776 11620 16804 11648
rect 16850 11636 16856 11688
rect 16908 11676 16914 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 16908 11648 18061 11676
rect 16908 11636 16914 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 2464 11580 2636 11608
rect 2464 11568 2470 11580
rect 2682 11568 2688 11620
rect 2740 11568 2746 11620
rect 3513 11611 3571 11617
rect 3513 11577 3525 11611
rect 3559 11608 3571 11611
rect 5350 11608 5356 11620
rect 3559 11580 5356 11608
rect 3559 11577 3571 11580
rect 3513 11571 3571 11577
rect 5350 11568 5356 11580
rect 5408 11568 5414 11620
rect 5552 11580 6040 11608
rect 2590 11540 2596 11552
rect 2551 11512 2596 11540
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 3660 11512 3705 11540
rect 3660 11500 3666 11512
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 4120 11512 4997 11540
rect 4120 11500 4126 11512
rect 4985 11509 4997 11512
rect 5031 11540 5043 11543
rect 5552 11540 5580 11580
rect 5718 11540 5724 11552
rect 5031 11512 5580 11540
rect 5679 11512 5724 11540
rect 5031 11509 5043 11512
rect 4985 11503 5043 11509
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 6012 11540 6040 11580
rect 6638 11568 6644 11620
rect 6696 11608 6702 11620
rect 7193 11611 7251 11617
rect 7193 11608 7205 11611
rect 6696 11580 7205 11608
rect 6696 11568 6702 11580
rect 7193 11577 7205 11580
rect 7239 11577 7251 11611
rect 7193 11571 7251 11577
rect 7282 11568 7288 11620
rect 7340 11608 7346 11620
rect 7340 11580 7385 11608
rect 7944 11580 8340 11608
rect 7340 11568 7346 11580
rect 7944 11540 7972 11580
rect 6012 11512 7972 11540
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 8076 11512 8217 11540
rect 8076 11500 8082 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8312 11540 8340 11580
rect 8570 11568 8576 11620
rect 8628 11608 8634 11620
rect 9309 11611 9367 11617
rect 9309 11608 9321 11611
rect 8628 11580 9321 11608
rect 8628 11568 8634 11580
rect 9309 11577 9321 11580
rect 9355 11608 9367 11611
rect 11422 11608 11428 11620
rect 9355 11580 11428 11608
rect 9355 11577 9367 11580
rect 9309 11571 9367 11577
rect 11422 11568 11428 11580
rect 11480 11568 11486 11620
rect 12618 11568 12624 11620
rect 12676 11608 12682 11620
rect 13630 11608 13636 11620
rect 12676 11580 13636 11608
rect 12676 11568 12682 11580
rect 13630 11568 13636 11580
rect 13688 11568 13694 11620
rect 13725 11611 13783 11617
rect 13725 11577 13737 11611
rect 13771 11608 13783 11611
rect 15286 11608 15292 11620
rect 13771 11580 15292 11608
rect 13771 11577 13783 11580
rect 13725 11571 13783 11577
rect 15286 11568 15292 11580
rect 15344 11568 15350 11620
rect 15381 11611 15439 11617
rect 15381 11577 15393 11611
rect 15427 11608 15439 11611
rect 15657 11611 15715 11617
rect 15657 11608 15669 11611
rect 15427 11580 15669 11608
rect 15427 11577 15439 11580
rect 15381 11571 15439 11577
rect 15657 11577 15669 11580
rect 15703 11577 15715 11611
rect 15657 11571 15715 11577
rect 16108 11611 16166 11617
rect 16108 11577 16120 11611
rect 16154 11608 16166 11611
rect 16574 11608 16580 11620
rect 16154 11580 16580 11608
rect 16154 11577 16166 11580
rect 16108 11571 16166 11577
rect 16574 11568 16580 11580
rect 16632 11568 16638 11620
rect 16758 11568 16764 11620
rect 16816 11568 16822 11620
rect 8938 11540 8944 11552
rect 8312 11512 8944 11540
rect 8205 11503 8263 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9214 11540 9220 11552
rect 9175 11512 9220 11540
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 9640 11512 11069 11540
rect 9640 11500 9646 11512
rect 11057 11509 11069 11512
rect 11103 11540 11115 11543
rect 13173 11543 13231 11549
rect 13173 11540 13185 11543
rect 11103 11512 13185 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 13173 11509 13185 11512
rect 13219 11509 13231 11543
rect 13354 11540 13360 11552
rect 13315 11512 13360 11540
rect 13173 11503 13231 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 13872 11512 13917 11540
rect 13872 11500 13878 11512
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 17092 11512 17233 11540
rect 17092 11500 17098 11512
rect 17221 11509 17233 11512
rect 17267 11509 17279 11543
rect 17221 11503 17279 11509
rect 17770 11500 17776 11552
rect 17828 11540 17834 11552
rect 18233 11543 18291 11549
rect 18233 11540 18245 11543
rect 17828 11512 18245 11540
rect 17828 11500 17834 11512
rect 18233 11509 18245 11512
rect 18279 11509 18291 11543
rect 18233 11503 18291 11509
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 2682 11336 2688 11348
rect 2372 11308 2688 11336
rect 2372 11296 2378 11308
rect 2682 11296 2688 11308
rect 2740 11336 2746 11348
rect 3513 11339 3571 11345
rect 3513 11336 3525 11339
rect 2740 11308 3525 11336
rect 2740 11296 2746 11308
rect 3513 11305 3525 11308
rect 3559 11305 3571 11339
rect 3513 11299 3571 11305
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 7469 11339 7527 11345
rect 5776 11308 7420 11336
rect 5776 11296 5782 11308
rect 5988 11271 6046 11277
rect 2148 11240 4108 11268
rect 1394 11160 1400 11212
rect 1452 11200 1458 11212
rect 2148 11209 2176 11240
rect 2406 11209 2412 11212
rect 2133 11203 2191 11209
rect 2133 11200 2145 11203
rect 1452 11172 2145 11200
rect 1452 11160 1458 11172
rect 2133 11169 2145 11172
rect 2179 11169 2191 11203
rect 2400 11200 2412 11209
rect 2367 11172 2412 11200
rect 2133 11163 2191 11169
rect 2400 11163 2412 11172
rect 2406 11160 2412 11163
rect 2464 11160 2470 11212
rect 4080 11209 4108 11240
rect 5988 11237 6000 11271
rect 6034 11268 6046 11271
rect 6362 11268 6368 11280
rect 6034 11240 6368 11268
rect 6034 11237 6046 11240
rect 5988 11231 6046 11237
rect 6362 11228 6368 11240
rect 6420 11228 6426 11280
rect 7392 11268 7420 11308
rect 7469 11305 7481 11339
rect 7515 11336 7527 11339
rect 9214 11336 9220 11348
rect 7515 11308 9220 11336
rect 7515 11305 7527 11308
rect 7469 11299 7527 11305
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 10594 11336 10600 11348
rect 9876 11308 10600 11336
rect 9876 11268 9904 11308
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 11057 11339 11115 11345
rect 11057 11305 11069 11339
rect 11103 11305 11115 11339
rect 11057 11299 11115 11305
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 11698 11336 11704 11348
rect 11379 11308 11704 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 7392 11240 9904 11268
rect 9944 11271 10002 11277
rect 9944 11237 9956 11271
rect 9990 11268 10002 11271
rect 10318 11268 10324 11280
rect 9990 11240 10324 11268
rect 9990 11237 10002 11240
rect 9944 11231 10002 11237
rect 10318 11228 10324 11240
rect 10376 11228 10382 11280
rect 4065 11203 4123 11209
rect 4065 11169 4077 11203
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 4332 11203 4390 11209
rect 4332 11169 4344 11203
rect 4378 11200 4390 11203
rect 4706 11200 4712 11212
rect 4378 11172 4712 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5721 11203 5779 11209
rect 5721 11169 5733 11203
rect 5767 11200 5779 11203
rect 5810 11200 5816 11212
rect 5767 11172 5816 11200
rect 5767 11169 5779 11172
rect 5721 11163 5779 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 8018 11200 8024 11212
rect 7432 11172 8024 11200
rect 7432 11160 7438 11172
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 8196 11203 8254 11209
rect 8196 11169 8208 11203
rect 8242 11200 8254 11203
rect 10686 11200 10692 11212
rect 8242 11172 10692 11200
rect 8242 11169 8254 11172
rect 8196 11163 8254 11169
rect 10686 11160 10692 11172
rect 10744 11200 10750 11212
rect 11072 11200 11100 11299
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 17126 11296 17132 11348
rect 17184 11336 17190 11348
rect 17221 11339 17279 11345
rect 17221 11336 17233 11339
rect 17184 11308 17233 11336
rect 17184 11296 17190 11308
rect 17221 11305 17233 11308
rect 17267 11305 17279 11339
rect 17221 11299 17279 11305
rect 12713 11271 12771 11277
rect 12713 11237 12725 11271
rect 12759 11268 12771 11271
rect 13998 11268 14004 11280
rect 12759 11240 14004 11268
rect 12759 11237 12771 11240
rect 12713 11231 12771 11237
rect 13998 11228 14004 11240
rect 14056 11228 14062 11280
rect 14182 11228 14188 11280
rect 14240 11268 14246 11280
rect 17589 11271 17647 11277
rect 17589 11268 17601 11271
rect 14240 11240 17601 11268
rect 14240 11228 14246 11240
rect 17589 11237 17601 11240
rect 17635 11237 17647 11271
rect 17589 11231 17647 11237
rect 10744 11172 11100 11200
rect 10744 11160 10750 11172
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 13538 11209 13544 11212
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 11388 11172 12633 11200
rect 11388 11160 11394 11172
rect 12621 11169 12633 11172
rect 12667 11169 12679 11203
rect 13532 11200 13544 11209
rect 13499 11172 13544 11200
rect 12621 11163 12679 11169
rect 13532 11163 13544 11172
rect 13538 11160 13544 11163
rect 13596 11160 13602 11212
rect 15562 11209 15568 11212
rect 15556 11200 15568 11209
rect 15212 11172 15568 11200
rect 1670 11132 1676 11144
rect 1631 11104 1676 11132
rect 1670 11092 1676 11104
rect 1728 11092 1734 11144
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 6972 11104 7941 11132
rect 6972 11092 6978 11104
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9490 11132 9496 11144
rect 9272 11104 9496 11132
rect 9272 11092 9278 11104
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11132 12955 11135
rect 13170 11132 13176 11144
rect 12943 11104 13176 11132
rect 12943 11101 12955 11104
rect 12897 11095 12955 11101
rect 5442 11064 5448 11076
rect 5403 11036 5448 11064
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 7558 11064 7564 11076
rect 7147 11036 7564 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 9309 11067 9367 11073
rect 9309 11033 9321 11067
rect 9355 11064 9367 11067
rect 9398 11064 9404 11076
rect 9355 11036 9404 11064
rect 9355 11033 9367 11036
rect 9309 11027 9367 11033
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 8570 10996 8576 11008
rect 3844 10968 8576 10996
rect 3844 10956 3850 10968
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 9692 10996 9720 11095
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11790 11064 11796 11076
rect 11020 11036 11796 11064
rect 11020 11024 11026 11036
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 10686 10996 10692 11008
rect 9692 10968 10692 10996
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 11606 10956 11612 11008
rect 11664 10996 11670 11008
rect 12253 10999 12311 11005
rect 12253 10996 12265 10999
rect 11664 10968 12265 10996
rect 11664 10956 11670 10968
rect 12253 10965 12265 10968
rect 12299 10965 12311 10999
rect 13280 10996 13308 11095
rect 14645 11067 14703 11073
rect 14645 11033 14657 11067
rect 14691 11064 14703 11067
rect 15212 11064 15240 11172
rect 15556 11163 15568 11172
rect 15562 11160 15568 11163
rect 15620 11160 15626 11212
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11101 15347 11135
rect 17678 11132 17684 11144
rect 17639 11104 17684 11132
rect 15289 11095 15347 11101
rect 14691 11036 15240 11064
rect 14691 11033 14703 11036
rect 14645 11027 14703 11033
rect 14734 10996 14740 11008
rect 13280 10968 14740 10996
rect 12253 10959 12311 10965
rect 14734 10956 14740 10968
rect 14792 10996 14798 11008
rect 15304 10996 15332 11095
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 17862 11132 17868 11144
rect 17823 11104 17868 11132
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 16574 11024 16580 11076
rect 16632 11064 16638 11076
rect 16669 11067 16727 11073
rect 16669 11064 16681 11067
rect 16632 11036 16681 11064
rect 16632 11024 16638 11036
rect 16669 11033 16681 11036
rect 16715 11064 16727 11067
rect 17880 11064 17908 11092
rect 16715 11036 17908 11064
rect 16715 11033 16727 11036
rect 16669 11027 16727 11033
rect 14792 10968 15332 10996
rect 14792 10956 14798 10968
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 2222 10792 2228 10804
rect 2179 10764 2228 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 3421 10795 3479 10801
rect 3421 10761 3433 10795
rect 3467 10792 3479 10795
rect 3602 10792 3608 10804
rect 3467 10764 3608 10792
rect 3467 10761 3479 10764
rect 3421 10755 3479 10761
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 5258 10792 5264 10804
rect 4304 10764 5264 10792
rect 4304 10752 4310 10764
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5350 10752 5356 10804
rect 5408 10792 5414 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 5408 10764 5457 10792
rect 5408 10752 5414 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 6825 10795 6883 10801
rect 6825 10761 6837 10795
rect 6871 10792 6883 10795
rect 9582 10792 9588 10804
rect 6871 10764 9588 10792
rect 6871 10761 6883 10764
rect 6825 10755 6883 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 9861 10795 9919 10801
rect 9861 10761 9873 10795
rect 9907 10792 9919 10795
rect 10318 10792 10324 10804
rect 9907 10764 10324 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 11146 10792 11152 10804
rect 11107 10764 11152 10792
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 13354 10792 13360 10804
rect 11808 10764 13360 10792
rect 3786 10724 3792 10736
rect 1596 10696 3792 10724
rect 1596 10597 1624 10696
rect 3786 10684 3792 10696
rect 3844 10684 3850 10736
rect 4080 10696 5488 10724
rect 2406 10616 2412 10668
rect 2464 10656 2470 10668
rect 4080 10665 4108 10696
rect 5460 10668 5488 10696
rect 6270 10684 6276 10736
rect 6328 10724 6334 10736
rect 6914 10724 6920 10736
rect 6328 10696 6920 10724
rect 6328 10684 6334 10696
rect 6914 10684 6920 10696
rect 6972 10724 6978 10736
rect 7837 10727 7895 10733
rect 7837 10724 7849 10727
rect 6972 10696 7849 10724
rect 6972 10684 6978 10696
rect 7837 10693 7849 10696
rect 7883 10724 7895 10727
rect 7883 10696 8524 10724
rect 7883 10693 7895 10696
rect 7837 10687 7895 10693
rect 2777 10659 2835 10665
rect 2777 10656 2789 10659
rect 2464 10628 2789 10656
rect 2464 10616 2470 10628
rect 2777 10625 2789 10628
rect 2823 10656 2835 10659
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 2823 10628 4077 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4706 10616 4712 10668
rect 4764 10656 4770 10668
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 4764 10628 4997 10656
rect 4764 10616 4770 10628
rect 4985 10625 4997 10628
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5500 10628 6009 10656
rect 5500 10616 5506 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6362 10616 6368 10668
rect 6420 10656 6426 10668
rect 6420 10628 6960 10656
rect 6420 10616 6426 10628
rect 1581 10591 1639 10597
rect 1581 10557 1593 10591
rect 1627 10557 1639 10591
rect 1581 10551 1639 10557
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 2501 10591 2559 10597
rect 2501 10588 2513 10591
rect 1728 10560 2513 10588
rect 1728 10548 1734 10560
rect 2501 10557 2513 10560
rect 2547 10557 2559 10591
rect 5534 10588 5540 10600
rect 2501 10551 2559 10557
rect 3712 10560 5540 10588
rect 2866 10520 2872 10532
rect 1780 10492 2872 10520
rect 1780 10461 1808 10492
rect 2866 10480 2872 10492
rect 2924 10480 2930 10532
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10421 1823 10455
rect 1765 10415 1823 10421
rect 2593 10455 2651 10461
rect 2593 10421 2605 10455
rect 2639 10452 2651 10455
rect 3712 10452 3740 10560
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 5902 10588 5908 10600
rect 5863 10560 5908 10588
rect 5902 10548 5908 10560
rect 5960 10548 5966 10600
rect 3789 10523 3847 10529
rect 3789 10489 3801 10523
rect 3835 10520 3847 10523
rect 4893 10523 4951 10529
rect 3835 10492 4476 10520
rect 3835 10489 3847 10492
rect 3789 10483 3847 10489
rect 3878 10452 3884 10464
rect 2639 10424 3740 10452
rect 3839 10424 3884 10452
rect 2639 10421 2651 10424
rect 2593 10415 2651 10421
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 4448 10461 4476 10492
rect 4893 10489 4905 10523
rect 4939 10520 4951 10523
rect 5350 10520 5356 10532
rect 4939 10492 5356 10520
rect 4939 10489 4951 10492
rect 4893 10483 4951 10489
rect 5350 10480 5356 10492
rect 5408 10480 5414 10532
rect 5718 10480 5724 10532
rect 5776 10520 5782 10532
rect 5813 10523 5871 10529
rect 5813 10520 5825 10523
rect 5776 10492 5825 10520
rect 5776 10480 5782 10492
rect 5813 10489 5825 10492
rect 5859 10489 5871 10523
rect 5813 10483 5871 10489
rect 6546 10480 6552 10532
rect 6604 10520 6610 10532
rect 6932 10520 6960 10628
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 7156 10628 7389 10656
rect 7156 10616 7162 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 8496 10665 8524 10696
rect 9490 10684 9496 10736
rect 9548 10724 9554 10736
rect 11238 10724 11244 10736
rect 9548 10696 11244 10724
rect 9548 10684 9554 10696
rect 11238 10684 11244 10696
rect 11296 10724 11302 10736
rect 11296 10696 11744 10724
rect 11296 10684 11302 10696
rect 8481 10659 8539 10665
rect 7616 10628 8248 10656
rect 7616 10616 7622 10628
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10588 7251 10591
rect 7282 10588 7288 10600
rect 7239 10560 7288 10588
rect 7239 10557 7251 10560
rect 7193 10551 7251 10557
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 8036 10520 8064 10551
rect 6604 10492 6776 10520
rect 6932 10492 8064 10520
rect 8220 10520 8248 10628
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 9858 10656 9864 10668
rect 9732 10628 9864 10656
rect 9732 10616 9738 10628
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 10594 10656 10600 10668
rect 10555 10628 10600 10656
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 9953 10591 10011 10597
rect 8588 10560 8892 10588
rect 8588 10520 8616 10560
rect 8220 10492 8616 10520
rect 8748 10523 8806 10529
rect 6604 10480 6610 10492
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10421 4491 10455
rect 4798 10452 4804 10464
rect 4759 10424 4804 10452
rect 4433 10415 4491 10421
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 6748 10452 6776 10492
rect 8748 10489 8760 10523
rect 8794 10489 8806 10523
rect 8864 10520 8892 10560
rect 9953 10557 9965 10591
rect 9999 10588 10011 10591
rect 10318 10588 10324 10600
rect 9999 10560 10324 10588
rect 9999 10557 10011 10560
rect 9953 10551 10011 10557
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 10502 10588 10508 10600
rect 10463 10560 10508 10588
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10704 10520 10732 10619
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 11716 10665 11744 10696
rect 11609 10659 11667 10665
rect 11609 10656 11621 10659
rect 11480 10628 11621 10656
rect 11480 10616 11486 10628
rect 11609 10625 11621 10628
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 11808 10588 11836 10764
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 13722 10752 13728 10804
rect 13780 10792 13786 10804
rect 13780 10764 15700 10792
rect 13780 10752 13786 10764
rect 15672 10724 15700 10764
rect 16666 10752 16672 10804
rect 16724 10792 16730 10804
rect 16945 10795 17003 10801
rect 16945 10792 16957 10795
rect 16724 10764 16957 10792
rect 16724 10752 16730 10764
rect 16945 10761 16957 10764
rect 16991 10761 17003 10795
rect 16945 10755 17003 10761
rect 15672 10696 18092 10724
rect 16850 10656 16856 10668
rect 15764 10628 16856 10656
rect 11296 10560 11836 10588
rect 11296 10548 11302 10560
rect 12158 10548 12164 10600
rect 12216 10588 12222 10600
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 12216 10560 12449 10588
rect 12216 10548 12222 10560
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 12704 10591 12762 10597
rect 12704 10557 12716 10591
rect 12750 10588 12762 10591
rect 13170 10588 13176 10600
rect 12750 10560 13176 10588
rect 12750 10557 12762 10560
rect 12704 10551 12762 10557
rect 13170 10548 13176 10560
rect 13228 10588 13234 10600
rect 13446 10588 13452 10600
rect 13228 10560 13452 10588
rect 13228 10548 13234 10560
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 14182 10588 14188 10600
rect 14143 10560 14188 10588
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 14734 10588 14740 10600
rect 14695 10560 14740 10588
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 15764 10588 15792 10628
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 17402 10656 17408 10668
rect 17363 10628 17408 10656
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 17589 10659 17647 10665
rect 17589 10625 17601 10659
rect 17635 10656 17647 10659
rect 17862 10656 17868 10668
rect 17635 10628 17868 10656
rect 17635 10625 17647 10628
rect 17589 10619 17647 10625
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 14936 10560 15792 10588
rect 8864 10492 10732 10520
rect 8748 10483 8806 10489
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 6748 10424 7297 10452
rect 7285 10421 7297 10424
rect 7331 10421 7343 10455
rect 7285 10415 7343 10421
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 8018 10452 8024 10464
rect 7800 10424 8024 10452
rect 7800 10412 7806 10424
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 8772 10452 8800 10483
rect 11790 10480 11796 10532
rect 11848 10520 11854 10532
rect 14936 10520 14964 10560
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 16393 10591 16451 10597
rect 16393 10588 16405 10591
rect 15896 10560 16405 10588
rect 15896 10548 15902 10560
rect 16393 10557 16405 10560
rect 16439 10557 16451 10591
rect 16393 10551 16451 10557
rect 16482 10548 16488 10600
rect 16540 10588 16546 10600
rect 17494 10588 17500 10600
rect 16540 10560 17500 10588
rect 16540 10548 16546 10560
rect 17494 10548 17500 10560
rect 17552 10548 17558 10600
rect 18064 10597 18092 10696
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 11848 10492 14964 10520
rect 15004 10523 15062 10529
rect 11848 10480 11854 10492
rect 15004 10489 15016 10523
rect 15050 10520 15062 10523
rect 17034 10520 17040 10532
rect 15050 10492 17040 10520
rect 15050 10489 15062 10492
rect 15004 10483 15062 10489
rect 17034 10480 17040 10492
rect 17092 10480 17098 10532
rect 8846 10452 8852 10464
rect 8772 10424 8852 10452
rect 8846 10412 8852 10424
rect 8904 10452 8910 10464
rect 9490 10452 9496 10464
rect 8904 10424 9496 10452
rect 8904 10412 8910 10424
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 9953 10455 10011 10461
rect 9953 10452 9965 10455
rect 9732 10424 9965 10452
rect 9732 10412 9738 10424
rect 9953 10421 9965 10424
rect 9999 10421 10011 10455
rect 9953 10415 10011 10421
rect 10137 10455 10195 10461
rect 10137 10421 10149 10455
rect 10183 10452 10195 10455
rect 10502 10452 10508 10464
rect 10183 10424 10508 10452
rect 10183 10421 10195 10424
rect 10137 10415 10195 10421
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 11422 10412 11428 10464
rect 11480 10452 11486 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 11480 10424 11529 10452
rect 11480 10412 11486 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 11517 10415 11575 10421
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 13538 10452 13544 10464
rect 12768 10424 13544 10452
rect 12768 10412 12774 10424
rect 13538 10412 13544 10424
rect 13596 10452 13602 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13596 10424 13829 10452
rect 13596 10412 13602 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 14369 10455 14427 10461
rect 14369 10421 14381 10455
rect 14415 10452 14427 10455
rect 15194 10452 15200 10464
rect 14415 10424 15200 10452
rect 14415 10421 14427 10424
rect 14369 10415 14427 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 15470 10412 15476 10464
rect 15528 10452 15534 10464
rect 15838 10452 15844 10464
rect 15528 10424 15844 10452
rect 15528 10412 15534 10424
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 16022 10412 16028 10464
rect 16080 10452 16086 10464
rect 16117 10455 16175 10461
rect 16117 10452 16129 10455
rect 16080 10424 16129 10452
rect 16080 10412 16086 10424
rect 16117 10421 16129 10424
rect 16163 10421 16175 10455
rect 16574 10452 16580 10464
rect 16535 10424 16580 10452
rect 16117 10415 16175 10421
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 17313 10455 17371 10461
rect 17313 10452 17325 10455
rect 16724 10424 17325 10452
rect 16724 10412 16730 10424
rect 17313 10421 17325 10424
rect 17359 10421 17371 10455
rect 17313 10415 17371 10421
rect 18233 10455 18291 10461
rect 18233 10421 18245 10455
rect 18279 10452 18291 10455
rect 18414 10452 18420 10464
rect 18279 10424 18420 10452
rect 18279 10421 18291 10424
rect 18233 10415 18291 10421
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 2958 10248 2964 10260
rect 2823 10220 2964 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 2958 10208 2964 10220
rect 3016 10248 3022 10260
rect 3418 10248 3424 10260
rect 3016 10220 3424 10248
rect 3016 10208 3022 10220
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 3878 10208 3884 10260
rect 3936 10248 3942 10260
rect 4433 10251 4491 10257
rect 4433 10248 4445 10251
rect 3936 10220 4445 10248
rect 3936 10208 3942 10220
rect 4433 10217 4445 10220
rect 4479 10217 4491 10251
rect 4433 10211 4491 10217
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5994 10248 6000 10260
rect 5592 10220 6000 10248
rect 5592 10208 5598 10220
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6178 10208 6184 10260
rect 6236 10248 6242 10260
rect 6730 10248 6736 10260
rect 6236 10220 6736 10248
rect 6236 10208 6242 10220
rect 6730 10208 6736 10220
rect 6788 10248 6794 10260
rect 9674 10248 9680 10260
rect 6788 10220 9680 10248
rect 6788 10208 6794 10220
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 9968 10220 10149 10248
rect 1664 10183 1722 10189
rect 1664 10149 1676 10183
rect 1710 10180 1722 10183
rect 2314 10180 2320 10192
rect 1710 10152 2320 10180
rect 1710 10149 1722 10152
rect 1664 10143 1722 10149
rect 2314 10140 2320 10152
rect 2372 10140 2378 10192
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 6632 10183 6690 10189
rect 4120 10152 6592 10180
rect 4120 10140 4126 10152
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10112 1458 10124
rect 1946 10112 1952 10124
rect 1452 10084 1952 10112
rect 1452 10072 1458 10084
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 3050 10112 3056 10124
rect 3011 10084 3056 10112
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 5074 10112 5080 10124
rect 4847 10084 5080 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 5074 10072 5080 10084
rect 5132 10112 5138 10124
rect 5132 10084 5488 10112
rect 5132 10072 5138 10084
rect 4890 10044 4896 10056
rect 4851 10016 4896 10044
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 5460 10044 5488 10084
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 5629 10115 5687 10121
rect 5629 10112 5641 10115
rect 5592 10084 5641 10112
rect 5592 10072 5598 10084
rect 5629 10081 5641 10084
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 6270 10112 6276 10124
rect 5868 10084 6276 10112
rect 5868 10072 5874 10084
rect 6270 10072 6276 10084
rect 6328 10112 6334 10124
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 6328 10084 6377 10112
rect 6328 10072 6334 10084
rect 6365 10081 6377 10084
rect 6411 10081 6423 10115
rect 6564 10112 6592 10152
rect 6632 10149 6644 10183
rect 6678 10180 6690 10183
rect 6914 10180 6920 10192
rect 6678 10152 6920 10180
rect 6678 10149 6690 10152
rect 6632 10143 6690 10149
rect 6914 10140 6920 10152
rect 6972 10180 6978 10192
rect 7466 10180 7472 10192
rect 6972 10152 7472 10180
rect 6972 10140 6978 10152
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 8478 10180 8484 10192
rect 8439 10152 8484 10180
rect 8478 10140 8484 10152
rect 8536 10140 8542 10192
rect 8570 10140 8576 10192
rect 8628 10180 8634 10192
rect 9968 10180 9996 10220
rect 10137 10217 10149 10220
rect 10183 10217 10195 10251
rect 10137 10211 10195 10217
rect 10318 10208 10324 10260
rect 10376 10248 10382 10260
rect 11422 10248 11428 10260
rect 10376 10220 11428 10248
rect 10376 10208 10382 10220
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 11977 10251 12035 10257
rect 11977 10217 11989 10251
rect 12023 10248 12035 10251
rect 12710 10248 12716 10260
rect 12023 10220 12716 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 13504 10220 13553 10248
rect 13504 10208 13510 10220
rect 13541 10217 13553 10220
rect 13587 10217 13599 10251
rect 13541 10211 13599 10217
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13872 10220 13921 10248
rect 13872 10208 13878 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 14274 10248 14280 10260
rect 14235 10220 14280 10248
rect 13909 10211 13967 10217
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 14366 10208 14372 10260
rect 14424 10248 14430 10260
rect 15102 10248 15108 10260
rect 14424 10220 15108 10248
rect 14424 10208 14430 10220
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15286 10248 15292 10260
rect 15247 10220 15292 10248
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 16301 10251 16359 10257
rect 15488 10220 16252 10248
rect 8628 10152 9996 10180
rect 10045 10183 10103 10189
rect 8628 10140 8634 10152
rect 10045 10149 10057 10183
rect 10091 10149 10103 10183
rect 10045 10143 10103 10149
rect 8389 10115 8447 10121
rect 6564 10084 8340 10112
rect 6365 10075 6423 10081
rect 6178 10044 6184 10056
rect 5460 10016 6184 10044
rect 4985 10007 5043 10013
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 5000 9976 5028 10007
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 4764 9948 5028 9976
rect 5445 9979 5503 9985
rect 4764 9936 4770 9948
rect 5445 9945 5457 9979
rect 5491 9976 5503 9979
rect 6362 9976 6368 9988
rect 5491 9948 6368 9976
rect 5491 9945 5503 9948
rect 5445 9939 5503 9945
rect 3142 9868 3148 9920
rect 3200 9908 3206 9920
rect 3237 9911 3295 9917
rect 3237 9908 3249 9911
rect 3200 9880 3249 9908
rect 3200 9868 3206 9880
rect 3237 9877 3249 9880
rect 3283 9877 3295 9911
rect 3237 9871 3295 9877
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 5460 9908 5488 9939
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 7466 9936 7472 9988
rect 7524 9976 7530 9988
rect 8021 9979 8079 9985
rect 8021 9976 8033 9979
rect 7524 9948 8033 9976
rect 7524 9936 7530 9948
rect 8021 9945 8033 9948
rect 8067 9945 8079 9979
rect 8312 9976 8340 10084
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 9674 10112 9680 10124
rect 8435 10084 9680 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 9858 10072 9864 10124
rect 9916 10112 9922 10124
rect 10060 10112 10088 10143
rect 11238 10140 11244 10192
rect 11296 10180 11302 10192
rect 11517 10183 11575 10189
rect 11517 10180 11529 10183
rect 11296 10152 11529 10180
rect 11296 10140 11302 10152
rect 11517 10149 11529 10152
rect 11563 10149 11575 10183
rect 11517 10143 11575 10149
rect 11606 10140 11612 10192
rect 11664 10180 11670 10192
rect 11664 10152 11709 10180
rect 12360 10152 15148 10180
rect 11664 10140 11670 10152
rect 9916 10084 10088 10112
rect 10965 10115 11023 10121
rect 9916 10072 9922 10084
rect 10965 10081 10977 10115
rect 11011 10081 11023 10115
rect 12360 10112 12388 10152
rect 10965 10075 11023 10081
rect 11716 10084 12388 10112
rect 12428 10115 12486 10121
rect 8570 10044 8576 10056
rect 8531 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 9232 10016 10241 10044
rect 9122 9976 9128 9988
rect 8312 9948 9128 9976
rect 8021 9939 8079 9945
rect 9122 9936 9128 9948
rect 9180 9936 9186 9988
rect 4580 9880 5488 9908
rect 7745 9911 7803 9917
rect 4580 9868 4586 9880
rect 7745 9877 7757 9911
rect 7791 9908 7803 9911
rect 8202 9908 8208 9920
rect 7791 9880 8208 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 8202 9868 8208 9880
rect 8260 9908 8266 9920
rect 9232 9908 9260 10016
rect 10229 10013 10241 10016
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 9858 9976 9864 9988
rect 9548 9948 9864 9976
rect 9548 9936 9554 9948
rect 9858 9936 9864 9948
rect 9916 9936 9922 9988
rect 9950 9936 9956 9988
rect 10008 9936 10014 9988
rect 10686 9936 10692 9988
rect 10744 9976 10750 9988
rect 10781 9979 10839 9985
rect 10781 9976 10793 9979
rect 10744 9948 10793 9976
rect 10744 9936 10750 9948
rect 10781 9945 10793 9948
rect 10827 9945 10839 9979
rect 10980 9976 11008 10075
rect 11054 9976 11060 9988
rect 10967 9948 11060 9976
rect 10781 9939 10839 9945
rect 11054 9936 11060 9948
rect 11112 9976 11118 9988
rect 11716 9976 11744 10084
rect 12428 10081 12440 10115
rect 12474 10112 12486 10115
rect 13262 10112 13268 10124
rect 12474 10084 13268 10112
rect 12474 10081 12486 10084
rect 12428 10075 12486 10081
rect 13262 10072 13268 10084
rect 13320 10112 13326 10124
rect 14550 10112 14556 10124
rect 13320 10084 14556 10112
rect 13320 10072 13326 10084
rect 11793 10047 11851 10053
rect 11793 10013 11805 10047
rect 11839 10044 11851 10047
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 11839 10016 11989 10044
rect 11839 10013 11851 10016
rect 11793 10007 11851 10013
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 12158 10044 12164 10056
rect 12119 10016 12164 10044
rect 11977 10007 12035 10013
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 14274 10004 14280 10056
rect 14332 10044 14338 10056
rect 14476 10053 14504 10084
rect 14550 10072 14556 10084
rect 14608 10112 14614 10124
rect 15120 10121 15148 10152
rect 15105 10115 15163 10121
rect 14608 10084 14688 10112
rect 14608 10072 14614 10084
rect 14369 10047 14427 10053
rect 14369 10044 14381 10047
rect 14332 10016 14381 10044
rect 14332 10004 14338 10016
rect 14369 10013 14381 10016
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 11112 9948 11744 9976
rect 14660 9976 14688 10084
rect 15105 10081 15117 10115
rect 15151 10081 15163 10115
rect 15105 10075 15163 10081
rect 15286 10072 15292 10124
rect 15344 10112 15350 10124
rect 15488 10112 15516 10220
rect 15562 10140 15568 10192
rect 15620 10180 15626 10192
rect 15620 10152 15976 10180
rect 15620 10140 15626 10152
rect 15654 10112 15660 10124
rect 15344 10084 15516 10112
rect 15615 10084 15660 10112
rect 15344 10072 15350 10084
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 15746 10072 15752 10124
rect 15804 10112 15810 10124
rect 15804 10084 15849 10112
rect 15804 10072 15810 10084
rect 15562 10004 15568 10056
rect 15620 10044 15626 10056
rect 15764 10044 15792 10072
rect 15620 10016 15792 10044
rect 15841 10047 15899 10053
rect 15620 10004 15626 10016
rect 15841 10013 15853 10047
rect 15887 10013 15899 10047
rect 15948 10044 15976 10152
rect 16224 10112 16252 10220
rect 16301 10217 16313 10251
rect 16347 10248 16359 10251
rect 17773 10251 17831 10257
rect 17773 10248 17785 10251
rect 16347 10220 17785 10248
rect 16347 10217 16359 10220
rect 16301 10211 16359 10217
rect 17773 10217 17785 10220
rect 17819 10217 17831 10251
rect 17773 10211 17831 10217
rect 16669 10183 16727 10189
rect 16669 10149 16681 10183
rect 16715 10180 16727 10183
rect 16942 10180 16948 10192
rect 16715 10152 16948 10180
rect 16715 10149 16727 10152
rect 16669 10143 16727 10149
rect 16942 10140 16948 10152
rect 17000 10140 17006 10192
rect 16761 10115 16819 10121
rect 16761 10112 16773 10115
rect 16224 10084 16773 10112
rect 16761 10081 16773 10084
rect 16807 10081 16819 10115
rect 16761 10075 16819 10081
rect 17402 10072 17408 10124
rect 17460 10112 17466 10124
rect 17681 10115 17739 10121
rect 17681 10112 17693 10115
rect 17460 10084 17693 10112
rect 17460 10072 17466 10084
rect 17681 10081 17693 10084
rect 17727 10081 17739 10115
rect 17681 10075 17739 10081
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 15948 10016 16865 10044
rect 15841 10007 15899 10013
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 17862 10044 17868 10056
rect 17823 10016 17868 10044
rect 16853 10007 16911 10013
rect 14660 9948 15424 9976
rect 11112 9936 11118 9948
rect 8260 9880 9260 9908
rect 9677 9911 9735 9917
rect 8260 9868 8266 9880
rect 9677 9877 9689 9911
rect 9723 9908 9735 9911
rect 9968 9908 9996 9936
rect 9723 9880 9996 9908
rect 11149 9911 11207 9917
rect 9723 9877 9735 9880
rect 9677 9871 9735 9877
rect 11149 9877 11161 9911
rect 11195 9908 11207 9911
rect 11422 9908 11428 9920
rect 11195 9880 11428 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 14182 9908 14188 9920
rect 14056 9880 14188 9908
rect 14056 9868 14062 9880
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 14921 9911 14979 9917
rect 14921 9908 14933 9911
rect 14792 9880 14933 9908
rect 14792 9868 14798 9880
rect 14921 9877 14933 9880
rect 14967 9908 14979 9911
rect 15102 9908 15108 9920
rect 14967 9880 15108 9908
rect 14967 9877 14979 9880
rect 14921 9871 14979 9877
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 15396 9908 15424 9948
rect 15847 9908 15875 10007
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 16022 9936 16028 9988
rect 16080 9936 16086 9988
rect 17310 9976 17316 9988
rect 17271 9948 17316 9976
rect 17310 9936 17316 9948
rect 17368 9936 17374 9988
rect 15396 9880 15875 9908
rect 16040 9908 16068 9936
rect 16482 9908 16488 9920
rect 16040 9880 16488 9908
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 4706 9664 4712 9716
rect 4764 9664 4770 9716
rect 4985 9707 5043 9713
rect 4985 9673 4997 9707
rect 5031 9704 5043 9707
rect 6457 9707 6515 9713
rect 5031 9676 6040 9704
rect 5031 9673 5043 9676
rect 4985 9667 5043 9673
rect 4724 9577 4752 9664
rect 6012 9636 6040 9676
rect 6457 9673 6469 9707
rect 6503 9704 6515 9707
rect 6914 9704 6920 9716
rect 6503 9676 6920 9704
rect 6503 9673 6515 9676
rect 6457 9667 6515 9673
rect 6914 9664 6920 9676
rect 6972 9664 6978 9716
rect 8846 9704 8852 9716
rect 7484 9676 8432 9704
rect 8807 9676 8852 9704
rect 7484 9636 7512 9676
rect 6012 9608 7512 9636
rect 8404 9636 8432 9676
rect 8846 9664 8852 9676
rect 8904 9664 8910 9716
rect 9122 9664 9128 9716
rect 9180 9704 9186 9716
rect 10686 9704 10692 9716
rect 9180 9676 10692 9704
rect 9180 9664 9186 9676
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 11606 9664 11612 9716
rect 11664 9704 11670 9716
rect 13722 9704 13728 9716
rect 11664 9676 13728 9704
rect 11664 9664 11670 9676
rect 13722 9664 13728 9676
rect 13780 9664 13786 9716
rect 15010 9704 15016 9716
rect 13832 9676 15016 9704
rect 11054 9636 11060 9648
rect 8404 9608 8524 9636
rect 11015 9608 11060 9636
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 6328 9540 7481 9568
rect 6328 9528 6334 9540
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 8496 9568 8524 9608
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 11330 9636 11336 9648
rect 11291 9608 11336 9636
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 12621 9639 12679 9645
rect 12621 9605 12633 9639
rect 12667 9636 12679 9639
rect 13832 9636 13860 9676
rect 15010 9664 15016 9676
rect 15068 9664 15074 9716
rect 16482 9664 16488 9716
rect 16540 9704 16546 9716
rect 16540 9676 16620 9704
rect 16540 9664 16546 9676
rect 12667 9608 13860 9636
rect 14001 9639 14059 9645
rect 12667 9605 12679 9608
rect 12621 9599 12679 9605
rect 14001 9605 14013 9639
rect 14047 9605 14059 9639
rect 14001 9599 14059 9605
rect 11977 9571 12035 9577
rect 8496 9540 9260 9568
rect 7469 9531 7527 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9469 1455 9503
rect 1946 9500 1952 9512
rect 1907 9472 1952 9500
rect 1397 9463 1455 9469
rect 1412 9432 1440 9463
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 2216 9503 2274 9509
rect 2216 9469 2228 9503
rect 2262 9500 2274 9503
rect 2958 9500 2964 9512
rect 2262 9472 2964 9500
rect 2262 9469 2274 9472
rect 2216 9463 2274 9469
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 3789 9503 3847 9509
rect 3108 9472 3648 9500
rect 3108 9460 3114 9472
rect 3510 9432 3516 9444
rect 1412 9404 3516 9432
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 3620 9432 3648 9472
rect 3789 9469 3801 9503
rect 3835 9500 3847 9503
rect 4522 9500 4528 9512
rect 3835 9472 4528 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 4522 9460 4528 9472
rect 4580 9460 4586 9512
rect 5074 9500 5080 9512
rect 5035 9472 5080 9500
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9500 7251 9503
rect 7374 9500 7380 9512
rect 7239 9472 7380 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 8570 9500 8576 9512
rect 7576 9472 8576 9500
rect 4985 9435 5043 9441
rect 4985 9432 4997 9435
rect 3620 9404 4997 9432
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 3326 9364 3332 9376
rect 3287 9336 3332 9364
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 3605 9367 3663 9373
rect 3605 9333 3617 9367
rect 3651 9364 3663 9367
rect 3786 9364 3792 9376
rect 3651 9336 3792 9364
rect 3651 9333 3663 9336
rect 3605 9327 3663 9333
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 4062 9364 4068 9376
rect 4023 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4430 9364 4436 9376
rect 4391 9336 4436 9364
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4540 9373 4568 9404
rect 4985 9401 4997 9404
rect 5031 9401 5043 9435
rect 4985 9395 5043 9401
rect 5344 9435 5402 9441
rect 5344 9401 5356 9435
rect 5390 9432 5402 9435
rect 5442 9432 5448 9444
rect 5390 9404 5448 9432
rect 5390 9401 5402 9404
rect 5344 9395 5402 9401
rect 5442 9392 5448 9404
rect 5500 9432 5506 9444
rect 7576 9432 7604 9472
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9232 9500 9260 9540
rect 10152 9540 11836 9568
rect 10152 9500 10180 9540
rect 11238 9500 11244 9512
rect 9232 9472 10180 9500
rect 11199 9472 11244 9500
rect 9125 9463 9183 9469
rect 7742 9441 7748 9444
rect 7736 9432 7748 9441
rect 5500 9404 7604 9432
rect 7703 9404 7748 9432
rect 5500 9392 5506 9404
rect 7736 9395 7748 9404
rect 7742 9392 7748 9395
rect 7800 9392 7806 9444
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9333 4583 9367
rect 4525 9327 4583 9333
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 5592 9336 7021 9364
rect 5592 9324 5598 9336
rect 7009 9333 7021 9336
rect 7055 9333 7067 9367
rect 9140 9364 9168 9463
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11664 9472 11713 9500
rect 11664 9460 11670 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11808 9500 11836 9540
rect 11977 9537 11989 9571
rect 12023 9568 12035 9571
rect 13262 9568 13268 9580
rect 12023 9540 13268 9568
rect 12023 9537 12035 9540
rect 11977 9531 12035 9537
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13722 9568 13728 9580
rect 13587 9540 13728 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 14016 9568 14044 9599
rect 14090 9596 14096 9648
rect 14148 9636 14154 9648
rect 14148 9608 14872 9636
rect 14148 9596 14154 9608
rect 14182 9568 14188 9580
rect 14016 9540 14188 9568
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 14550 9568 14556 9580
rect 14511 9540 14556 9568
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 14844 9512 14872 9608
rect 15102 9528 15108 9580
rect 15160 9568 15166 9580
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 15160 9540 15577 9568
rect 15160 9528 15166 9540
rect 15565 9537 15577 9540
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 12066 9500 12072 9512
rect 11808 9472 12072 9500
rect 11701 9463 11759 9469
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12216 9472 12449 9500
rect 12216 9460 12222 9472
rect 12437 9469 12449 9472
rect 12483 9500 12495 9503
rect 12894 9500 12900 9512
rect 12483 9472 12900 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 14826 9460 14832 9512
rect 14884 9500 14890 9512
rect 15838 9509 15844 9512
rect 15013 9503 15071 9509
rect 15013 9500 15025 9503
rect 14884 9472 15025 9500
rect 14884 9460 14890 9472
rect 15013 9469 15025 9472
rect 15059 9469 15071 9503
rect 15832 9500 15844 9509
rect 15751 9472 15844 9500
rect 15013 9463 15071 9469
rect 15832 9463 15844 9472
rect 15896 9500 15902 9512
rect 16592 9500 16620 9676
rect 15896 9472 16620 9500
rect 15838 9460 15844 9463
rect 15896 9460 15902 9472
rect 16758 9460 16764 9512
rect 16816 9500 16822 9512
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 16816 9472 17233 9500
rect 16816 9460 16822 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17310 9460 17316 9512
rect 17368 9500 17374 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17368 9472 18061 9500
rect 17368 9460 17374 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 9306 9392 9312 9444
rect 9364 9441 9370 9444
rect 9364 9435 9428 9441
rect 9364 9401 9382 9435
rect 9416 9401 9428 9435
rect 10594 9432 10600 9444
rect 9364 9395 9428 9401
rect 9499 9404 10600 9432
rect 9364 9392 9370 9395
rect 9499 9364 9527 9404
rect 10594 9392 10600 9404
rect 10652 9392 10658 9444
rect 10686 9392 10692 9444
rect 10744 9432 10750 9444
rect 12710 9432 12716 9444
rect 10744 9404 12716 9432
rect 10744 9392 10750 9404
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 14461 9435 14519 9441
rect 14461 9432 14473 9435
rect 13004 9404 14473 9432
rect 9140 9336 9527 9364
rect 7009 9327 7067 9333
rect 9582 9324 9588 9376
rect 9640 9364 9646 9376
rect 10318 9364 10324 9376
rect 9640 9336 10324 9364
rect 9640 9324 9646 9336
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10505 9367 10563 9373
rect 10505 9333 10517 9367
rect 10551 9364 10563 9367
rect 10778 9364 10784 9376
rect 10551 9336 10784 9364
rect 10551 9333 10563 9336
rect 10505 9327 10563 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 13004 9373 13032 9404
rect 14461 9401 14473 9404
rect 14507 9401 14519 9435
rect 17494 9432 17500 9444
rect 17455 9404 17500 9432
rect 14461 9395 14519 9401
rect 17494 9392 17500 9404
rect 17552 9392 17558 9444
rect 12989 9367 13047 9373
rect 11848 9336 11893 9364
rect 11848 9324 11854 9336
rect 12989 9333 13001 9367
rect 13035 9333 13047 9367
rect 12989 9327 13047 9333
rect 13170 9324 13176 9376
rect 13228 9364 13234 9376
rect 13357 9367 13415 9373
rect 13357 9364 13369 9367
rect 13228 9336 13369 9364
rect 13228 9324 13234 9336
rect 13357 9333 13369 9336
rect 13403 9333 13415 9367
rect 13357 9327 13415 9333
rect 13449 9367 13507 9373
rect 13449 9333 13461 9367
rect 13495 9364 13507 9367
rect 13538 9364 13544 9376
rect 13495 9336 13544 9364
rect 13495 9333 13507 9336
rect 13449 9327 13507 9333
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 14366 9364 14372 9376
rect 14327 9336 14372 9364
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 16390 9364 16396 9376
rect 15243 9336 16396 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 16945 9367 17003 9373
rect 16945 9333 16957 9367
rect 16991 9364 17003 9367
rect 17218 9364 17224 9376
rect 16991 9336 17224 9364
rect 16991 9333 17003 9336
rect 16945 9327 17003 9333
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 17862 9324 17868 9376
rect 17920 9364 17926 9376
rect 18233 9367 18291 9373
rect 18233 9364 18245 9367
rect 17920 9336 18245 9364
rect 17920 9324 17926 9336
rect 18233 9333 18245 9336
rect 18279 9333 18291 9367
rect 18233 9327 18291 9333
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 4614 9160 4620 9172
rect 2188 9132 4620 9160
rect 2188 9120 2194 9132
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 5442 9160 5448 9172
rect 5403 9132 5448 9160
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 5721 9163 5779 9169
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 7282 9160 7288 9172
rect 5767 9132 7288 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7926 9160 7932 9172
rect 7887 9132 7932 9160
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 8018 9120 8024 9172
rect 8076 9160 8082 9172
rect 8076 9132 8524 9160
rect 8076 9120 8082 9132
rect 1664 9095 1722 9101
rect 1664 9061 1676 9095
rect 1710 9092 1722 9095
rect 3326 9092 3332 9104
rect 1710 9064 3332 9092
rect 1710 9061 1722 9064
rect 1664 9055 1722 9061
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 4430 9052 4436 9104
rect 4488 9092 4494 9104
rect 8389 9095 8447 9101
rect 8389 9092 8401 9095
rect 4488 9064 8401 9092
rect 4488 9052 4494 9064
rect 8389 9061 8401 9064
rect 8435 9061 8447 9095
rect 8389 9055 8447 9061
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1946 9024 1952 9036
rect 1443 8996 1952 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 1946 8984 1952 8996
rect 2004 9024 2010 9036
rect 2004 8996 2452 9024
rect 2004 8984 2010 8996
rect 2424 8968 2452 8996
rect 2682 8984 2688 9036
rect 2740 9024 2746 9036
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2740 8996 2881 9024
rect 2740 8984 2746 8996
rect 2869 8993 2881 8996
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 3053 9027 3111 9033
rect 3053 9024 3065 9027
rect 3016 8996 3065 9024
rect 3016 8984 3022 8996
rect 3053 8993 3065 8996
rect 3099 9024 3111 9027
rect 3694 9024 3700 9036
rect 3099 8996 3700 9024
rect 3099 8993 3111 8996
rect 3053 8987 3111 8993
rect 3694 8984 3700 8996
rect 3752 8984 3758 9036
rect 4338 9033 4344 9036
rect 4332 9024 4344 9033
rect 4251 8996 4344 9024
rect 4332 8987 4344 8996
rect 4396 9024 4402 9036
rect 6270 9024 6276 9036
rect 4396 8996 5304 9024
rect 6231 8996 6276 9024
rect 4338 8984 4344 8987
rect 4396 8984 4402 8996
rect 2406 8916 2412 8968
rect 2464 8956 2470 8968
rect 3786 8956 3792 8968
rect 2464 8928 3792 8956
rect 2464 8916 2470 8928
rect 3786 8916 3792 8928
rect 3844 8956 3850 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3844 8928 4077 8956
rect 3844 8916 3850 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 3237 8891 3295 8897
rect 3237 8888 3249 8891
rect 2332 8860 3249 8888
rect 1118 8780 1124 8832
rect 1176 8820 1182 8832
rect 2332 8820 2360 8860
rect 3237 8857 3249 8860
rect 3283 8857 3295 8891
rect 3237 8851 3295 8857
rect 1176 8792 2360 8820
rect 2777 8823 2835 8829
rect 1176 8780 1182 8792
rect 2777 8789 2789 8823
rect 2823 8820 2835 8823
rect 2869 8823 2927 8829
rect 2869 8820 2881 8823
rect 2823 8792 2881 8820
rect 2823 8789 2835 8792
rect 2777 8783 2835 8789
rect 2869 8789 2881 8792
rect 2915 8789 2927 8823
rect 4080 8820 4108 8919
rect 5074 8820 5080 8832
rect 4080 8792 5080 8820
rect 2869 8783 2927 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5276 8820 5304 8996
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 6540 9027 6598 9033
rect 6540 8993 6552 9027
rect 6586 9024 6598 9027
rect 7558 9024 7564 9036
rect 6586 8996 7564 9024
rect 6586 8993 6598 8996
rect 6540 8987 6598 8993
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 8294 9024 8300 9036
rect 8255 8996 8300 9024
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 8496 9024 8524 9132
rect 8938 9120 8944 9172
rect 8996 9160 9002 9172
rect 9122 9160 9128 9172
rect 8996 9132 9128 9160
rect 8996 9120 9002 9132
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10137 9163 10195 9169
rect 10137 9129 10149 9163
rect 10183 9160 10195 9163
rect 10870 9160 10876 9172
rect 10183 9132 10876 9160
rect 10183 9129 10195 9132
rect 10137 9123 10195 9129
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 11425 9163 11483 9169
rect 11425 9129 11437 9163
rect 11471 9160 11483 9163
rect 11790 9160 11796 9172
rect 11471 9132 11796 9160
rect 11471 9129 11483 9132
rect 11425 9123 11483 9129
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 12437 9163 12495 9169
rect 12437 9129 12449 9163
rect 12483 9160 12495 9163
rect 14366 9160 14372 9172
rect 12483 9132 14372 9160
rect 12483 9129 12495 9132
rect 12437 9123 12495 9129
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 14550 9120 14556 9172
rect 14608 9160 14614 9172
rect 14829 9163 14887 9169
rect 14829 9160 14841 9163
rect 14608 9132 14841 9160
rect 14608 9120 14614 9132
rect 14829 9129 14841 9132
rect 14875 9129 14887 9163
rect 14829 9123 14887 9129
rect 14918 9120 14924 9172
rect 14976 9160 14982 9172
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 14976 9132 15761 9160
rect 14976 9120 14982 9132
rect 15749 9129 15761 9132
rect 15795 9129 15807 9163
rect 15749 9123 15807 9129
rect 15841 9163 15899 9169
rect 15841 9129 15853 9163
rect 15887 9160 15899 9163
rect 16298 9160 16304 9172
rect 15887 9132 16304 9160
rect 15887 9129 15899 9132
rect 15841 9123 15899 9129
rect 16298 9120 16304 9132
rect 16356 9120 16362 9172
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 9493 9095 9551 9101
rect 9493 9092 9505 9095
rect 8628 9064 9505 9092
rect 8628 9052 8634 9064
rect 9493 9061 9505 9064
rect 9539 9061 9551 9095
rect 9493 9055 9551 9061
rect 9582 9052 9588 9104
rect 9640 9092 9646 9104
rect 10045 9095 10103 9101
rect 10045 9092 10057 9095
rect 9640 9064 10057 9092
rect 9640 9052 9646 9064
rect 10045 9061 10057 9064
rect 10091 9061 10103 9095
rect 10045 9055 10103 9061
rect 10965 9095 11023 9101
rect 10965 9061 10977 9095
rect 11011 9092 11023 9095
rect 12342 9092 12348 9104
rect 11011 9064 12348 9092
rect 11011 9061 11023 9064
rect 10965 9055 11023 9061
rect 12342 9052 12348 9064
rect 12400 9052 12406 9104
rect 12897 9095 12955 9101
rect 12897 9061 12909 9095
rect 12943 9092 12955 9095
rect 13262 9092 13268 9104
rect 12943 9064 13268 9092
rect 12943 9061 12955 9064
rect 12897 9055 12955 9061
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 8496 8996 10701 9024
rect 10689 8993 10701 8996
rect 10735 8993 10747 9027
rect 10689 8987 10747 8993
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 9024 11851 9027
rect 12526 9024 12532 9036
rect 11839 8996 12532 9024
rect 11839 8993 11851 8996
rect 11793 8987 11851 8993
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 12618 8984 12624 9036
rect 12676 9024 12682 9036
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 12676 8996 12817 9024
rect 12676 8984 12682 8996
rect 12805 8993 12817 8996
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 8662 8956 8668 8968
rect 8619 8928 8668 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8662 8916 8668 8928
rect 8720 8956 8726 8968
rect 8846 8956 8852 8968
rect 8720 8928 8852 8956
rect 8720 8916 8726 8928
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 8938 8916 8944 8968
rect 8996 8956 9002 8968
rect 10042 8956 10048 8968
rect 8996 8928 10048 8956
rect 8996 8916 9002 8928
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 9493 8891 9551 8897
rect 7208 8860 8248 8888
rect 7208 8820 7236 8860
rect 5276 8792 7236 8820
rect 7653 8823 7711 8829
rect 7653 8789 7665 8823
rect 7699 8820 7711 8823
rect 8110 8820 8116 8832
rect 7699 8792 8116 8820
rect 7699 8789 7711 8792
rect 7653 8783 7711 8789
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 8220 8820 8248 8860
rect 9493 8857 9505 8891
rect 9539 8888 9551 8891
rect 10134 8888 10140 8900
rect 9539 8860 10140 8888
rect 9539 8857 9551 8860
rect 9493 8851 9551 8857
rect 10134 8848 10140 8860
rect 10192 8848 10198 8900
rect 10244 8820 10272 8919
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 11112 8928 11897 8956
rect 11112 8916 11118 8928
rect 11885 8925 11897 8928
rect 11931 8956 11943 8959
rect 11974 8956 11980 8968
rect 11931 8928 11980 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 12069 8959 12127 8965
rect 12069 8925 12081 8959
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 12084 8888 12112 8919
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 12434 8956 12440 8968
rect 12216 8928 12440 8956
rect 12216 8916 12222 8928
rect 12434 8916 12440 8928
rect 12492 8956 12498 8968
rect 12912 8956 12940 9055
rect 13262 9052 13268 9064
rect 13320 9052 13326 9104
rect 16684 9092 16712 9120
rect 16684 9064 18092 9092
rect 18064 9036 18092 9064
rect 13722 9033 13728 9036
rect 13716 9024 13728 9033
rect 13096 8996 13728 9024
rect 13096 8965 13124 8996
rect 13716 8987 13728 8996
rect 13722 8984 13728 8987
rect 13780 8984 13786 9036
rect 15102 8984 15108 9036
rect 15160 9024 15166 9036
rect 16393 9027 16451 9033
rect 16393 9024 16405 9027
rect 15160 8996 16405 9024
rect 15160 8984 15166 8996
rect 16393 8993 16405 8996
rect 16439 8993 16451 9027
rect 16393 8987 16451 8993
rect 16660 9027 16718 9033
rect 16660 8993 16672 9027
rect 16706 9024 16718 9027
rect 17218 9024 17224 9036
rect 16706 8996 17224 9024
rect 16706 8993 16718 8996
rect 16660 8987 16718 8993
rect 17218 8984 17224 8996
rect 17276 8984 17282 9036
rect 18046 9024 18052 9036
rect 17959 8996 18052 9024
rect 18046 8984 18052 8996
rect 18104 8984 18110 9036
rect 12492 8928 12940 8956
rect 13081 8959 13139 8965
rect 12492 8916 12498 8928
rect 13081 8925 13093 8959
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 13096 8888 13124 8919
rect 12084 8860 13124 8888
rect 8220 8792 10272 8820
rect 10686 8780 10692 8832
rect 10744 8820 10750 8832
rect 12342 8820 12348 8832
rect 10744 8792 12348 8820
rect 10744 8780 10750 8792
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 13464 8820 13492 8919
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 15933 8959 15991 8965
rect 15933 8956 15945 8959
rect 15896 8928 15945 8956
rect 15896 8916 15902 8928
rect 15933 8925 15945 8928
rect 15979 8925 15991 8959
rect 15933 8919 15991 8925
rect 15102 8888 15108 8900
rect 14384 8860 15108 8888
rect 14384 8820 14412 8860
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 13464 8792 14412 8820
rect 15010 8780 15016 8832
rect 15068 8820 15074 8832
rect 15381 8823 15439 8829
rect 15381 8820 15393 8823
rect 15068 8792 15393 8820
rect 15068 8780 15074 8792
rect 15381 8789 15393 8792
rect 15427 8789 15439 8823
rect 15381 8783 15439 8789
rect 16758 8780 16764 8832
rect 16816 8820 16822 8832
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 16816 8792 17785 8820
rect 16816 8780 16822 8792
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 17773 8783 17831 8789
rect 18233 8823 18291 8829
rect 18233 8789 18245 8823
rect 18279 8820 18291 8823
rect 18322 8820 18328 8832
rect 18279 8792 18328 8820
rect 18279 8789 18291 8792
rect 18233 8783 18291 8789
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 3234 8576 3240 8628
rect 3292 8576 3298 8628
rect 3973 8619 4031 8625
rect 3973 8585 3985 8619
rect 4019 8616 4031 8619
rect 8294 8616 8300 8628
rect 4019 8588 8300 8616
rect 4019 8585 4031 8588
rect 3973 8579 4031 8585
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 9088 8588 9229 8616
rect 9088 8576 9094 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 11054 8616 11060 8628
rect 9217 8579 9275 8585
rect 10060 8588 11060 8616
rect 1857 8551 1915 8557
rect 1857 8517 1869 8551
rect 1903 8517 1915 8551
rect 3252 8548 3280 8576
rect 3697 8551 3755 8557
rect 3697 8548 3709 8551
rect 3252 8520 3709 8548
rect 1857 8511 1915 8517
rect 3697 8517 3709 8520
rect 3743 8548 3755 8551
rect 4338 8548 4344 8560
rect 3743 8520 4344 8548
rect 3743 8517 3755 8520
rect 3697 8511 3755 8517
rect 1872 8480 1900 8511
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 4985 8551 5043 8557
rect 4985 8517 4997 8551
rect 5031 8548 5043 8551
rect 6730 8548 6736 8560
rect 5031 8520 6736 8548
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 8570 8508 8576 8560
rect 8628 8548 8634 8560
rect 10060 8548 10088 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 12158 8616 12164 8628
rect 11164 8588 12164 8616
rect 8628 8520 10088 8548
rect 8628 8508 8634 8520
rect 1872 8452 2452 8480
rect 1670 8412 1676 8424
rect 1631 8384 1676 8412
rect 1670 8372 1676 8384
rect 1728 8372 1734 8424
rect 2314 8412 2320 8424
rect 2275 8384 2320 8412
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 2424 8412 2452 8452
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 3384 8452 4537 8480
rect 3384 8440 3390 8452
rect 4525 8449 4537 8452
rect 4571 8480 4583 8483
rect 4614 8480 4620 8492
rect 4571 8452 4620 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4614 8440 4620 8452
rect 4672 8480 4678 8492
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 4672 8452 5549 8480
rect 4672 8440 4678 8452
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 6638 8480 6644 8492
rect 6328 8452 6644 8480
rect 6328 8440 6334 8452
rect 6638 8440 6644 8452
rect 6696 8480 6702 8492
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 6696 8452 7573 8480
rect 6696 8440 6702 8452
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 9306 8480 9312 8492
rect 8996 8452 9312 8480
rect 8996 8440 9002 8452
rect 9306 8440 9312 8452
rect 9364 8480 9370 8492
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9364 8452 9781 8480
rect 9364 8440 9370 8452
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 5994 8412 6000 8424
rect 2424 8384 3280 8412
rect 5955 8384 6000 8412
rect 3252 8356 3280 8384
rect 5994 8372 6000 8384
rect 6052 8372 6058 8424
rect 8662 8412 8668 8424
rect 7760 8384 8668 8412
rect 2590 8353 2596 8356
rect 2584 8344 2596 8353
rect 2551 8316 2596 8344
rect 2584 8307 2596 8316
rect 2590 8304 2596 8307
rect 2648 8304 2654 8356
rect 3234 8304 3240 8356
rect 3292 8304 3298 8356
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 5445 8347 5503 8353
rect 5445 8344 5457 8347
rect 4304 8316 5457 8344
rect 4304 8304 4310 8316
rect 5445 8313 5457 8316
rect 5491 8344 5503 8347
rect 6454 8344 6460 8356
rect 5491 8316 6460 8344
rect 5491 8313 5503 8316
rect 5445 8307 5503 8313
rect 6454 8304 6460 8316
rect 6512 8304 6518 8356
rect 7101 8347 7159 8353
rect 7101 8313 7113 8347
rect 7147 8344 7159 8347
rect 7760 8344 7788 8384
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 9030 8372 9036 8424
rect 9088 8412 9094 8424
rect 9585 8415 9643 8421
rect 9585 8412 9597 8415
rect 9088 8384 9597 8412
rect 9088 8372 9094 8384
rect 9585 8381 9597 8384
rect 9631 8412 9643 8415
rect 10042 8412 10048 8424
rect 9631 8384 9812 8412
rect 10003 8384 10048 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 7147 8316 7788 8344
rect 7828 8347 7886 8353
rect 7147 8313 7159 8316
rect 7101 8307 7159 8313
rect 7828 8313 7840 8347
rect 7874 8344 7886 8347
rect 8110 8344 8116 8356
rect 7874 8316 8116 8344
rect 7874 8313 7886 8316
rect 7828 8307 7886 8313
rect 8110 8304 8116 8316
rect 8168 8304 8174 8356
rect 8570 8304 8576 8356
rect 8628 8344 8634 8356
rect 9677 8347 9735 8353
rect 9677 8344 9689 8347
rect 8628 8316 9689 8344
rect 8628 8304 8634 8316
rect 9677 8313 9689 8316
rect 9723 8313 9735 8347
rect 9677 8307 9735 8313
rect 2406 8236 2412 8288
rect 2464 8276 2470 8288
rect 2958 8276 2964 8288
rect 2464 8248 2964 8276
rect 2464 8236 2470 8248
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 3602 8276 3608 8288
rect 3108 8248 3608 8276
rect 3108 8236 3114 8248
rect 3602 8236 3608 8248
rect 3660 8236 3666 8288
rect 4338 8276 4344 8288
rect 4299 8248 4344 8276
rect 4338 8236 4344 8248
rect 4396 8236 4402 8288
rect 4433 8279 4491 8285
rect 4433 8245 4445 8279
rect 4479 8276 4491 8279
rect 4522 8276 4528 8288
rect 4479 8248 4528 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4522 8236 4528 8248
rect 4580 8276 4586 8288
rect 5258 8276 5264 8288
rect 4580 8248 5264 8276
rect 4580 8236 4586 8248
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 6178 8276 6184 8288
rect 5408 8248 5453 8276
rect 6139 8248 6184 8276
rect 5408 8236 5414 8248
rect 6178 8236 6184 8248
rect 6236 8236 6242 8288
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 8938 8276 8944 8288
rect 6604 8248 8944 8276
rect 6604 8236 6610 8248
rect 8938 8236 8944 8248
rect 8996 8236 9002 8288
rect 9784 8276 9812 8384
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10312 8415 10370 8421
rect 10312 8381 10324 8415
rect 10358 8412 10370 8415
rect 10870 8412 10876 8424
rect 10358 8384 10876 8412
rect 10358 8381 10370 8384
rect 10312 8375 10370 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11164 8412 11192 8588
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 12342 8576 12348 8628
rect 12400 8616 12406 8628
rect 12400 8588 18092 8616
rect 12400 8576 12406 8588
rect 11330 8508 11336 8560
rect 11388 8548 11394 8560
rect 11425 8551 11483 8557
rect 11425 8548 11437 8551
rect 11388 8520 11437 8548
rect 11388 8508 11394 8520
rect 11425 8517 11437 8520
rect 11471 8517 11483 8551
rect 11425 8511 11483 8517
rect 11517 8551 11575 8557
rect 11517 8517 11529 8551
rect 11563 8517 11575 8551
rect 13541 8551 13599 8557
rect 13541 8548 13553 8551
rect 11517 8511 11575 8517
rect 11900 8520 13553 8548
rect 11072 8384 11192 8412
rect 9858 8304 9864 8356
rect 9916 8344 9922 8356
rect 10686 8344 10692 8356
rect 9916 8316 10692 8344
rect 9916 8304 9922 8316
rect 10686 8304 10692 8316
rect 10744 8344 10750 8356
rect 10962 8344 10968 8356
rect 10744 8316 10968 8344
rect 10744 8304 10750 8316
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 11072 8276 11100 8384
rect 11532 8344 11560 8511
rect 11900 8421 11928 8520
rect 13541 8517 13553 8520
rect 13587 8517 13599 8551
rect 13541 8511 13599 8517
rect 13906 8508 13912 8560
rect 13964 8548 13970 8560
rect 14182 8548 14188 8560
rect 13964 8520 14188 8548
rect 13964 8508 13970 8520
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 12066 8480 12072 8492
rect 12027 8452 12072 8480
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 12216 8452 12848 8480
rect 12216 8440 12222 8452
rect 11885 8415 11943 8421
rect 11885 8381 11897 8415
rect 11931 8381 11943 8415
rect 11885 8375 11943 8381
rect 11977 8415 12035 8421
rect 11977 8381 11989 8415
rect 12023 8412 12035 8415
rect 12710 8412 12716 8424
rect 12023 8384 12716 8412
rect 12023 8381 12035 8384
rect 11977 8375 12035 8381
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 12820 8421 12848 8452
rect 12894 8440 12900 8492
rect 12952 8440 12958 8492
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8480 13139 8483
rect 13262 8480 13268 8492
rect 13127 8452 13268 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 13446 8440 13452 8492
rect 13504 8480 13510 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13504 8452 14105 8480
rect 13504 8440 13510 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8480 14611 8483
rect 17218 8480 17224 8492
rect 14599 8452 15148 8480
rect 17179 8452 17224 8480
rect 14599 8449 14611 8452
rect 14553 8443 14611 8449
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8381 12863 8415
rect 12912 8412 12940 8440
rect 13909 8415 13967 8421
rect 13909 8412 13921 8415
rect 12912 8384 13921 8412
rect 12805 8375 12863 8381
rect 13909 8381 13921 8384
rect 13955 8412 13967 8415
rect 14366 8412 14372 8424
rect 13955 8384 14372 8412
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 15013 8415 15071 8421
rect 15013 8381 15025 8415
rect 15059 8381 15071 8415
rect 15120 8412 15148 8452
rect 17218 8440 17224 8452
rect 17276 8440 17282 8492
rect 15654 8412 15660 8424
rect 15120 8384 15660 8412
rect 15013 8375 15071 8381
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 11532 8316 12909 8344
rect 12897 8313 12909 8316
rect 12943 8313 12955 8347
rect 12897 8307 12955 8313
rect 14001 8347 14059 8353
rect 14001 8313 14013 8347
rect 14047 8344 14059 8347
rect 14918 8344 14924 8356
rect 14047 8316 14924 8344
rect 14047 8313 14059 8316
rect 14001 8307 14059 8313
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 15028 8344 15056 8375
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 17037 8415 17095 8421
rect 17037 8412 17049 8415
rect 16540 8384 17049 8412
rect 16540 8372 16546 8384
rect 17037 8381 17049 8384
rect 17083 8381 17095 8415
rect 17037 8375 17095 8381
rect 17126 8372 17132 8424
rect 17184 8412 17190 8424
rect 18064 8421 18092 8588
rect 18230 8548 18236 8560
rect 18191 8520 18236 8548
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 18049 8415 18107 8421
rect 17184 8384 17229 8412
rect 17184 8372 17190 8384
rect 18049 8381 18061 8415
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 15102 8344 15108 8356
rect 15028 8316 15108 8344
rect 15102 8304 15108 8316
rect 15160 8304 15166 8356
rect 15280 8347 15338 8353
rect 15280 8313 15292 8347
rect 15326 8344 15338 8347
rect 16758 8344 16764 8356
rect 15326 8316 16764 8344
rect 15326 8313 15338 8316
rect 15280 8307 15338 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 17218 8304 17224 8356
rect 17276 8344 17282 8356
rect 17678 8344 17684 8356
rect 17276 8316 17684 8344
rect 17276 8304 17282 8316
rect 17678 8304 17684 8316
rect 17736 8304 17742 8356
rect 9784 8248 11100 8276
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11882 8276 11888 8288
rect 11204 8248 11888 8276
rect 11204 8236 11210 8248
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 12492 8248 12537 8276
rect 12492 8236 12498 8248
rect 12618 8236 12624 8288
rect 12676 8276 12682 8288
rect 16206 8276 16212 8288
rect 12676 8248 16212 8276
rect 12676 8236 12682 8248
rect 16206 8236 16212 8248
rect 16264 8236 16270 8288
rect 16298 8236 16304 8288
rect 16356 8276 16362 8288
rect 16393 8279 16451 8285
rect 16393 8276 16405 8279
rect 16356 8248 16405 8276
rect 16356 8236 16362 8248
rect 16393 8245 16405 8248
rect 16439 8245 16451 8279
rect 16666 8276 16672 8288
rect 16627 8248 16672 8276
rect 16393 8239 16451 8245
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 2317 8075 2375 8081
rect 2317 8041 2329 8075
rect 2363 8072 2375 8075
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2363 8044 2973 8072
rect 2363 8041 2375 8044
rect 2317 8035 2375 8041
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 3510 8072 3516 8084
rect 3467 8044 3516 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8072 4123 8075
rect 4430 8072 4436 8084
rect 4111 8044 4436 8072
rect 4111 8041 4123 8044
rect 4065 8035 4123 8041
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 7650 8072 7656 8084
rect 5276 8044 7656 8072
rect 5276 8004 5304 8044
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 8386 8072 8392 8084
rect 8347 8044 8392 8072
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8478 8032 8484 8084
rect 8536 8072 8542 8084
rect 8757 8075 8815 8081
rect 8757 8072 8769 8075
rect 8536 8044 8769 8072
rect 8536 8032 8542 8044
rect 8757 8041 8769 8044
rect 8803 8072 8815 8075
rect 9858 8072 9864 8084
rect 8803 8044 9864 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 10321 8075 10379 8081
rect 10321 8041 10333 8075
rect 10367 8072 10379 8075
rect 12158 8072 12164 8084
rect 10367 8044 12164 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 12618 8072 12624 8084
rect 12400 8044 12624 8072
rect 12400 8032 12406 8044
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12759 8044 12909 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 12897 8035 12955 8041
rect 13722 8032 13728 8084
rect 13780 8072 13786 8084
rect 14369 8075 14427 8081
rect 14369 8072 14381 8075
rect 13780 8044 14381 8072
rect 13780 8032 13786 8044
rect 14369 8041 14381 8044
rect 14415 8041 14427 8075
rect 14369 8035 14427 8041
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 17405 8075 17463 8081
rect 17405 8072 17417 8075
rect 16264 8044 17417 8072
rect 16264 8032 16270 8044
rect 17405 8041 17417 8044
rect 17451 8072 17463 8075
rect 17954 8072 17960 8084
rect 17451 8044 17960 8072
rect 17451 8041 17463 8044
rect 17405 8035 17463 8041
rect 17954 8032 17960 8044
rect 18012 8032 18018 8084
rect 1412 7976 5304 8004
rect 5344 8007 5402 8013
rect 1412 7945 1440 7976
rect 5344 7973 5356 8007
rect 5390 8004 5402 8007
rect 6546 8004 6552 8016
rect 5390 7976 6552 8004
rect 5390 7973 5402 7976
rect 5344 7967 5402 7973
rect 6546 7964 6552 7976
rect 6604 7964 6610 8016
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 8849 8007 8907 8013
rect 8849 8004 8861 8007
rect 6788 7976 8861 8004
rect 6788 7964 6794 7976
rect 8849 7973 8861 7976
rect 8895 7973 8907 8007
rect 11882 8004 11888 8016
rect 8849 7967 8907 7973
rect 9692 7976 11888 8004
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 1397 7899 1455 7905
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7905 3387 7939
rect 3329 7899 3387 7905
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 5074 7936 5080 7948
rect 4479 7908 4936 7936
rect 5035 7908 5080 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7868 2467 7871
rect 2498 7868 2504 7880
rect 2455 7840 2504 7868
rect 2455 7837 2467 7840
rect 2409 7831 2467 7837
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 3050 7868 3056 7880
rect 2639 7840 3056 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 1581 7803 1639 7809
rect 1581 7769 1593 7803
rect 1627 7800 1639 7803
rect 1627 7772 2268 7800
rect 1627 7769 1639 7772
rect 1581 7763 1639 7769
rect 1946 7732 1952 7744
rect 1907 7704 1952 7732
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 2240 7732 2268 7772
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 3344 7800 3372 7899
rect 3513 7871 3571 7877
rect 3513 7837 3525 7871
rect 3559 7837 3571 7871
rect 3513 7831 3571 7837
rect 2372 7772 3372 7800
rect 2372 7760 2378 7772
rect 3418 7760 3424 7812
rect 3476 7800 3482 7812
rect 3528 7800 3556 7831
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 3844 7840 4537 7868
rect 3844 7828 3850 7840
rect 4525 7837 4537 7840
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4614 7828 4620 7880
rect 4672 7868 4678 7880
rect 4672 7840 4717 7868
rect 4672 7828 4678 7840
rect 3476 7772 3556 7800
rect 3476 7760 3482 7772
rect 3510 7732 3516 7744
rect 2240 7704 3516 7732
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 4908 7732 4936 7908
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 7000 7939 7058 7945
rect 7000 7936 7012 7939
rect 6472 7908 7012 7936
rect 6472 7809 6500 7908
rect 7000 7905 7012 7908
rect 7046 7936 7058 7939
rect 7374 7936 7380 7948
rect 7046 7908 7380 7936
rect 7046 7905 7058 7908
rect 7000 7899 7058 7905
rect 7374 7896 7380 7908
rect 7432 7936 7438 7948
rect 8018 7936 8024 7948
rect 7432 7908 8024 7936
rect 7432 7896 7438 7908
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 9692 7945 9720 7976
rect 11882 7964 11888 7976
rect 11940 7964 11946 8016
rect 12250 7964 12256 8016
rect 12308 8004 12314 8016
rect 12308 7976 18000 8004
rect 12308 7964 12314 7976
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7905 9735 7939
rect 10686 7936 10692 7948
rect 10647 7908 10692 7936
rect 9677 7899 9735 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 11600 7939 11658 7945
rect 11600 7936 11612 7939
rect 10980 7908 11612 7936
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6696 7840 6745 7868
rect 6696 7828 6702 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8904 7840 8953 7868
rect 8904 7828 8910 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9398 7828 9404 7880
rect 9456 7868 9462 7880
rect 9861 7871 9919 7877
rect 9861 7868 9873 7871
rect 9456 7840 9873 7868
rect 9456 7828 9462 7840
rect 9861 7837 9873 7840
rect 9907 7837 9919 7871
rect 10778 7868 10784 7880
rect 10739 7840 10784 7868
rect 9861 7831 9919 7837
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 10980 7877 11008 7908
rect 11600 7905 11612 7908
rect 11646 7936 11658 7939
rect 12066 7936 12072 7948
rect 11646 7908 12072 7936
rect 11646 7905 11658 7908
rect 11600 7899 11658 7905
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 13262 7945 13268 7948
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7936 12955 7939
rect 13245 7939 13268 7945
rect 13245 7936 13257 7939
rect 12943 7908 13257 7936
rect 12943 7905 12955 7908
rect 12897 7899 12955 7905
rect 13245 7905 13257 7908
rect 13320 7936 13326 7948
rect 13320 7908 13393 7936
rect 13245 7899 13268 7905
rect 13262 7896 13268 7899
rect 13320 7896 13326 7908
rect 14366 7896 14372 7948
rect 14424 7936 14430 7948
rect 14645 7939 14703 7945
rect 14645 7936 14657 7939
rect 14424 7908 14657 7936
rect 14424 7896 14430 7908
rect 14645 7905 14657 7908
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 15556 7939 15614 7945
rect 15556 7905 15568 7939
rect 15602 7936 15614 7939
rect 16298 7936 16304 7948
rect 15602 7908 16304 7936
rect 15602 7905 15614 7908
rect 15556 7899 15614 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 17310 7936 17316 7948
rect 16408 7908 17316 7936
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 12996 7871 13054 7877
rect 12996 7837 13008 7871
rect 13042 7837 13054 7871
rect 12996 7831 13054 7837
rect 6457 7803 6515 7809
rect 6457 7769 6469 7803
rect 6503 7769 6515 7803
rect 8386 7800 8392 7812
rect 6457 7763 6515 7769
rect 7668 7772 8392 7800
rect 7668 7732 7696 7772
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 10594 7800 10600 7812
rect 10100 7772 10600 7800
rect 10100 7760 10106 7772
rect 10594 7760 10600 7772
rect 10652 7800 10658 7812
rect 11348 7800 11376 7831
rect 13004 7800 13032 7831
rect 15102 7828 15108 7880
rect 15160 7868 15166 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15160 7840 15301 7868
rect 15160 7828 15166 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 10652 7772 11376 7800
rect 10652 7760 10658 7772
rect 4908 7704 7696 7732
rect 7742 7692 7748 7744
rect 7800 7732 7806 7744
rect 8113 7735 8171 7741
rect 8113 7732 8125 7735
rect 7800 7704 8125 7732
rect 7800 7692 7806 7704
rect 8113 7701 8125 7704
rect 8159 7701 8171 7735
rect 11348 7732 11376 7772
rect 12544 7772 13032 7800
rect 12544 7732 12572 7772
rect 11348 7704 12572 7732
rect 8113 7695 8171 7701
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 14550 7732 14556 7744
rect 13412 7704 14556 7732
rect 13412 7692 13418 7704
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 14829 7735 14887 7741
rect 14829 7701 14841 7735
rect 14875 7732 14887 7735
rect 15194 7732 15200 7744
rect 14875 7704 15200 7732
rect 14875 7701 14887 7704
rect 14829 7695 14887 7701
rect 15194 7692 15200 7704
rect 15252 7692 15258 7744
rect 15562 7692 15568 7744
rect 15620 7732 15626 7744
rect 16408 7732 16436 7908
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 17972 7945 18000 7976
rect 17957 7939 18015 7945
rect 17957 7905 17969 7939
rect 18003 7905 18015 7939
rect 17957 7899 18015 7905
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 16758 7760 16764 7812
rect 16816 7800 16822 7812
rect 17512 7800 17540 7831
rect 17678 7800 17684 7812
rect 16816 7772 17684 7800
rect 16816 7760 16822 7772
rect 17678 7760 17684 7772
rect 17736 7760 17742 7812
rect 15620 7704 16436 7732
rect 15620 7692 15626 7704
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 16669 7735 16727 7741
rect 16669 7732 16681 7735
rect 16632 7704 16681 7732
rect 16632 7692 16638 7704
rect 16669 7701 16681 7704
rect 16715 7701 16727 7735
rect 16942 7732 16948 7744
rect 16903 7704 16948 7732
rect 16669 7695 16727 7701
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 17770 7692 17776 7744
rect 17828 7732 17834 7744
rect 18141 7735 18199 7741
rect 18141 7732 18153 7735
rect 17828 7704 18153 7732
rect 17828 7692 17834 7704
rect 18141 7701 18153 7704
rect 18187 7701 18199 7735
rect 18141 7695 18199 7701
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 2498 7488 2504 7540
rect 2556 7528 2562 7540
rect 2869 7531 2927 7537
rect 2869 7528 2881 7531
rect 2556 7500 2881 7528
rect 2556 7488 2562 7500
rect 2869 7497 2881 7500
rect 2915 7497 2927 7531
rect 2869 7491 2927 7497
rect 3694 7488 3700 7540
rect 3752 7528 3758 7540
rect 4522 7528 4528 7540
rect 3752 7500 4528 7528
rect 3752 7488 3758 7500
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 4706 7488 4712 7540
rect 4764 7528 4770 7540
rect 5905 7531 5963 7537
rect 5905 7528 5917 7531
rect 4764 7500 5917 7528
rect 4764 7488 4770 7500
rect 5905 7497 5917 7500
rect 5951 7497 5963 7531
rect 5905 7491 5963 7497
rect 10229 7531 10287 7537
rect 10229 7497 10241 7531
rect 10275 7528 10287 7531
rect 10318 7528 10324 7540
rect 10275 7500 10324 7528
rect 10275 7497 10287 7500
rect 10229 7491 10287 7497
rect 10318 7488 10324 7500
rect 10376 7528 10382 7540
rect 10376 7500 11192 7528
rect 10376 7488 10382 7500
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 4338 7460 4344 7472
rect 1903 7432 4344 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 4338 7420 4344 7432
rect 4396 7420 4402 7472
rect 7834 7420 7840 7472
rect 7892 7420 7898 7472
rect 10594 7420 10600 7472
rect 10652 7460 10658 7472
rect 10962 7460 10968 7472
rect 10652 7432 10968 7460
rect 10652 7420 10658 7432
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 11164 7460 11192 7500
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11974 7528 11980 7540
rect 11296 7500 11980 7528
rect 11296 7488 11302 7500
rect 11974 7488 11980 7500
rect 12032 7528 12038 7540
rect 12621 7531 12679 7537
rect 12621 7528 12633 7531
rect 12032 7500 12633 7528
rect 12032 7488 12038 7500
rect 12621 7497 12633 7500
rect 12667 7497 12679 7531
rect 12621 7491 12679 7497
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 12897 7531 12955 7537
rect 12897 7528 12909 7531
rect 12768 7500 12909 7528
rect 12768 7488 12774 7500
rect 12897 7497 12909 7500
rect 12943 7497 12955 7531
rect 12897 7491 12955 7497
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 13504 7500 15301 7528
rect 13504 7488 13510 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 11333 7463 11391 7469
rect 11164 7432 11284 7460
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7392 1455 7395
rect 2314 7392 2320 7404
rect 1443 7364 2320 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 3050 7392 3056 7404
rect 2547 7364 3056 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 3418 7392 3424 7404
rect 3379 7364 3424 7392
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 6270 7392 6276 7404
rect 6104 7364 6276 7392
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7324 3755 7327
rect 3881 7327 3939 7333
rect 3881 7324 3893 7327
rect 3743 7296 3893 7324
rect 3743 7293 3755 7296
rect 3697 7287 3755 7293
rect 3881 7293 3893 7296
rect 3927 7324 3939 7327
rect 4522 7324 4528 7336
rect 3927 7296 4384 7324
rect 4483 7296 4528 7324
rect 3927 7293 3939 7296
rect 3881 7287 3939 7293
rect 2866 7216 2872 7268
rect 2924 7256 2930 7268
rect 4356 7256 4384 7296
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 4792 7327 4850 7333
rect 4792 7293 4804 7327
rect 4838 7324 4850 7327
rect 6104 7324 6132 7364
rect 6270 7352 6276 7364
rect 6328 7392 6334 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 6328 7364 7389 7392
rect 6328 7352 6334 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7852 7392 7880 7420
rect 8018 7392 8024 7404
rect 7377 7355 7435 7361
rect 7668 7364 8024 7392
rect 4838 7296 6132 7324
rect 6181 7327 6239 7333
rect 4838 7293 4850 7296
rect 4792 7287 4850 7293
rect 6181 7293 6193 7327
rect 6227 7324 6239 7327
rect 7668 7324 7696 7364
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 11146 7392 11152 7404
rect 8956 7364 11152 7392
rect 7834 7324 7840 7336
rect 6227 7296 7696 7324
rect 7795 7296 7840 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 8956 7333 8984 7364
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11256 7392 11284 7432
rect 11333 7429 11345 7463
rect 11379 7460 11391 7463
rect 12250 7460 12256 7472
rect 11379 7432 12256 7460
rect 11379 7429 11391 7432
rect 11333 7423 11391 7429
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 16390 7420 16396 7472
rect 16448 7460 16454 7472
rect 16448 7432 17080 7460
rect 16448 7420 16454 7432
rect 11977 7395 12035 7401
rect 11256 7364 11376 7392
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 11238 7324 11244 7336
rect 9180 7296 11244 7324
rect 9180 7284 9186 7296
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 11348 7324 11376 7364
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12526 7392 12532 7404
rect 12023 7364 12532 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12526 7352 12532 7364
rect 12584 7352 12590 7404
rect 13446 7392 13452 7404
rect 13407 7364 13452 7392
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7392 13783 7395
rect 13814 7392 13820 7404
rect 13771 7364 13820 7392
rect 13771 7361 13783 7364
rect 13725 7355 13783 7361
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 16577 7395 16635 7401
rect 16577 7361 16589 7395
rect 16623 7392 16635 7395
rect 16758 7392 16764 7404
rect 16623 7364 16764 7392
rect 16623 7361 16635 7364
rect 16577 7355 16635 7361
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 11348 7296 12817 7324
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 13909 7327 13967 7333
rect 13909 7293 13921 7327
rect 13955 7324 13967 7327
rect 15102 7324 15108 7336
rect 13955 7296 15108 7324
rect 13955 7293 13967 7296
rect 13909 7287 13967 7293
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 15194 7284 15200 7336
rect 15252 7324 15258 7336
rect 16114 7324 16120 7336
rect 15252 7296 16120 7324
rect 15252 7284 15258 7296
rect 16114 7284 16120 7296
rect 16172 7284 16178 7336
rect 16206 7284 16212 7336
rect 16264 7324 16270 7336
rect 16485 7327 16543 7333
rect 16264 7296 16344 7324
rect 16264 7284 16270 7296
rect 6730 7256 6736 7268
rect 2924 7228 4108 7256
rect 4356 7228 6736 7256
rect 2924 7216 2930 7228
rect 2222 7188 2228 7200
rect 2183 7160 2228 7188
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 2314 7148 2320 7200
rect 2372 7188 2378 7200
rect 2372 7160 2417 7188
rect 2372 7148 2378 7160
rect 2958 7148 2964 7200
rect 3016 7188 3022 7200
rect 4080 7197 4108 7228
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 7193 7259 7251 7265
rect 7193 7225 7205 7259
rect 7239 7256 7251 7259
rect 7558 7256 7564 7268
rect 7239 7228 7564 7256
rect 7239 7225 7251 7228
rect 7193 7219 7251 7225
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 7650 7216 7656 7268
rect 7708 7256 7714 7268
rect 8113 7259 8171 7265
rect 8113 7256 8125 7259
rect 7708 7228 8125 7256
rect 7708 7216 7714 7228
rect 8113 7225 8125 7228
rect 8159 7225 8171 7259
rect 8113 7219 8171 7225
rect 9030 7216 9036 7268
rect 9088 7256 9094 7268
rect 11054 7256 11060 7268
rect 9088 7228 11060 7256
rect 9088 7216 9094 7228
rect 11054 7216 11060 7228
rect 11112 7216 11118 7268
rect 11701 7259 11759 7265
rect 11701 7225 11713 7259
rect 11747 7256 11759 7259
rect 12710 7256 12716 7268
rect 11747 7228 12716 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 13265 7259 13323 7265
rect 13265 7225 13277 7259
rect 13311 7256 13323 7259
rect 13725 7259 13783 7265
rect 13725 7256 13737 7259
rect 13311 7228 13737 7256
rect 13311 7225 13323 7228
rect 13265 7219 13323 7225
rect 13725 7225 13737 7228
rect 13771 7225 13783 7259
rect 13725 7219 13783 7225
rect 14176 7259 14234 7265
rect 14176 7225 14188 7259
rect 14222 7256 14234 7259
rect 14458 7256 14464 7268
rect 14222 7228 14464 7256
rect 14222 7225 14234 7228
rect 14176 7219 14234 7225
rect 14458 7216 14464 7228
rect 14516 7216 14522 7268
rect 14550 7216 14556 7268
rect 14608 7256 14614 7268
rect 16316 7256 16344 7296
rect 16485 7293 16497 7327
rect 16531 7324 16543 7327
rect 16666 7324 16672 7336
rect 16531 7296 16672 7324
rect 16531 7293 16543 7296
rect 16485 7287 16543 7293
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 17052 7333 17080 7432
rect 17037 7327 17095 7333
rect 17037 7293 17049 7327
rect 17083 7293 17095 7327
rect 18046 7324 18052 7336
rect 18007 7296 18052 7324
rect 17037 7287 17095 7293
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 17313 7259 17371 7265
rect 17313 7256 17325 7259
rect 14608 7228 16252 7256
rect 16316 7228 17325 7256
rect 14608 7216 14614 7228
rect 3237 7191 3295 7197
rect 3237 7188 3249 7191
rect 3016 7160 3249 7188
rect 3016 7148 3022 7160
rect 3237 7157 3249 7160
rect 3283 7157 3295 7191
rect 3237 7151 3295 7157
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7188 3387 7191
rect 3697 7191 3755 7197
rect 3697 7188 3709 7191
rect 3375 7160 3709 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 3697 7157 3709 7160
rect 3743 7157 3755 7191
rect 3697 7151 3755 7157
rect 4065 7191 4123 7197
rect 4065 7157 4077 7191
rect 4111 7157 4123 7191
rect 4065 7151 4123 7157
rect 5626 7148 5632 7200
rect 5684 7188 5690 7200
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 5684 7160 6377 7188
rect 5684 7148 5690 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6604 7160 6837 7188
rect 6604 7148 6610 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 7282 7188 7288 7200
rect 7243 7160 7288 7188
rect 6825 7151 6883 7157
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 10781 7191 10839 7197
rect 10781 7157 10793 7191
rect 10827 7188 10839 7191
rect 10962 7188 10968 7200
rect 10827 7160 10968 7188
rect 10827 7157 10839 7160
rect 10781 7151 10839 7157
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 11790 7188 11796 7200
rect 11751 7160 11796 7188
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 13357 7191 13415 7197
rect 13357 7157 13369 7191
rect 13403 7188 13415 7191
rect 13998 7188 14004 7200
rect 13403 7160 14004 7188
rect 13403 7157 13415 7160
rect 13357 7151 13415 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 15562 7188 15568 7200
rect 15523 7160 15568 7188
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 16025 7191 16083 7197
rect 16025 7157 16037 7191
rect 16071 7188 16083 7191
rect 16114 7188 16120 7200
rect 16071 7160 16120 7188
rect 16071 7157 16083 7160
rect 16025 7151 16083 7157
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 16224 7188 16252 7228
rect 17313 7225 17325 7228
rect 17359 7225 17371 7259
rect 17313 7219 17371 7225
rect 16393 7191 16451 7197
rect 16393 7188 16405 7191
rect 16224 7160 16405 7188
rect 16393 7157 16405 7160
rect 16439 7188 16451 7191
rect 16482 7188 16488 7200
rect 16439 7160 16488 7188
rect 16439 7157 16451 7160
rect 16393 7151 16451 7157
rect 16482 7148 16488 7160
rect 16540 7148 16546 7200
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 18233 7191 18291 7197
rect 18233 7188 18245 7191
rect 17920 7160 18245 7188
rect 17920 7148 17926 7160
rect 18233 7157 18245 7160
rect 18279 7157 18291 7191
rect 18233 7151 18291 7157
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 4430 6984 4436 6996
rect 2004 6956 4436 6984
rect 2004 6944 2010 6956
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 6270 6984 6276 6996
rect 6231 6956 6276 6984
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 6454 6944 6460 6996
rect 6512 6984 6518 6996
rect 7558 6984 7564 6996
rect 6512 6956 7420 6984
rect 7519 6956 7564 6984
rect 6512 6944 6518 6956
rect 3418 6916 3424 6928
rect 2976 6888 3424 6916
rect 2976 6860 3004 6888
rect 3418 6876 3424 6888
rect 3476 6876 3482 6928
rect 5534 6916 5540 6928
rect 5092 6888 5540 6916
rect 1664 6851 1722 6857
rect 1664 6817 1676 6851
rect 1710 6848 1722 6851
rect 2958 6848 2964 6860
rect 1710 6820 2964 6848
rect 1710 6817 1722 6820
rect 1664 6811 1722 6817
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 3053 6851 3111 6857
rect 3053 6817 3065 6851
rect 3099 6848 3111 6851
rect 3326 6848 3332 6860
rect 3099 6820 3332 6848
rect 3099 6817 3111 6820
rect 3053 6811 3111 6817
rect 3326 6808 3332 6820
rect 3384 6808 3390 6860
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6817 3847 6851
rect 4062 6848 4068 6860
rect 4023 6820 4068 6848
rect 3789 6811 3847 6817
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1412 6644 1440 6743
rect 2777 6715 2835 6721
rect 2777 6681 2789 6715
rect 2823 6712 2835 6715
rect 3050 6712 3056 6724
rect 2823 6684 3056 6712
rect 2823 6681 2835 6684
rect 2777 6675 2835 6681
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 3237 6715 3295 6721
rect 3237 6681 3249 6715
rect 3283 6712 3295 6715
rect 3694 6712 3700 6724
rect 3283 6684 3700 6712
rect 3283 6681 3295 6684
rect 3237 6675 3295 6681
rect 3694 6672 3700 6684
rect 3752 6672 3758 6724
rect 3804 6712 3832 6811
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4801 6851 4859 6857
rect 4801 6817 4813 6851
rect 4847 6848 4859 6851
rect 5092 6848 5120 6888
rect 5534 6876 5540 6888
rect 5592 6876 5598 6928
rect 6840 6888 7144 6916
rect 4847 6820 5120 6848
rect 5160 6851 5218 6857
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 5160 6817 5172 6851
rect 5206 6848 5218 6851
rect 6840 6848 6868 6888
rect 5206 6820 6868 6848
rect 6917 6851 6975 6857
rect 5206 6817 5218 6820
rect 5160 6811 5218 6817
rect 6917 6817 6929 6851
rect 6963 6817 6975 6851
rect 6917 6811 6975 6817
rect 4522 6740 4528 6792
rect 4580 6780 4586 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4580 6752 4905 6780
rect 4580 6740 4586 6752
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 4893 6743 4951 6749
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6932 6780 6960 6811
rect 7116 6789 7144 6888
rect 7392 6848 7420 6956
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 8110 6944 8116 6996
rect 8168 6984 8174 6996
rect 8168 6956 8248 6984
rect 8168 6944 8174 6956
rect 7926 6916 7932 6928
rect 7887 6888 7932 6916
rect 7926 6876 7932 6888
rect 7984 6876 7990 6928
rect 8220 6916 8248 6956
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8444 6956 8953 6984
rect 8444 6944 8450 6956
rect 8941 6953 8953 6956
rect 8987 6984 8999 6987
rect 9030 6984 9036 6996
rect 8987 6956 9036 6984
rect 8987 6953 8999 6956
rect 8941 6947 8999 6953
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 10505 6987 10563 6993
rect 10505 6953 10517 6987
rect 10551 6984 10563 6987
rect 10686 6984 10692 6996
rect 10551 6956 10692 6984
rect 10551 6953 10563 6956
rect 10505 6947 10563 6953
rect 10686 6944 10692 6956
rect 10744 6944 10750 6996
rect 10873 6987 10931 6993
rect 10873 6953 10885 6987
rect 10919 6984 10931 6987
rect 11238 6984 11244 6996
rect 10919 6956 11244 6984
rect 10919 6953 10931 6956
rect 10873 6947 10931 6953
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 13446 6984 13452 6996
rect 11788 6956 13452 6984
rect 8220 6888 8800 6916
rect 8772 6848 8800 6888
rect 9214 6876 9220 6928
rect 9272 6916 9278 6928
rect 9582 6916 9588 6928
rect 9272 6888 9588 6916
rect 9272 6876 9278 6888
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 9677 6851 9735 6857
rect 7392 6820 8708 6848
rect 8772 6820 9168 6848
rect 6696 6752 6960 6780
rect 7009 6783 7067 6789
rect 6696 6740 6702 6752
rect 7009 6749 7021 6783
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 8018 6780 8024 6792
rect 7147 6752 7880 6780
rect 7979 6752 8024 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 7024 6712 7052 6743
rect 7374 6712 7380 6724
rect 3804 6684 4660 6712
rect 7024 6684 7380 6712
rect 2498 6644 2504 6656
rect 1412 6616 2504 6644
rect 2498 6604 2504 6616
rect 2556 6644 2562 6656
rect 3602 6644 3608 6656
rect 2556 6616 3608 6644
rect 2556 6604 2562 6616
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 3786 6604 3792 6656
rect 3844 6644 3850 6656
rect 4632 6653 4660 6684
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 7852 6712 7880 6752
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 8128 6712 8156 6743
rect 8202 6712 8208 6724
rect 7852 6684 8208 6712
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 8570 6712 8576 6724
rect 8531 6684 8576 6712
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 8680 6712 8708 6820
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 9140 6789 9168 6820
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 10410 6848 10416 6860
rect 9723 6820 10416 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 11788 6857 11816 6956
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 13909 6987 13967 6993
rect 13909 6984 13921 6987
rect 13872 6956 13921 6984
rect 13872 6944 13878 6956
rect 13909 6953 13921 6956
rect 13955 6953 13967 6987
rect 13909 6947 13967 6953
rect 14182 6944 14188 6996
rect 14240 6984 14246 6996
rect 14277 6987 14335 6993
rect 14277 6984 14289 6987
rect 14240 6956 14289 6984
rect 14240 6944 14246 6956
rect 14277 6953 14289 6956
rect 14323 6953 14335 6987
rect 14277 6947 14335 6953
rect 14366 6944 14372 6996
rect 14424 6984 14430 6996
rect 14424 6956 14469 6984
rect 14424 6944 14430 6956
rect 13722 6876 13728 6928
rect 13780 6916 13786 6928
rect 18046 6916 18052 6928
rect 13780 6888 18052 6916
rect 13780 6876 13786 6888
rect 18046 6876 18052 6888
rect 18104 6876 18110 6928
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10888 6820 10977 6848
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8904 6752 9045 6780
rect 8904 6740 8910 6752
rect 9033 6749 9045 6752
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9272 6752 9873 6780
rect 9272 6740 9278 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10888 6780 10916 6820
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 11773 6851 11831 6857
rect 11773 6848 11785 6851
rect 10965 6811 11023 6817
rect 11072 6820 11785 6848
rect 11072 6792 11100 6820
rect 11773 6817 11785 6820
rect 11819 6817 11831 6851
rect 11773 6811 11831 6817
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 13173 6851 13231 6857
rect 12124 6820 12940 6848
rect 12124 6808 12130 6820
rect 11054 6780 11060 6792
rect 10376 6752 10916 6780
rect 11015 6752 11060 6780
rect 10376 6740 10382 6752
rect 10410 6712 10416 6724
rect 8680 6684 10416 6712
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 10888 6712 10916 6752
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 11204 6752 11529 6780
rect 11204 6740 11210 6752
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 12912 6721 12940 6820
rect 13173 6817 13185 6851
rect 13219 6848 13231 6851
rect 13262 6848 13268 6860
rect 13219 6820 13268 6848
rect 13219 6817 13231 6820
rect 13173 6811 13231 6817
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 15740 6851 15798 6857
rect 15740 6817 15752 6851
rect 15786 6848 15798 6851
rect 16574 6848 16580 6860
rect 15786 6820 16580 6848
rect 15786 6817 15798 6820
rect 15740 6811 15798 6817
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 17126 6808 17132 6860
rect 17184 6848 17190 6860
rect 17497 6851 17555 6857
rect 17497 6848 17509 6851
rect 17184 6820 17509 6848
rect 17184 6808 17190 6820
rect 17497 6817 17509 6820
rect 17543 6817 17555 6851
rect 17497 6811 17555 6817
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13357 6783 13415 6789
rect 13357 6780 13369 6783
rect 13136 6752 13369 6780
rect 13136 6740 13142 6752
rect 13357 6749 13369 6752
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 14516 6752 14561 6780
rect 14516 6740 14522 6752
rect 15102 6740 15108 6792
rect 15160 6780 15166 6792
rect 15473 6783 15531 6789
rect 15473 6780 15485 6783
rect 15160 6752 15485 6780
rect 15160 6740 15166 6752
rect 15473 6749 15485 6752
rect 15519 6749 15531 6783
rect 15473 6743 15531 6749
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 17276 6752 17601 6780
rect 17276 6740 17282 6752
rect 17589 6749 17601 6752
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 17678 6740 17684 6792
rect 17736 6780 17742 6792
rect 18138 6780 18144 6792
rect 17736 6752 17781 6780
rect 18099 6752 18144 6780
rect 17736 6740 17742 6752
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 12897 6715 12955 6721
rect 10888 6684 11376 6712
rect 4249 6647 4307 6653
rect 4249 6644 4261 6647
rect 3844 6616 4261 6644
rect 3844 6604 3850 6616
rect 4249 6613 4261 6616
rect 4295 6613 4307 6647
rect 4249 6607 4307 6613
rect 4617 6647 4675 6653
rect 4617 6613 4629 6647
rect 4663 6644 4675 6647
rect 5994 6644 6000 6656
rect 4663 6616 6000 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 7190 6644 7196 6656
rect 6595 6616 7196 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7558 6604 7564 6656
rect 7616 6644 7622 6656
rect 11238 6644 11244 6656
rect 7616 6616 11244 6644
rect 7616 6604 7622 6616
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 11348 6644 11376 6684
rect 12897 6681 12909 6715
rect 12943 6681 12955 6715
rect 12897 6675 12955 6681
rect 12986 6672 12992 6724
rect 13044 6712 13050 6724
rect 14366 6712 14372 6724
rect 13044 6684 14372 6712
rect 13044 6672 13050 6684
rect 14366 6672 14372 6684
rect 14424 6672 14430 6724
rect 16758 6712 16764 6724
rect 16408 6684 16764 6712
rect 16408 6644 16436 6684
rect 16758 6672 16764 6684
rect 16816 6672 16822 6724
rect 16850 6644 16856 6656
rect 11348 6616 16436 6644
rect 16811 6616 16856 6644
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17218 6644 17224 6656
rect 17175 6616 17224 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 2222 6440 2228 6452
rect 1811 6412 2228 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 6178 6440 6184 6452
rect 3476 6412 6184 6440
rect 3476 6400 3482 6412
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 7466 6440 7472 6452
rect 6328 6412 7472 6440
rect 6328 6400 6334 6412
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 8202 6440 8208 6452
rect 8163 6412 8208 6440
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8294 6400 8300 6452
rect 8352 6400 8358 6452
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 13998 6440 14004 6452
rect 10468 6412 13124 6440
rect 13959 6412 14004 6440
rect 10468 6400 10474 6412
rect 2498 6372 2504 6384
rect 2240 6344 2504 6372
rect 2240 6316 2268 6344
rect 2498 6332 2504 6344
rect 2556 6372 2562 6384
rect 2556 6344 2820 6372
rect 2556 6332 2562 6344
rect 2222 6264 2228 6316
rect 2280 6264 2286 6316
rect 2792 6313 2820 6344
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6304 2467 6307
rect 2777 6307 2835 6313
rect 2455 6276 2728 6304
rect 2455 6273 2467 6276
rect 2409 6267 2467 6273
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6236 2191 6239
rect 2590 6236 2596 6248
rect 2179 6208 2596 6236
rect 2179 6205 2191 6208
rect 2133 6199 2191 6205
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 2700 6168 2728 6276
rect 2777 6273 2789 6307
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 5810 6304 5816 6316
rect 5592 6276 5816 6304
rect 5592 6264 5598 6276
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8312 6304 8340 6400
rect 10045 6375 10103 6381
rect 10045 6341 10057 6375
rect 10091 6372 10103 6375
rect 10134 6372 10140 6384
rect 10091 6344 10140 6372
rect 10091 6341 10103 6344
rect 10045 6335 10103 6341
rect 10134 6332 10140 6344
rect 10192 6332 10198 6384
rect 12710 6332 12716 6384
rect 12768 6372 12774 6384
rect 12989 6375 13047 6381
rect 12989 6372 13001 6375
rect 12768 6344 13001 6372
rect 12768 6332 12774 6344
rect 12989 6341 13001 6344
rect 13035 6341 13047 6375
rect 13096 6372 13124 6412
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 14366 6400 14372 6452
rect 14424 6440 14430 6452
rect 15378 6440 15384 6452
rect 14424 6412 15384 6440
rect 14424 6400 14430 6412
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 13096 6344 15700 6372
rect 12989 6335 13047 6341
rect 8260 6276 8340 6304
rect 10152 6304 10180 6332
rect 10152 6276 10272 6304
rect 8260 6264 8266 6276
rect 3050 6245 3056 6248
rect 3044 6199 3056 6245
rect 3108 6236 3114 6248
rect 3108 6208 3144 6236
rect 3050 6196 3056 6199
rect 3108 6196 3114 6208
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 4433 6239 4491 6245
rect 4433 6236 4445 6239
rect 3660 6208 4445 6236
rect 3660 6196 3666 6208
rect 4433 6205 4445 6208
rect 4479 6236 4491 6239
rect 4522 6236 4528 6248
rect 4479 6208 4528 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6236 6147 6239
rect 6454 6236 6460 6248
rect 6135 6208 6460 6236
rect 6135 6205 6147 6208
rect 6089 6199 6147 6205
rect 6454 6196 6460 6208
rect 6512 6196 6518 6248
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 2958 6168 2964 6180
rect 2700 6140 2964 6168
rect 2958 6128 2964 6140
rect 3016 6168 3022 6180
rect 4614 6168 4620 6180
rect 3016 6140 3096 6168
rect 3016 6128 3022 6140
rect 3068 6112 3096 6140
rect 4172 6140 4620 6168
rect 2225 6103 2283 6109
rect 2225 6069 2237 6103
rect 2271 6100 2283 6103
rect 2866 6100 2872 6112
rect 2271 6072 2872 6100
rect 2271 6069 2283 6072
rect 2225 6063 2283 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 3050 6060 3056 6112
rect 3108 6060 3114 6112
rect 4172 6109 4200 6140
rect 4614 6128 4620 6140
rect 4672 6177 4678 6180
rect 4672 6171 4736 6177
rect 4672 6137 4690 6171
rect 4724 6137 4736 6171
rect 4672 6131 4736 6137
rect 4816 6140 6316 6168
rect 4672 6128 4678 6131
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6069 4215 6103
rect 4157 6063 4215 6069
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 4816 6100 4844 6140
rect 4580 6072 4844 6100
rect 5813 6103 5871 6109
rect 4580 6060 4586 6072
rect 5813 6069 5825 6103
rect 5859 6100 5871 6103
rect 5902 6100 5908 6112
rect 5859 6072 5908 6100
rect 5859 6069 5871 6072
rect 5813 6063 5871 6069
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 6288 6109 6316 6140
rect 6273 6103 6331 6109
rect 6273 6069 6285 6103
rect 6319 6069 6331 6103
rect 6273 6063 6331 6069
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 6840 6100 6868 6199
rect 8570 6196 8576 6248
rect 8628 6236 8634 6248
rect 8665 6239 8723 6245
rect 8665 6236 8677 6239
rect 8628 6208 8677 6236
rect 8628 6196 8634 6208
rect 8665 6205 8677 6208
rect 8711 6205 8723 6239
rect 10137 6239 10195 6245
rect 10137 6236 10149 6239
rect 8665 6199 8723 6205
rect 8772 6208 10149 6236
rect 7092 6171 7150 6177
rect 7092 6137 7104 6171
rect 7138 6168 7150 6171
rect 7466 6168 7472 6180
rect 7138 6140 7472 6168
rect 7138 6137 7150 6140
rect 7092 6131 7150 6137
rect 7466 6128 7472 6140
rect 7524 6128 7530 6180
rect 8772 6168 8800 6208
rect 10137 6205 10149 6208
rect 10183 6205 10195 6239
rect 10244 6236 10272 6276
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 12216 6276 12449 6304
rect 12216 6264 12222 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 13633 6307 13691 6313
rect 13633 6273 13645 6307
rect 13679 6304 13691 6307
rect 13722 6304 13728 6316
rect 13679 6276 13728 6304
rect 13679 6273 13691 6276
rect 13633 6267 13691 6273
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 14458 6264 14464 6316
rect 14516 6304 14522 6316
rect 14553 6307 14611 6313
rect 14553 6304 14565 6307
rect 14516 6276 14565 6304
rect 14516 6264 14522 6276
rect 14553 6273 14565 6276
rect 14599 6304 14611 6307
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 14599 6276 15577 6304
rect 14599 6273 14611 6276
rect 14553 6267 14611 6273
rect 15565 6273 15577 6276
rect 15611 6273 15623 6307
rect 15672 6304 15700 6344
rect 15672 6276 16436 6304
rect 15565 6267 15623 6273
rect 10393 6239 10451 6245
rect 10393 6236 10405 6239
rect 10244 6208 10405 6236
rect 10137 6199 10195 6205
rect 10393 6205 10405 6208
rect 10439 6205 10451 6239
rect 10393 6199 10451 6205
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6205 12311 6239
rect 12253 6199 12311 6205
rect 7576 6140 8800 6168
rect 8932 6171 8990 6177
rect 7576 6100 7604 6140
rect 8932 6137 8944 6171
rect 8978 6168 8990 6171
rect 11330 6168 11336 6180
rect 8978 6140 11336 6168
rect 8978 6137 8990 6140
rect 8932 6131 8990 6137
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 11974 6128 11980 6180
rect 12032 6168 12038 6180
rect 12268 6168 12296 6199
rect 15102 6196 15108 6248
rect 15160 6236 15166 6248
rect 16301 6239 16359 6245
rect 16301 6236 16313 6239
rect 15160 6208 16313 6236
rect 15160 6196 15166 6208
rect 16301 6205 16313 6208
rect 16347 6205 16359 6239
rect 16408 6236 16436 6276
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 16408 6208 18061 6236
rect 16301 6199 16359 6205
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 12032 6140 12296 6168
rect 13357 6171 13415 6177
rect 12032 6128 12038 6140
rect 13357 6137 13369 6171
rect 13403 6168 13415 6171
rect 13630 6168 13636 6180
rect 13403 6140 13636 6168
rect 13403 6137 13415 6140
rect 13357 6131 13415 6137
rect 13630 6128 13636 6140
rect 13688 6128 13694 6180
rect 13814 6128 13820 6180
rect 13872 6168 13878 6180
rect 15470 6168 15476 6180
rect 13872 6140 15476 6168
rect 13872 6128 13878 6140
rect 15470 6128 15476 6140
rect 15528 6128 15534 6180
rect 16568 6171 16626 6177
rect 16568 6137 16580 6171
rect 16614 6168 16626 6171
rect 16850 6168 16856 6180
rect 16614 6140 16856 6168
rect 16614 6137 16626 6140
rect 16568 6131 16626 6137
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 17310 6128 17316 6180
rect 17368 6168 17374 6180
rect 17368 6140 17816 6168
rect 17368 6128 17374 6140
rect 17788 6112 17816 6140
rect 6788 6072 7604 6100
rect 6788 6060 6794 6072
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 11238 6100 11244 6112
rect 8536 6072 11244 6100
rect 8536 6060 8542 6072
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 11517 6103 11575 6109
rect 11517 6069 11529 6103
rect 11563 6100 11575 6103
rect 11606 6100 11612 6112
rect 11563 6072 11612 6100
rect 11563 6069 11575 6072
rect 11517 6063 11575 6069
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 12066 6100 12072 6112
rect 12027 6072 12072 6100
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 13446 6100 13452 6112
rect 13407 6072 13452 6100
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 13906 6060 13912 6112
rect 13964 6100 13970 6112
rect 14090 6100 14096 6112
rect 13964 6072 14096 6100
rect 13964 6060 13970 6072
rect 14090 6060 14096 6072
rect 14148 6100 14154 6112
rect 14369 6103 14427 6109
rect 14369 6100 14381 6103
rect 14148 6072 14381 6100
rect 14148 6060 14154 6072
rect 14369 6069 14381 6072
rect 14415 6069 14427 6103
rect 14369 6063 14427 6069
rect 14461 6103 14519 6109
rect 14461 6069 14473 6103
rect 14507 6100 14519 6103
rect 14550 6100 14556 6112
rect 14507 6072 14556 6100
rect 14507 6069 14519 6072
rect 14461 6063 14519 6069
rect 14550 6060 14556 6072
rect 14608 6100 14614 6112
rect 14734 6100 14740 6112
rect 14608 6072 14740 6100
rect 14608 6060 14614 6072
rect 14734 6060 14740 6072
rect 14792 6060 14798 6112
rect 14918 6060 14924 6112
rect 14976 6100 14982 6112
rect 15013 6103 15071 6109
rect 15013 6100 15025 6103
rect 14976 6072 15025 6100
rect 14976 6060 14982 6072
rect 15013 6069 15025 6072
rect 15059 6069 15071 6103
rect 15013 6063 15071 6069
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 15378 6100 15384 6112
rect 15252 6072 15384 6100
rect 15252 6060 15258 6072
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 15654 6060 15660 6112
rect 15712 6100 15718 6112
rect 17681 6103 17739 6109
rect 17681 6100 17693 6103
rect 15712 6072 17693 6100
rect 15712 6060 15718 6072
rect 17681 6069 17693 6072
rect 17727 6069 17739 6103
rect 17681 6063 17739 6069
rect 17770 6060 17776 6112
rect 17828 6060 17834 6112
rect 18230 6100 18236 6112
rect 18191 6072 18236 6100
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 1857 5899 1915 5905
rect 1857 5865 1869 5899
rect 1903 5896 1915 5899
rect 2314 5896 2320 5908
rect 1903 5868 2320 5896
rect 1903 5865 1915 5868
rect 1857 5859 1915 5865
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 2866 5896 2872 5908
rect 2827 5868 2872 5896
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 4028 5868 4077 5896
rect 4028 5856 4034 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4430 5896 4436 5908
rect 4391 5868 4436 5896
rect 4065 5859 4123 5865
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 4982 5856 4988 5908
rect 5040 5896 5046 5908
rect 5445 5899 5503 5905
rect 5445 5896 5457 5899
rect 5040 5868 5457 5896
rect 5040 5856 5046 5868
rect 5445 5865 5457 5868
rect 5491 5865 5503 5899
rect 5445 5859 5503 5865
rect 6638 5856 6644 5908
rect 6696 5896 6702 5908
rect 6917 5899 6975 5905
rect 6917 5896 6929 5899
rect 6696 5868 6929 5896
rect 6696 5856 6702 5868
rect 6917 5865 6929 5868
rect 6963 5865 6975 5899
rect 6917 5859 6975 5865
rect 7929 5899 7987 5905
rect 7929 5865 7941 5899
rect 7975 5896 7987 5899
rect 8018 5896 8024 5908
rect 7975 5868 8024 5896
rect 7975 5865 7987 5868
rect 7929 5859 7987 5865
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 9861 5899 9919 5905
rect 9861 5896 9873 5899
rect 8128 5868 9873 5896
rect 1762 5788 1768 5840
rect 1820 5828 1826 5840
rect 3329 5831 3387 5837
rect 3329 5828 3341 5831
rect 1820 5800 3341 5828
rect 1820 5788 1826 5800
rect 3329 5797 3341 5800
rect 3375 5797 3387 5831
rect 3329 5791 3387 5797
rect 4246 5788 4252 5840
rect 4304 5828 4310 5840
rect 8128 5828 8156 5868
rect 9861 5865 9873 5868
rect 9907 5865 9919 5899
rect 9861 5859 9919 5865
rect 10321 5899 10379 5905
rect 10321 5865 10333 5899
rect 10367 5896 10379 5899
rect 10778 5896 10784 5908
rect 10367 5868 10784 5896
rect 10367 5865 10379 5868
rect 10321 5859 10379 5865
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 11238 5856 11244 5908
rect 11296 5896 11302 5908
rect 12618 5896 12624 5908
rect 11296 5868 12624 5896
rect 11296 5856 11302 5868
rect 12618 5856 12624 5868
rect 12676 5896 12682 5908
rect 13170 5896 13176 5908
rect 12676 5868 13176 5896
rect 12676 5856 12682 5868
rect 13170 5856 13176 5868
rect 13228 5856 13234 5908
rect 14185 5899 14243 5905
rect 14185 5865 14197 5899
rect 14231 5896 14243 5899
rect 14458 5896 14464 5908
rect 14231 5868 14464 5896
rect 14231 5865 14243 5868
rect 14185 5859 14243 5865
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 15841 5899 15899 5905
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16114 5896 16120 5908
rect 15887 5868 16120 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 17313 5899 17371 5905
rect 17313 5865 17325 5899
rect 17359 5896 17371 5899
rect 18138 5896 18144 5908
rect 17359 5868 18144 5896
rect 17359 5865 17371 5868
rect 17313 5859 17371 5865
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 4304 5800 8156 5828
rect 8297 5831 8355 5837
rect 4304 5788 4310 5800
rect 8297 5797 8309 5831
rect 8343 5828 8355 5831
rect 8938 5828 8944 5840
rect 8343 5800 8944 5828
rect 8343 5797 8355 5800
rect 8297 5791 8355 5797
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 9030 5788 9036 5840
rect 9088 5828 9094 5840
rect 10045 5831 10103 5837
rect 10045 5828 10057 5831
rect 9088 5800 10057 5828
rect 9088 5788 9094 5800
rect 10045 5797 10057 5800
rect 10091 5797 10103 5831
rect 10045 5791 10103 5797
rect 10410 5788 10416 5840
rect 10468 5828 10474 5840
rect 10468 5800 10824 5828
rect 10468 5788 10474 5800
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 3142 5760 3148 5772
rect 2271 5732 3148 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 3142 5720 3148 5732
rect 3200 5720 3206 5772
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 3283 5732 4108 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 2314 5692 2320 5704
rect 2275 5664 2320 5692
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5692 2559 5695
rect 3050 5692 3056 5704
rect 2547 5664 3056 5692
rect 2547 5661 2559 5664
rect 2501 5655 2559 5661
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 2866 5624 2872 5636
rect 2740 5596 2872 5624
rect 2740 5584 2746 5596
rect 2866 5584 2872 5596
rect 2924 5584 2930 5636
rect 2498 5516 2504 5568
rect 2556 5556 2562 5568
rect 3326 5556 3332 5568
rect 2556 5528 3332 5556
rect 2556 5516 2562 5528
rect 3326 5516 3332 5528
rect 3384 5556 3390 5568
rect 3436 5556 3464 5655
rect 3602 5584 3608 5636
rect 3660 5624 3666 5636
rect 3970 5624 3976 5636
rect 3660 5596 3976 5624
rect 3660 5584 3666 5596
rect 3970 5584 3976 5596
rect 4028 5584 4034 5636
rect 3384 5528 3464 5556
rect 4080 5556 4108 5732
rect 4338 5720 4344 5772
rect 4396 5760 4402 5772
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 4396 5732 4537 5760
rect 4396 5720 4402 5732
rect 4525 5729 4537 5732
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 4890 5720 4896 5772
rect 4948 5760 4954 5772
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 4948 5732 5549 5760
rect 4948 5720 4954 5732
rect 5537 5729 5549 5732
rect 5583 5729 5595 5763
rect 5902 5760 5908 5772
rect 5537 5723 5595 5729
rect 5736 5732 5908 5760
rect 4614 5652 4620 5704
rect 4672 5692 4678 5704
rect 4672 5664 4717 5692
rect 4672 5652 4678 5664
rect 4798 5652 4804 5704
rect 4856 5692 4862 5704
rect 5350 5692 5356 5704
rect 4856 5664 5356 5692
rect 4856 5652 4862 5664
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5736 5701 5764 5732
rect 5902 5720 5908 5732
rect 5960 5720 5966 5772
rect 6089 5763 6147 5769
rect 6089 5729 6101 5763
rect 6135 5760 6147 5763
rect 6178 5760 6184 5772
rect 6135 5732 6184 5760
rect 6135 5729 6147 5732
rect 6089 5723 6147 5729
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 6362 5720 6368 5772
rect 6420 5760 6426 5772
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 6420 5732 7297 5760
rect 6420 5720 6426 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 9122 5760 9128 5772
rect 7285 5723 7343 5729
rect 7392 5732 8708 5760
rect 9083 5732 9128 5760
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 7392 5701 7420 5732
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 5868 5664 6285 5692
rect 5868 5652 5874 5664
rect 6273 5661 6285 5664
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 7392 5624 7420 5655
rect 7466 5652 7472 5704
rect 7524 5692 7530 5704
rect 8389 5695 8447 5701
rect 7524 5664 7569 5692
rect 7524 5652 7530 5664
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 8478 5692 8484 5704
rect 8435 5664 8484 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5661 8631 5695
rect 8680 5692 8708 5732
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 9677 5763 9735 5769
rect 9232 5732 9527 5760
rect 9232 5701 9260 5732
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 8680 5664 9229 5692
rect 8573 5655 8631 5661
rect 9217 5661 9229 5664
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 4764 5596 7420 5624
rect 7484 5624 7512 5652
rect 8588 5624 8616 5655
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 9499 5692 9527 5732
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10318 5760 10324 5772
rect 9723 5732 10324 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 10796 5769 10824 5800
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 13050 5831 13108 5837
rect 13050 5828 13062 5831
rect 12584 5800 13062 5828
rect 12584 5788 12590 5800
rect 13050 5797 13062 5800
rect 13096 5797 13108 5831
rect 15102 5828 15108 5840
rect 13050 5791 13108 5797
rect 14384 5800 15108 5828
rect 10689 5763 10747 5769
rect 10689 5729 10701 5763
rect 10735 5729 10747 5763
rect 10689 5723 10747 5729
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5729 10839 5763
rect 11146 5760 11152 5772
rect 11107 5732 11152 5760
rect 10781 5723 10839 5729
rect 10410 5692 10416 5704
rect 9364 5664 9409 5692
rect 9499 5664 10416 5692
rect 9364 5652 9370 5664
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10704 5692 10732 5723
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 11416 5763 11474 5769
rect 11416 5729 11428 5763
rect 11462 5760 11474 5763
rect 12158 5760 12164 5772
rect 11462 5732 12164 5760
rect 11462 5729 11474 5732
rect 11416 5723 11474 5729
rect 12158 5720 12164 5732
rect 12216 5720 12222 5772
rect 12805 5763 12863 5769
rect 12805 5729 12817 5763
rect 12851 5760 12863 5763
rect 14384 5760 14412 5800
rect 15102 5788 15108 5800
rect 15160 5788 15166 5840
rect 15749 5831 15807 5837
rect 15749 5797 15761 5831
rect 15795 5828 15807 5831
rect 16942 5828 16948 5840
rect 15795 5800 16948 5828
rect 15795 5797 15807 5800
rect 15749 5791 15807 5797
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 17402 5788 17408 5840
rect 17460 5788 17466 5840
rect 12851 5732 14412 5760
rect 14461 5763 14519 5769
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 14461 5729 14473 5763
rect 14507 5760 14519 5763
rect 15010 5760 15016 5772
rect 14507 5732 15016 5760
rect 14507 5729 14519 5732
rect 14461 5723 14519 5729
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 16393 5763 16451 5769
rect 16393 5760 16405 5763
rect 15528 5732 16405 5760
rect 15528 5720 15534 5732
rect 16393 5729 16405 5732
rect 16439 5729 16451 5763
rect 17420 5760 17448 5788
rect 17957 5763 18015 5769
rect 17957 5760 17969 5763
rect 17420 5732 17969 5760
rect 16393 5723 16451 5729
rect 17957 5729 17969 5732
rect 18003 5729 18015 5763
rect 17957 5723 18015 5729
rect 10965 5695 11023 5701
rect 10704 5664 10916 5692
rect 7484 5596 8616 5624
rect 4764 5584 4770 5596
rect 8938 5584 8944 5636
rect 8996 5624 9002 5636
rect 9324 5624 9352 5652
rect 8996 5596 9352 5624
rect 8996 5584 9002 5596
rect 4798 5556 4804 5568
rect 4080 5528 4804 5556
rect 3384 5516 3390 5528
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 5074 5556 5080 5568
rect 5035 5528 5080 5556
rect 5074 5516 5080 5528
rect 5132 5516 5138 5568
rect 5994 5516 6000 5568
rect 6052 5556 6058 5568
rect 7190 5556 7196 5568
rect 6052 5528 7196 5556
rect 6052 5516 6058 5528
rect 7190 5516 7196 5528
rect 7248 5516 7254 5568
rect 7558 5516 7564 5568
rect 7616 5556 7622 5568
rect 8018 5556 8024 5568
rect 7616 5528 8024 5556
rect 7616 5516 7622 5528
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 8757 5559 8815 5565
rect 8757 5556 8769 5559
rect 8260 5528 8769 5556
rect 8260 5516 8266 5528
rect 8757 5525 8769 5528
rect 8803 5525 8815 5559
rect 10888 5556 10916 5664
rect 10965 5661 10977 5695
rect 11011 5692 11023 5695
rect 11054 5692 11060 5704
rect 11011 5664 11060 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 13964 5664 14657 5692
rect 13964 5652 13970 5664
rect 14645 5661 14657 5664
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 14734 5652 14740 5704
rect 14792 5692 14798 5704
rect 16025 5695 16083 5701
rect 14792 5664 15976 5692
rect 14792 5652 14798 5664
rect 12526 5624 12532 5636
rect 12487 5596 12532 5624
rect 12526 5584 12532 5596
rect 12584 5584 12590 5636
rect 14182 5584 14188 5636
rect 14240 5624 14246 5636
rect 14918 5624 14924 5636
rect 14240 5596 14924 5624
rect 14240 5584 14246 5596
rect 14918 5584 14924 5596
rect 14976 5584 14982 5636
rect 11054 5556 11060 5568
rect 10888 5528 11060 5556
rect 8757 5519 8815 5525
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 15378 5556 15384 5568
rect 15339 5528 15384 5556
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 15948 5556 15976 5664
rect 16025 5661 16037 5695
rect 16071 5692 16083 5695
rect 16298 5692 16304 5704
rect 16071 5664 16304 5692
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 16298 5652 16304 5664
rect 16356 5692 16362 5704
rect 17310 5692 17316 5704
rect 16356 5664 17316 5692
rect 16356 5652 16362 5664
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5692 17647 5695
rect 17678 5692 17684 5704
rect 17635 5664 17684 5692
rect 17635 5661 17647 5664
rect 17589 5655 17647 5661
rect 17420 5624 17448 5655
rect 17678 5652 17684 5664
rect 17736 5652 17742 5704
rect 16408 5596 17448 5624
rect 16408 5556 16436 5596
rect 16574 5556 16580 5568
rect 15948 5528 16436 5556
rect 16535 5528 16580 5556
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 16942 5556 16948 5568
rect 16903 5528 16948 5556
rect 16942 5516 16948 5528
rect 17000 5516 17006 5568
rect 17862 5516 17868 5568
rect 17920 5556 17926 5568
rect 18141 5559 18199 5565
rect 18141 5556 18153 5559
rect 17920 5528 18153 5556
rect 17920 5516 17926 5528
rect 18141 5525 18153 5528
rect 18187 5525 18199 5559
rect 18141 5519 18199 5525
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3697 5355 3755 5361
rect 3697 5352 3709 5355
rect 3108 5324 3709 5352
rect 3108 5312 3114 5324
rect 3697 5321 3709 5324
rect 3743 5321 3755 5355
rect 4982 5352 4988 5364
rect 3697 5315 3755 5321
rect 3896 5324 4988 5352
rect 3896 5296 3924 5324
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 5350 5312 5356 5364
rect 5408 5352 5414 5364
rect 6641 5355 6699 5361
rect 6641 5352 6653 5355
rect 5408 5324 6653 5352
rect 5408 5312 5414 5324
rect 6641 5321 6653 5324
rect 6687 5321 6699 5355
rect 6641 5315 6699 5321
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 7374 5352 7380 5364
rect 6871 5324 7380 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 7837 5355 7895 5361
rect 7837 5321 7849 5355
rect 7883 5352 7895 5355
rect 7926 5352 7932 5364
rect 7883 5324 7932 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 11333 5355 11391 5361
rect 11333 5321 11345 5355
rect 11379 5352 11391 5355
rect 11790 5352 11796 5364
rect 11379 5324 11796 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 13504 5324 13553 5352
rect 13504 5312 13510 5324
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 13541 5315 13599 5321
rect 14182 5312 14188 5364
rect 14240 5352 14246 5364
rect 14550 5352 14556 5364
rect 14240 5324 14556 5352
rect 14240 5312 14246 5324
rect 14550 5312 14556 5324
rect 14608 5352 14614 5364
rect 17954 5352 17960 5364
rect 14608 5324 17960 5352
rect 14608 5312 14614 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 3878 5244 3884 5296
rect 3936 5244 3942 5296
rect 9030 5284 9036 5296
rect 8496 5256 9036 5284
rect 4430 5216 4436 5228
rect 1688 5188 2452 5216
rect 1688 5157 1716 5188
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5117 1731 5151
rect 1673 5111 1731 5117
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5117 2375 5151
rect 2424 5148 2452 5188
rect 3896 5188 4436 5216
rect 3896 5148 3924 5188
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 4614 5216 4620 5228
rect 4575 5188 4620 5216
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 5902 5216 5908 5228
rect 5644 5188 5908 5216
rect 2424 5120 3924 5148
rect 3973 5151 4031 5157
rect 2317 5111 2375 5117
rect 3973 5117 3985 5151
rect 4019 5148 4031 5151
rect 4884 5151 4942 5157
rect 4019 5120 4844 5148
rect 4019 5117 4031 5120
rect 3973 5111 4031 5117
rect 1394 5040 1400 5092
rect 1452 5080 1458 5092
rect 2222 5080 2228 5092
rect 1452 5052 2228 5080
rect 1452 5040 1458 5052
rect 2222 5040 2228 5052
rect 2280 5080 2286 5092
rect 2332 5080 2360 5111
rect 4816 5092 4844 5120
rect 4884 5117 4896 5151
rect 4930 5148 4942 5151
rect 5644 5148 5672 5188
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 7466 5176 7472 5188
rect 7524 5216 7530 5228
rect 8386 5216 8392 5228
rect 7524 5188 8392 5216
rect 7524 5176 7530 5188
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 4930 5120 5672 5148
rect 8205 5151 8263 5157
rect 4930 5117 4942 5120
rect 4884 5111 4942 5117
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8496 5148 8524 5256
rect 9030 5244 9036 5256
rect 9088 5244 9094 5296
rect 10410 5284 10416 5296
rect 10323 5256 10416 5284
rect 10410 5244 10416 5256
rect 10468 5284 10474 5296
rect 12158 5284 12164 5296
rect 10468 5256 11008 5284
rect 10468 5244 10474 5256
rect 8251 5120 8524 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8570 5108 8576 5160
rect 8628 5148 8634 5160
rect 9030 5148 9036 5160
rect 8628 5120 9036 5148
rect 8628 5108 8634 5120
rect 9030 5108 9036 5120
rect 9088 5108 9094 5160
rect 10980 5148 11008 5256
rect 11992 5256 12164 5284
rect 11992 5225 12020 5256
rect 12158 5244 12164 5256
rect 12216 5284 12222 5296
rect 13722 5284 13728 5296
rect 12216 5256 13728 5284
rect 12216 5244 12222 5256
rect 13722 5244 13728 5256
rect 13780 5244 13786 5296
rect 16482 5244 16488 5296
rect 16540 5284 16546 5296
rect 16540 5256 18092 5284
rect 16540 5244 16546 5256
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 12894 5216 12900 5228
rect 12855 5188 12900 5216
rect 11977 5179 12035 5185
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 13127 5188 14197 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 14185 5185 14197 5188
rect 14231 5216 14243 5219
rect 14274 5216 14280 5228
rect 14231 5188 14280 5216
rect 14231 5185 14243 5188
rect 14185 5179 14243 5185
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 15102 5216 15108 5228
rect 15063 5188 15108 5216
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 13262 5148 13268 5160
rect 10980 5120 13268 5148
rect 13262 5108 13268 5120
rect 13320 5108 13326 5160
rect 13446 5108 13452 5160
rect 13504 5148 13510 5160
rect 13909 5151 13967 5157
rect 13504 5120 13676 5148
rect 13504 5108 13510 5120
rect 2280 5052 2360 5080
rect 2280 5040 2286 5052
rect 2498 5040 2504 5092
rect 2556 5089 2562 5092
rect 2556 5083 2620 5089
rect 2556 5049 2574 5083
rect 2608 5049 2620 5083
rect 2556 5043 2620 5049
rect 2556 5040 2562 5043
rect 4798 5040 4804 5092
rect 4856 5040 4862 5092
rect 9300 5083 9358 5089
rect 9300 5049 9312 5083
rect 9346 5080 9358 5083
rect 11606 5080 11612 5092
rect 9346 5052 11612 5080
rect 9346 5049 9358 5052
rect 9300 5043 9358 5049
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 11701 5083 11759 5089
rect 11701 5049 11713 5083
rect 11747 5080 11759 5083
rect 12805 5083 12863 5089
rect 11747 5052 12480 5080
rect 11747 5049 11759 5052
rect 11701 5043 11759 5049
rect 1857 5015 1915 5021
rect 1857 4981 1869 5015
rect 1903 5012 1915 5015
rect 3050 5012 3056 5024
rect 1903 4984 3056 5012
rect 1903 4981 1915 4984
rect 1857 4975 1915 4981
rect 3050 4972 3056 4984
rect 3108 4972 3114 5024
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 5012 4215 5015
rect 4338 5012 4344 5024
rect 4203 4984 4344 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 4614 5012 4620 5024
rect 4488 4984 4620 5012
rect 4488 4972 4494 4984
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 5994 5012 6000 5024
rect 5955 4984 6000 5012
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 6687 4984 7205 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 7193 4981 7205 4984
rect 7239 4981 7251 5015
rect 7193 4975 7251 4981
rect 7282 4972 7288 5024
rect 7340 5012 7346 5024
rect 7340 4984 7385 5012
rect 7340 4972 7346 4984
rect 8202 4972 8208 5024
rect 8260 5012 8266 5024
rect 8297 5015 8355 5021
rect 8297 5012 8309 5015
rect 8260 4984 8309 5012
rect 8260 4972 8266 4984
rect 8297 4981 8309 4984
rect 8343 5012 8355 5015
rect 8570 5012 8576 5024
rect 8343 4984 8576 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 8570 4972 8576 4984
rect 8628 4972 8634 5024
rect 9122 4972 9128 5024
rect 9180 5012 9186 5024
rect 10873 5015 10931 5021
rect 10873 5012 10885 5015
rect 9180 4984 10885 5012
rect 9180 4972 9186 4984
rect 10873 4981 10885 4984
rect 10919 4981 10931 5015
rect 11790 5012 11796 5024
rect 11751 4984 11796 5012
rect 10873 4975 10931 4981
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 12452 5021 12480 5052
rect 12805 5049 12817 5083
rect 12851 5080 12863 5083
rect 13538 5080 13544 5092
rect 12851 5052 13544 5080
rect 12851 5049 12863 5052
rect 12805 5043 12863 5049
rect 13538 5040 13544 5052
rect 13596 5040 13602 5092
rect 13648 5080 13676 5120
rect 13909 5117 13921 5151
rect 13955 5148 13967 5151
rect 14366 5148 14372 5160
rect 13955 5120 14372 5148
rect 13955 5117 13967 5120
rect 13909 5111 13967 5117
rect 14366 5108 14372 5120
rect 14424 5108 14430 5160
rect 15372 5151 15430 5157
rect 15372 5117 15384 5151
rect 15418 5148 15430 5151
rect 15654 5148 15660 5160
rect 15418 5120 15660 5148
rect 15418 5117 15430 5120
rect 15372 5111 15430 5117
rect 15654 5108 15660 5120
rect 15712 5108 15718 5160
rect 16500 5080 16528 5244
rect 17218 5216 17224 5228
rect 17179 5188 17224 5216
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 17310 5176 17316 5228
rect 17368 5216 17374 5228
rect 17368 5188 17413 5216
rect 17368 5176 17374 5188
rect 16574 5108 16580 5160
rect 16632 5148 16638 5160
rect 16758 5148 16764 5160
rect 16632 5120 16764 5148
rect 16632 5108 16638 5120
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 16942 5108 16948 5160
rect 17000 5148 17006 5160
rect 18064 5157 18092 5256
rect 17129 5151 17187 5157
rect 17129 5148 17141 5151
rect 17000 5120 17141 5148
rect 17000 5108 17006 5120
rect 17129 5117 17141 5120
rect 17175 5117 17187 5151
rect 17129 5111 17187 5117
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 13648 5052 16528 5080
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 4981 12495 5015
rect 12437 4975 12495 4981
rect 13170 4972 13176 5024
rect 13228 5012 13234 5024
rect 14001 5015 14059 5021
rect 14001 5012 14013 5015
rect 13228 4984 14013 5012
rect 13228 4972 13234 4984
rect 14001 4981 14013 4984
rect 14047 4981 14059 5015
rect 14550 5012 14556 5024
rect 14511 4984 14556 5012
rect 14001 4975 14059 4981
rect 14550 4972 14556 4984
rect 14608 4972 14614 5024
rect 16482 5012 16488 5024
rect 16443 4984 16488 5012
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 16758 5012 16764 5024
rect 16719 4984 16764 5012
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 2314 4768 2320 4820
rect 2372 4808 2378 4820
rect 2593 4811 2651 4817
rect 2593 4808 2605 4811
rect 2372 4780 2605 4808
rect 2372 4768 2378 4780
rect 2593 4777 2605 4780
rect 2639 4777 2651 4811
rect 2593 4771 2651 4777
rect 3142 4768 3148 4820
rect 3200 4808 3206 4820
rect 4065 4811 4123 4817
rect 4065 4808 4077 4811
rect 3200 4780 4077 4808
rect 3200 4768 3206 4780
rect 4065 4777 4077 4780
rect 4111 4777 4123 4811
rect 4430 4808 4436 4820
rect 4391 4780 4436 4808
rect 4065 4771 4123 4777
rect 4430 4768 4436 4780
rect 4488 4808 4494 4820
rect 4706 4808 4712 4820
rect 4488 4780 4712 4808
rect 4488 4768 4494 4780
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 5074 4768 5080 4820
rect 5132 4808 5138 4820
rect 5537 4811 5595 4817
rect 5537 4808 5549 4811
rect 5132 4780 5549 4808
rect 5132 4768 5138 4780
rect 5537 4777 5549 4780
rect 5583 4777 5595 4811
rect 5537 4771 5595 4777
rect 8386 4768 8392 4820
rect 8444 4808 8450 4820
rect 8481 4811 8539 4817
rect 8481 4808 8493 4811
rect 8444 4780 8493 4808
rect 8444 4768 8450 4780
rect 8481 4777 8493 4780
rect 8527 4777 8539 4811
rect 8481 4771 8539 4777
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 12158 4808 12164 4820
rect 8628 4780 12164 4808
rect 8628 4768 8634 4780
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 13446 4808 13452 4820
rect 12759 4780 13452 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 13722 4768 13728 4820
rect 13780 4808 13786 4820
rect 14921 4811 14979 4817
rect 14921 4808 14933 4811
rect 13780 4780 14933 4808
rect 13780 4768 13786 4780
rect 14921 4777 14933 4780
rect 14967 4777 14979 4811
rect 14921 4771 14979 4777
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4777 15347 4811
rect 15289 4771 15347 4777
rect 3878 4740 3884 4752
rect 2056 4712 3884 4740
rect 1486 4672 1492 4684
rect 1447 4644 1492 4672
rect 1486 4632 1492 4644
rect 1544 4632 1550 4684
rect 2056 4681 2084 4712
rect 3878 4700 3884 4712
rect 3936 4700 3942 4752
rect 3970 4700 3976 4752
rect 4028 4740 4034 4752
rect 5626 4740 5632 4752
rect 4028 4712 5632 4740
rect 4028 4700 4034 4712
rect 5626 4700 5632 4712
rect 5684 4700 5690 4752
rect 6362 4700 6368 4752
rect 6420 4740 6426 4752
rect 9033 4743 9091 4749
rect 9033 4740 9045 4743
rect 6420 4712 9045 4740
rect 6420 4700 6426 4712
rect 9033 4709 9045 4712
rect 9079 4709 9091 4743
rect 9033 4703 9091 4709
rect 10036 4743 10094 4749
rect 10036 4709 10048 4743
rect 10082 4740 10094 4743
rect 10410 4740 10416 4752
rect 10082 4712 10416 4740
rect 10082 4709 10094 4712
rect 10036 4703 10094 4709
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 13538 4740 13544 4752
rect 11480 4712 13544 4740
rect 11480 4700 11486 4712
rect 13538 4700 13544 4712
rect 13596 4700 13602 4752
rect 14090 4700 14096 4752
rect 14148 4740 14154 4752
rect 14366 4740 14372 4752
rect 14148 4712 14372 4740
rect 14148 4700 14154 4712
rect 14366 4700 14372 4712
rect 14424 4740 14430 4752
rect 14424 4712 15240 4740
rect 14424 4700 14430 4712
rect 2041 4675 2099 4681
rect 2041 4641 2053 4675
rect 2087 4641 2099 4675
rect 2041 4635 2099 4641
rect 2409 4675 2467 4681
rect 2409 4641 2421 4675
rect 2455 4672 2467 4675
rect 2590 4672 2596 4684
rect 2455 4644 2596 4672
rect 2455 4641 2467 4644
rect 2409 4635 2467 4641
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 2682 4632 2688 4684
rect 2740 4672 2746 4684
rect 2961 4675 3019 4681
rect 2961 4672 2973 4675
rect 2740 4644 2973 4672
rect 2740 4632 2746 4644
rect 2961 4641 2973 4644
rect 3007 4641 3019 4675
rect 2961 4635 3019 4641
rect 4525 4675 4583 4681
rect 4525 4641 4537 4675
rect 4571 4672 4583 4675
rect 5166 4672 5172 4684
rect 4571 4644 5172 4672
rect 4571 4641 4583 4644
rect 4525 4635 4583 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5442 4672 5448 4684
rect 5403 4644 5448 4672
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 6454 4672 6460 4684
rect 6415 4644 6460 4672
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 7101 4675 7159 4681
rect 7101 4672 7113 4675
rect 6972 4644 7113 4672
rect 6972 4632 6978 4644
rect 7101 4641 7113 4644
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 7368 4675 7426 4681
rect 7368 4641 7380 4675
rect 7414 4672 7426 4675
rect 8202 4672 8208 4684
rect 7414 4644 8208 4672
rect 7414 4641 7426 4644
rect 7368 4635 7426 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 10502 4672 10508 4684
rect 8803 4644 10508 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 11609 4675 11667 4681
rect 11609 4641 11621 4675
rect 11655 4672 11667 4675
rect 12434 4672 12440 4684
rect 11655 4644 12440 4672
rect 11655 4641 11667 4644
rect 11609 4635 11667 4641
rect 12434 4632 12440 4644
rect 12492 4632 12498 4684
rect 13808 4675 13866 4681
rect 13808 4672 13820 4675
rect 13004 4644 13820 4672
rect 1946 4564 1952 4616
rect 2004 4604 2010 4616
rect 3050 4604 3056 4616
rect 2004 4576 3056 4604
rect 2004 4564 2010 4576
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 5994 4604 6000 4616
rect 5767 4576 6000 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 2225 4539 2283 4545
rect 2225 4505 2237 4539
rect 2271 4536 2283 4539
rect 2409 4539 2467 4545
rect 2409 4536 2421 4539
rect 2271 4508 2421 4536
rect 2271 4505 2283 4508
rect 2225 4499 2283 4505
rect 2409 4505 2421 4508
rect 2455 4505 2467 4539
rect 2958 4536 2964 4548
rect 2409 4499 2467 4505
rect 2516 4508 2964 4536
rect 1673 4471 1731 4477
rect 1673 4437 1685 4471
rect 1719 4468 1731 4471
rect 2516 4468 2544 4508
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 3252 4536 3280 4567
rect 3326 4536 3332 4548
rect 3252 4508 3332 4536
rect 3326 4496 3332 4508
rect 3384 4536 3390 4548
rect 4632 4536 4660 4567
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6730 4604 6736 4616
rect 6691 4576 6736 4604
rect 6549 4567 6607 4573
rect 3384 4508 4660 4536
rect 5077 4539 5135 4545
rect 3384 4496 3390 4508
rect 5077 4505 5089 4539
rect 5123 4536 5135 4539
rect 6564 4536 6592 4567
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4604 11943 4607
rect 12158 4604 12164 4616
rect 11931 4576 12164 4604
rect 11931 4573 11943 4576
rect 11885 4567 11943 4573
rect 5123 4508 6592 4536
rect 5123 4505 5135 4508
rect 5077 4499 5135 4505
rect 1719 4440 2544 4468
rect 1719 4437 1731 4440
rect 1673 4431 1731 4437
rect 2590 4428 2596 4480
rect 2648 4468 2654 4480
rect 3418 4468 3424 4480
rect 2648 4440 3424 4468
rect 2648 4428 2654 4440
rect 3418 4428 3424 4440
rect 3476 4428 3482 4480
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 5684 4440 6101 4468
rect 5684 4428 5690 4440
rect 6089 4437 6101 4440
rect 6135 4437 6147 4471
rect 6089 4431 6147 4437
rect 9030 4428 9036 4480
rect 9088 4468 9094 4480
rect 9306 4468 9312 4480
rect 9088 4440 9312 4468
rect 9088 4428 9094 4440
rect 9306 4428 9312 4440
rect 9364 4468 9370 4480
rect 9784 4468 9812 4567
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 12802 4604 12808 4616
rect 12763 4576 12808 4604
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 13004 4613 13032 4644
rect 13808 4641 13820 4644
rect 13854 4672 13866 4675
rect 14274 4672 14280 4684
rect 13854 4644 14280 4672
rect 13854 4641 13866 4644
rect 13808 4635 13866 4641
rect 14274 4632 14280 4644
rect 14332 4632 14338 4684
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4573 13047 4607
rect 12989 4567 13047 4573
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4573 13599 4607
rect 15212 4604 15240 4712
rect 15304 4672 15332 4771
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 15749 4811 15807 4817
rect 15749 4808 15761 4811
rect 15436 4780 15761 4808
rect 15436 4768 15442 4780
rect 15749 4777 15761 4780
rect 15795 4777 15807 4811
rect 15749 4771 15807 4777
rect 15838 4768 15844 4820
rect 15896 4808 15902 4820
rect 17497 4811 17555 4817
rect 17497 4808 17509 4811
rect 15896 4780 17509 4808
rect 15896 4768 15902 4780
rect 17497 4777 17509 4780
rect 17543 4777 17555 4811
rect 17497 4771 17555 4777
rect 17589 4811 17647 4817
rect 17589 4777 17601 4811
rect 17635 4808 17647 4811
rect 17954 4808 17960 4820
rect 17635 4780 17960 4808
rect 17635 4777 17647 4780
rect 17589 4771 17647 4777
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 15657 4743 15715 4749
rect 15657 4709 15669 4743
rect 15703 4740 15715 4743
rect 16758 4740 16764 4752
rect 15703 4712 16764 4740
rect 15703 4709 15715 4712
rect 15657 4703 15715 4709
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 16301 4675 16359 4681
rect 16301 4672 16313 4675
rect 15304 4644 16313 4672
rect 16301 4641 16313 4644
rect 16347 4641 16359 4675
rect 16666 4672 16672 4684
rect 16301 4635 16359 4641
rect 16408 4644 16672 4672
rect 15838 4604 15844 4616
rect 15212 4576 15844 4604
rect 13541 4567 13599 4573
rect 10778 4496 10784 4548
rect 10836 4536 10842 4548
rect 10836 4508 11192 4536
rect 10836 4496 10842 4508
rect 11054 4468 11060 4480
rect 9364 4440 11060 4468
rect 9364 4428 9370 4440
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11164 4477 11192 4508
rect 11790 4496 11796 4548
rect 11848 4536 11854 4548
rect 12345 4539 12403 4545
rect 12345 4536 12357 4539
rect 11848 4508 12357 4536
rect 11848 4496 11854 4508
rect 12345 4505 12357 4508
rect 12391 4505 12403 4539
rect 13446 4536 13452 4548
rect 12345 4499 12403 4505
rect 12452 4508 13452 4536
rect 11149 4471 11207 4477
rect 11149 4437 11161 4471
rect 11195 4468 11207 4471
rect 12452 4468 12480 4508
rect 13446 4496 13452 4508
rect 13504 4496 13510 4548
rect 11195 4440 12480 4468
rect 11195 4437 11207 4440
rect 11149 4431 11207 4437
rect 12710 4428 12716 4480
rect 12768 4468 12774 4480
rect 13556 4468 13584 4567
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16408 4604 16436 4644
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 15979 4576 16436 4604
rect 16485 4607 16543 4613
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 16485 4573 16497 4607
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4573 17739 4607
rect 17681 4567 17739 4573
rect 15010 4496 15016 4548
rect 15068 4536 15074 4548
rect 16500 4536 16528 4567
rect 15068 4508 16528 4536
rect 15068 4496 15074 4508
rect 16850 4496 16856 4548
rect 16908 4536 16914 4548
rect 17402 4536 17408 4548
rect 16908 4508 17408 4536
rect 16908 4496 16914 4508
rect 17402 4496 17408 4508
rect 17460 4536 17466 4548
rect 17696 4536 17724 4567
rect 17460 4508 17724 4536
rect 17460 4496 17466 4508
rect 15102 4468 15108 4480
rect 12768 4440 15108 4468
rect 12768 4428 12774 4440
rect 15102 4428 15108 4440
rect 15160 4428 15166 4480
rect 17126 4468 17132 4480
rect 17087 4440 17132 4468
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 6178 4264 6184 4276
rect 3068 4236 6184 4264
rect 3068 4196 3096 4236
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 7558 4264 7564 4276
rect 7064 4236 7564 4264
rect 7064 4224 7070 4236
rect 7558 4224 7564 4236
rect 7616 4264 7622 4276
rect 8202 4264 8208 4276
rect 7616 4236 7880 4264
rect 8163 4236 8208 4264
rect 7616 4224 7622 4236
rect 2148 4168 3096 4196
rect 2148 4137 2176 4168
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 2222 4088 2228 4140
rect 2280 4128 2286 4140
rect 3068 4137 3096 4168
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 4764 4168 5396 4196
rect 4764 4156 4770 4168
rect 3053 4131 3111 4137
rect 2280 4100 2912 4128
rect 2280 4088 2286 4100
rect 1854 4060 1860 4072
rect 1815 4032 1860 4060
rect 1854 4020 1860 4032
rect 1912 4020 1918 4072
rect 2884 4069 2912 4100
rect 3053 4097 3065 4131
rect 3099 4097 3111 4131
rect 5368 4128 5396 4168
rect 5442 4156 5448 4208
rect 5500 4196 5506 4208
rect 5994 4196 6000 4208
rect 5500 4168 6000 4196
rect 5500 4156 5506 4168
rect 5828 4137 5856 4168
rect 5994 4156 6000 4168
rect 6052 4156 6058 4208
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 5368 4100 5641 4128
rect 3053 4091 3111 4097
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4097 5871 4131
rect 6196 4128 6224 4224
rect 6549 4199 6607 4205
rect 6549 4165 6561 4199
rect 6595 4196 6607 4199
rect 6638 4196 6644 4208
rect 6595 4168 6644 4196
rect 6595 4165 6607 4168
rect 6549 4159 6607 4165
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 7852 4128 7880 4236
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 8846 4224 8852 4276
rect 8904 4264 8910 4276
rect 12529 4267 12587 4273
rect 8904 4236 9527 4264
rect 8904 4224 8910 4236
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 6196 4100 6960 4128
rect 7852 4100 8493 4128
rect 5813 4091 5871 4097
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4029 3571 4063
rect 3513 4023 3571 4029
rect 3780 4063 3838 4069
rect 3780 4029 3792 4063
rect 3826 4060 3838 4063
rect 4798 4060 4804 4072
rect 3826 4032 4804 4060
rect 3826 4029 3838 4032
rect 3780 4023 3838 4029
rect 1394 3952 1400 4004
rect 1452 3992 1458 4004
rect 3528 3992 3556 4023
rect 4798 4020 4804 4032
rect 4856 4060 4862 4072
rect 5442 4060 5448 4072
rect 4856 4032 5448 4060
rect 4856 4020 4862 4032
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5994 4020 6000 4072
rect 6052 4060 6058 4072
rect 6181 4063 6239 4069
rect 6181 4060 6193 4063
rect 6052 4032 6193 4060
rect 6052 4020 6058 4032
rect 6181 4029 6193 4032
rect 6227 4060 6239 4063
rect 6549 4063 6607 4069
rect 6549 4060 6561 4063
rect 6227 4032 6561 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6549 4029 6561 4032
rect 6595 4029 6607 4063
rect 6822 4060 6828 4072
rect 6783 4032 6828 4060
rect 6549 4023 6607 4029
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 6932 4060 6960 4100
rect 8481 4097 8493 4100
rect 8527 4097 8539 4131
rect 9499 4128 9527 4236
rect 11256 4236 12020 4264
rect 10318 4196 10324 4208
rect 10279 4168 10324 4196
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 11256 4196 11284 4236
rect 11698 4196 11704 4208
rect 11072 4168 11284 4196
rect 11624 4168 11704 4196
rect 10226 4128 10232 4140
rect 9499 4100 10232 4128
rect 8481 4091 8539 4097
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 8737 4063 8795 4069
rect 8737 4060 8749 4063
rect 6932 4032 8749 4060
rect 8737 4029 8749 4032
rect 8783 4060 8795 4063
rect 10778 4060 10784 4072
rect 8783 4032 10784 4060
rect 8783 4029 8795 4032
rect 8737 4023 8795 4029
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 10870 4020 10876 4072
rect 10928 4060 10934 4072
rect 10980 4060 11008 4091
rect 10928 4032 11008 4060
rect 10928 4020 10934 4032
rect 6454 3992 6460 4004
rect 1452 3964 3556 3992
rect 5184 3964 6460 3992
rect 1452 3952 1458 3964
rect 1489 3927 1547 3933
rect 1489 3893 1501 3927
rect 1535 3924 1547 3927
rect 1762 3924 1768 3936
rect 1535 3896 1768 3924
rect 1535 3893 1547 3896
rect 1489 3887 1547 3893
rect 1762 3884 1768 3896
rect 1820 3884 1826 3936
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3924 2007 3927
rect 2406 3924 2412 3936
rect 1995 3896 2412 3924
rect 1995 3893 2007 3896
rect 1949 3887 2007 3893
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3924 2559 3927
rect 2774 3924 2780 3936
rect 2547 3896 2780 3924
rect 2547 3893 2559 3896
rect 2501 3887 2559 3893
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3924 3019 3927
rect 4706 3924 4712 3936
rect 3007 3896 4712 3924
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 4890 3924 4896 3936
rect 4851 3896 4896 3924
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5184 3933 5212 3964
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 6638 3952 6644 4004
rect 6696 3992 6702 4004
rect 7070 3995 7128 4001
rect 7070 3992 7082 3995
rect 6696 3964 7082 3992
rect 6696 3952 6702 3964
rect 7070 3961 7082 3964
rect 7116 3961 7128 3995
rect 7070 3955 7128 3961
rect 10502 3952 10508 4004
rect 10560 3992 10566 4004
rect 10689 3995 10747 4001
rect 10689 3992 10701 3995
rect 10560 3964 10701 3992
rect 10560 3952 10566 3964
rect 10689 3961 10701 3964
rect 10735 3992 10747 3995
rect 11072 3992 11100 4168
rect 11624 4060 11652 4168
rect 11698 4156 11704 4168
rect 11756 4156 11762 4208
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11848 4100 11897 4128
rect 11848 4088 11854 4100
rect 11885 4097 11897 4100
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11624 4032 11713 4060
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11992 4060 12020 4236
rect 12529 4233 12541 4267
rect 12575 4264 12587 4267
rect 12802 4264 12808 4276
rect 12575 4236 12808 4264
rect 12575 4233 12587 4236
rect 12529 4227 12587 4233
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 13998 4196 14004 4208
rect 13004 4168 14004 4196
rect 13004 4137 13032 4168
rect 13998 4156 14004 4168
rect 14056 4156 14062 4208
rect 14645 4199 14703 4205
rect 14645 4165 14657 4199
rect 14691 4165 14703 4199
rect 14645 4159 14703 4165
rect 12161 4131 12219 4137
rect 12161 4097 12173 4131
rect 12207 4128 12219 4131
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12207 4100 13001 4128
rect 12207 4097 12219 4100
rect 12161 4091 12219 4097
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 13170 4128 13176 4140
rect 13131 4100 13176 4128
rect 12989 4091 13047 4097
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 14274 4128 14280 4140
rect 14235 4100 14280 4128
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 14660 4128 14688 4159
rect 15102 4128 15108 4140
rect 14660 4100 15108 4128
rect 15102 4088 15108 4100
rect 15160 4128 15166 4140
rect 15197 4131 15255 4137
rect 15197 4128 15209 4131
rect 15160 4100 15209 4128
rect 15160 4088 15166 4100
rect 15197 4097 15209 4100
rect 15243 4097 15255 4131
rect 15197 4091 15255 4097
rect 17402 4088 17408 4140
rect 17460 4128 17466 4140
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 17460 4100 17509 4128
rect 17460 4088 17466 4100
rect 17497 4097 17509 4100
rect 17543 4097 17555 4131
rect 17497 4091 17555 4097
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 11992 4032 12909 4060
rect 11701 4023 11759 4029
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 14001 4063 14059 4069
rect 14001 4029 14013 4063
rect 14047 4060 14059 4063
rect 14550 4060 14556 4072
rect 14047 4032 14556 4060
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 15470 4069 15476 4072
rect 14829 4063 14887 4069
rect 14829 4029 14841 4063
rect 14875 4029 14887 4063
rect 15464 4060 15476 4069
rect 15383 4032 15476 4060
rect 14829 4023 14887 4029
rect 15464 4023 15476 4032
rect 15528 4060 15534 4072
rect 16482 4060 16488 4072
rect 15528 4032 16488 4060
rect 11793 3995 11851 4001
rect 10735 3964 11100 3992
rect 11256 3964 11744 3992
rect 10735 3961 10747 3964
rect 10689 3955 10747 3961
rect 5169 3927 5227 3933
rect 5169 3893 5181 3927
rect 5215 3893 5227 3927
rect 5534 3924 5540 3936
rect 5495 3896 5540 3924
rect 5169 3887 5227 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 5960 3896 6377 3924
rect 5960 3884 5966 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 8386 3884 8392 3936
rect 8444 3924 8450 3936
rect 9214 3924 9220 3936
rect 8444 3896 9220 3924
rect 8444 3884 8450 3896
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9548 3896 9873 3924
rect 9548 3884 9554 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 10781 3927 10839 3933
rect 10781 3924 10793 3927
rect 10284 3896 10793 3924
rect 10284 3884 10290 3896
rect 10781 3893 10793 3896
rect 10827 3924 10839 3927
rect 11256 3924 11284 3964
rect 10827 3896 11284 3924
rect 11333 3927 11391 3933
rect 10827 3893 10839 3896
rect 10781 3887 10839 3893
rect 11333 3893 11345 3927
rect 11379 3924 11391 3927
rect 11514 3924 11520 3936
rect 11379 3896 11520 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 11716 3924 11744 3964
rect 11793 3961 11805 3995
rect 11839 3992 11851 3995
rect 12250 3992 12256 4004
rect 11839 3964 12256 3992
rect 11839 3961 11851 3964
rect 11793 3955 11851 3961
rect 12250 3952 12256 3964
rect 12308 3952 12314 4004
rect 12526 3952 12532 4004
rect 12584 3992 12590 4004
rect 14844 3992 14872 4023
rect 15470 4020 15476 4023
rect 15528 4020 15534 4032
rect 16482 4020 16488 4032
rect 16540 4020 16546 4072
rect 17310 4020 17316 4072
rect 17368 4060 17374 4072
rect 17368 4032 17448 4060
rect 17368 4020 17374 4032
rect 12584 3964 14872 3992
rect 12584 3952 12590 3964
rect 14918 3952 14924 4004
rect 14976 3992 14982 4004
rect 17420 4001 17448 4032
rect 17954 4020 17960 4072
rect 18012 4060 18018 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 18012 4032 18061 4060
rect 18012 4020 18018 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 17405 3995 17463 4001
rect 14976 3964 17356 3992
rect 14976 3952 14982 3964
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 11716 3896 12173 3924
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 13630 3924 13636 3936
rect 13591 3896 13636 3924
rect 12161 3887 12219 3893
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 14093 3927 14151 3933
rect 14093 3893 14105 3927
rect 14139 3924 14151 3927
rect 14642 3924 14648 3936
rect 14139 3896 14648 3924
rect 14139 3893 14151 3896
rect 14093 3887 14151 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 16577 3927 16635 3933
rect 16577 3924 16589 3927
rect 14792 3896 16589 3924
rect 14792 3884 14798 3896
rect 16577 3893 16589 3896
rect 16623 3893 16635 3927
rect 16942 3924 16948 3936
rect 16903 3896 16948 3924
rect 16577 3887 16635 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17328 3933 17356 3964
rect 17405 3961 17417 3995
rect 17451 3961 17463 3995
rect 17405 3955 17463 3961
rect 17313 3927 17371 3933
rect 17313 3893 17325 3927
rect 17359 3893 17371 3927
rect 18230 3924 18236 3936
rect 18191 3896 18236 3924
rect 17313 3887 17371 3893
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 2777 3723 2835 3729
rect 2777 3720 2789 3723
rect 2556 3692 2789 3720
rect 2556 3680 2562 3692
rect 2777 3689 2789 3692
rect 2823 3689 2835 3723
rect 2777 3683 2835 3689
rect 4617 3723 4675 3729
rect 4617 3689 4629 3723
rect 4663 3720 4675 3723
rect 6270 3720 6276 3732
rect 4663 3692 6276 3720
rect 4663 3689 4675 3692
rect 4617 3683 4675 3689
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 6917 3723 6975 3729
rect 6917 3720 6929 3723
rect 6512 3692 6929 3720
rect 6512 3680 6518 3692
rect 6917 3689 6929 3692
rect 6963 3689 6975 3723
rect 7282 3720 7288 3732
rect 7243 3692 7288 3720
rect 6917 3683 6975 3689
rect 2406 3612 2412 3664
rect 2464 3652 2470 3664
rect 4709 3655 4767 3661
rect 4709 3652 4721 3655
rect 2464 3624 4721 3652
rect 2464 3612 2470 3624
rect 4709 3621 4721 3624
rect 4755 3621 4767 3655
rect 4709 3615 4767 3621
rect 4890 3612 4896 3664
rect 4948 3652 4954 3664
rect 5166 3652 5172 3664
rect 4948 3624 5172 3652
rect 4948 3612 4954 3624
rect 5166 3612 5172 3624
rect 5224 3652 5230 3664
rect 5528 3655 5586 3661
rect 5528 3652 5540 3655
rect 5224 3624 5540 3652
rect 5224 3612 5230 3624
rect 5528 3621 5540 3624
rect 5574 3652 5586 3655
rect 6730 3652 6736 3664
rect 5574 3624 6736 3652
rect 5574 3621 5586 3624
rect 5528 3615 5586 3621
rect 6730 3612 6736 3624
rect 6788 3612 6794 3664
rect 6932 3652 6960 3683
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 7926 3720 7932 3732
rect 7791 3692 7932 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 8662 3720 8668 3732
rect 8623 3692 8668 3720
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 8757 3723 8815 3729
rect 8757 3689 8769 3723
rect 8803 3720 8815 3723
rect 11422 3720 11428 3732
rect 8803 3692 11428 3720
rect 8803 3689 8815 3692
rect 8757 3683 8815 3689
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 12066 3720 12072 3732
rect 11532 3692 12072 3720
rect 7558 3652 7564 3664
rect 6932 3624 7564 3652
rect 7558 3612 7564 3624
rect 7616 3612 7622 3664
rect 11532 3652 11560 3692
rect 12066 3680 12072 3692
rect 12124 3720 12130 3732
rect 12526 3720 12532 3732
rect 12124 3692 12532 3720
rect 12124 3680 12130 3692
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 14274 3720 14280 3732
rect 12728 3692 13308 3720
rect 14235 3692 14280 3720
rect 9508 3624 11560 3652
rect 382 3544 388 3596
rect 440 3584 446 3596
rect 1653 3587 1711 3593
rect 1653 3584 1665 3587
rect 440 3556 1665 3584
rect 440 3544 446 3556
rect 1653 3553 1665 3556
rect 1699 3553 1711 3587
rect 1653 3547 1711 3553
rect 3237 3587 3295 3593
rect 3237 3553 3249 3587
rect 3283 3584 3295 3587
rect 4154 3584 4160 3596
rect 3283 3556 4160 3584
rect 3283 3553 3295 3556
rect 3237 3547 3295 3553
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 7101 3587 7159 3593
rect 5000 3556 6316 3584
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 3421 3519 3479 3525
rect 3421 3516 3433 3519
rect 3108 3488 3433 3516
rect 3108 3476 3114 3488
rect 3421 3485 3433 3488
rect 3467 3485 3479 3519
rect 4798 3516 4804 3528
rect 4759 3488 4804 3516
rect 3421 3479 3479 3485
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 3234 3408 3240 3460
rect 3292 3448 3298 3460
rect 5000 3448 5028 3556
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 5132 3488 5273 3516
rect 5132 3476 5138 3488
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 3292 3420 5028 3448
rect 6288 3448 6316 3556
rect 7101 3553 7113 3587
rect 7147 3584 7159 3587
rect 7374 3584 7380 3596
rect 7147 3556 7380 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 7653 3587 7711 3593
rect 7653 3553 7665 3587
rect 7699 3584 7711 3587
rect 8294 3584 8300 3596
rect 7699 3556 8300 3584
rect 7699 3553 7711 3556
rect 7653 3547 7711 3553
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 7668 3516 7696 3547
rect 8294 3544 8300 3556
rect 8352 3584 8358 3596
rect 9508 3593 9536 3624
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 12728 3652 12756 3692
rect 13170 3661 13176 3664
rect 11756 3624 12756 3652
rect 12805 3655 12863 3661
rect 11756 3612 11762 3624
rect 12805 3621 12817 3655
rect 12851 3652 12863 3655
rect 13164 3652 13176 3661
rect 12851 3624 13176 3652
rect 12851 3621 12863 3624
rect 12805 3615 12863 3621
rect 13164 3615 13176 3624
rect 13170 3612 13176 3615
rect 13228 3612 13234 3664
rect 13280 3652 13308 3692
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 14826 3680 14832 3732
rect 14884 3720 14890 3732
rect 16393 3723 16451 3729
rect 16393 3720 16405 3723
rect 14884 3692 16405 3720
rect 14884 3680 14890 3692
rect 16393 3689 16405 3692
rect 16439 3689 16451 3723
rect 16393 3683 16451 3689
rect 16485 3723 16543 3729
rect 16485 3689 16497 3723
rect 16531 3720 16543 3723
rect 17037 3723 17095 3729
rect 17037 3720 17049 3723
rect 16531 3692 17049 3720
rect 16531 3689 16543 3692
rect 16485 3683 16543 3689
rect 17037 3689 17049 3692
rect 17083 3689 17095 3723
rect 17037 3683 17095 3689
rect 17405 3723 17463 3729
rect 17405 3689 17417 3723
rect 17451 3720 17463 3723
rect 17770 3720 17776 3732
rect 17451 3692 17776 3720
rect 17451 3689 17463 3692
rect 17405 3683 17463 3689
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 18046 3680 18052 3732
rect 18104 3680 18110 3732
rect 18230 3720 18236 3732
rect 18191 3692 18236 3720
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 16666 3652 16672 3664
rect 13280 3624 16672 3652
rect 16666 3612 16672 3624
rect 16724 3612 16730 3664
rect 17497 3655 17555 3661
rect 17497 3621 17509 3655
rect 17543 3652 17555 3655
rect 18064 3652 18092 3680
rect 17543 3624 18092 3652
rect 17543 3621 17555 3624
rect 17497 3615 17555 3621
rect 9493 3587 9551 3593
rect 8352 3556 9076 3584
rect 8352 3544 8358 3556
rect 6512 3488 7696 3516
rect 7929 3519 7987 3525
rect 6512 3476 6518 3488
rect 7929 3485 7941 3519
rect 7975 3516 7987 3519
rect 8202 3516 8208 3528
rect 7975 3488 8208 3516
rect 7975 3485 7987 3488
rect 7929 3479 7987 3485
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8938 3516 8944 3528
rect 8536 3488 8944 3516
rect 8536 3476 8542 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 9048 3516 9076 3556
rect 9493 3553 9505 3587
rect 9539 3553 9551 3587
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9493 3547 9551 3553
rect 9674 3544 9680 3556
rect 9732 3584 9738 3596
rect 10597 3587 10655 3593
rect 10597 3584 10609 3587
rect 9732 3556 10609 3584
rect 9732 3544 9738 3556
rect 10597 3553 10609 3556
rect 10643 3553 10655 3587
rect 10597 3547 10655 3553
rect 10689 3587 10747 3593
rect 10689 3553 10701 3587
rect 10735 3584 10747 3587
rect 10778 3584 10784 3596
rect 10735 3556 10784 3584
rect 10735 3553 10747 3556
rect 10689 3547 10747 3553
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 11241 3587 11299 3593
rect 11241 3584 11253 3587
rect 11204 3556 11253 3584
rect 11204 3544 11210 3556
rect 11241 3553 11253 3556
rect 11287 3553 11299 3587
rect 11241 3547 11299 3553
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 11497 3587 11555 3593
rect 11497 3584 11509 3587
rect 11388 3556 11509 3584
rect 11388 3544 11394 3556
rect 11497 3553 11509 3556
rect 11543 3553 11555 3587
rect 11497 3547 11555 3553
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 13596 3556 15301 3584
rect 13596 3544 13602 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 15289 3547 15347 3553
rect 15387 3556 18061 3584
rect 10502 3516 10508 3528
rect 9048 3488 10508 3516
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 10870 3516 10876 3528
rect 10831 3488 10876 3516
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 12710 3476 12716 3528
rect 12768 3516 12774 3528
rect 12897 3519 12955 3525
rect 12897 3516 12909 3519
rect 12768 3488 12909 3516
rect 12768 3476 12774 3488
rect 12897 3485 12909 3488
rect 12943 3485 12955 3519
rect 12897 3479 12955 3485
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 15387 3516 15415 3556
rect 18049 3553 18061 3556
rect 18095 3553 18107 3587
rect 18049 3547 18107 3553
rect 14056 3488 15415 3516
rect 15473 3519 15531 3525
rect 14056 3476 14062 3488
rect 15473 3485 15485 3519
rect 15519 3485 15531 3519
rect 15473 3479 15531 3485
rect 9861 3451 9919 3457
rect 9861 3448 9873 3451
rect 6288 3420 9873 3448
rect 3292 3408 3298 3420
rect 9861 3417 9873 3420
rect 9907 3417 9919 3451
rect 10226 3448 10232 3460
rect 10187 3420 10232 3448
rect 9861 3411 9919 3417
rect 10226 3408 10232 3420
rect 10284 3408 10290 3460
rect 12621 3451 12679 3457
rect 12621 3417 12633 3451
rect 12667 3448 12679 3451
rect 12805 3451 12863 3457
rect 12805 3448 12817 3451
rect 12667 3420 12817 3448
rect 12667 3417 12679 3420
rect 12621 3411 12679 3417
rect 12805 3417 12817 3420
rect 12851 3417 12863 3451
rect 12805 3411 12863 3417
rect 14090 3408 14096 3460
rect 14148 3448 14154 3460
rect 14918 3448 14924 3460
rect 14148 3420 14924 3448
rect 14148 3408 14154 3420
rect 14918 3408 14924 3420
rect 14976 3408 14982 3460
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 3326 3380 3332 3392
rect 1820 3352 3332 3380
rect 1820 3340 1826 3352
rect 3326 3340 3332 3352
rect 3384 3340 3390 3392
rect 4249 3383 4307 3389
rect 4249 3349 4261 3383
rect 4295 3380 4307 3383
rect 4890 3380 4896 3392
rect 4295 3352 4896 3380
rect 4295 3349 4307 3352
rect 4249 3343 4307 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 6638 3380 6644 3392
rect 5500 3352 6644 3380
rect 5500 3340 5506 3352
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 8294 3380 8300 3392
rect 8255 3352 8300 3380
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 9306 3380 9312 3392
rect 9267 3352 9312 3380
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 12894 3380 12900 3392
rect 9640 3352 12900 3380
rect 9640 3340 9646 3352
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13170 3340 13176 3392
rect 13228 3380 13234 3392
rect 15488 3380 15516 3479
rect 15654 3476 15660 3528
rect 15712 3516 15718 3528
rect 16298 3516 16304 3528
rect 15712 3488 16304 3516
rect 15712 3476 15718 3488
rect 16298 3476 16304 3488
rect 16356 3516 16362 3528
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 16356 3488 16589 3516
rect 16356 3476 16362 3488
rect 16577 3485 16589 3488
rect 16623 3485 16635 3519
rect 16577 3479 16635 3485
rect 17589 3519 17647 3525
rect 17589 3485 17601 3519
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 17402 3408 17408 3460
rect 17460 3448 17466 3460
rect 17604 3448 17632 3479
rect 17460 3420 17632 3448
rect 17460 3408 17466 3420
rect 13228 3352 15516 3380
rect 16025 3383 16083 3389
rect 13228 3340 13234 3352
rect 16025 3349 16037 3383
rect 16071 3380 16083 3383
rect 16850 3380 16856 3392
rect 16071 3352 16856 3380
rect 16071 3349 16083 3352
rect 16025 3343 16083 3349
rect 16850 3340 16856 3352
rect 16908 3340 16914 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 3252 3148 6040 3176
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 3252 3040 3280 3148
rect 5718 3108 5724 3120
rect 3344 3080 5724 3108
rect 3344 3049 3372 3080
rect 5718 3068 5724 3080
rect 5776 3068 5782 3120
rect 6012 3108 6040 3148
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 7892 3148 8125 3176
rect 7892 3136 7898 3148
rect 8113 3145 8125 3148
rect 8159 3145 8171 3179
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 8113 3139 8171 3145
rect 8220 3148 10609 3176
rect 8220 3108 8248 3148
rect 10597 3145 10609 3148
rect 10643 3176 10655 3179
rect 11330 3176 11336 3188
rect 10643 3148 11336 3176
rect 10643 3145 10655 3148
rect 10597 3139 10655 3145
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 12032 3148 12449 3176
rect 12032 3136 12038 3148
rect 12437 3145 12449 3148
rect 12483 3145 12495 3179
rect 12437 3139 12495 3145
rect 13725 3179 13783 3185
rect 13725 3145 13737 3179
rect 13771 3176 13783 3179
rect 16390 3176 16396 3188
rect 13771 3148 16396 3176
rect 13771 3145 13783 3148
rect 13725 3139 13783 3145
rect 16390 3136 16396 3148
rect 16448 3136 16454 3188
rect 11790 3108 11796 3120
rect 6012 3080 8248 3108
rect 11440 3080 11796 3108
rect 2547 3012 3280 3040
rect 3329 3043 3387 3049
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 3329 3009 3341 3043
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 3970 3040 3976 3052
rect 3559 3012 3976 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 3970 3000 3976 3012
rect 4028 3040 4034 3052
rect 4430 3040 4436 3052
rect 4028 3012 4436 3040
rect 4028 3000 4034 3012
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3040 4583 3043
rect 5442 3040 5448 3052
rect 4571 3012 5448 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 7653 3043 7711 3049
rect 5592 3012 5637 3040
rect 5592 3000 5598 3012
rect 7653 3009 7665 3043
rect 7699 3009 7711 3043
rect 7653 3003 7711 3009
rect 1210 2932 1216 2984
rect 1268 2972 1274 2984
rect 4062 2972 4068 2984
rect 1268 2944 4068 2972
rect 1268 2932 1274 2944
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 4341 2975 4399 2981
rect 4341 2941 4353 2975
rect 4387 2972 4399 2975
rect 5626 2972 5632 2984
rect 4387 2944 5632 2972
rect 4387 2941 4399 2944
rect 4341 2935 4399 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 5997 2975 6055 2981
rect 5997 2941 6009 2975
rect 6043 2972 6055 2975
rect 6546 2972 6552 2984
rect 6043 2944 6552 2972
rect 6043 2941 6055 2944
rect 5997 2935 6055 2941
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 7668 2972 7696 3003
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 7800 3012 8677 3040
rect 7800 3000 7806 3012
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 11440 3049 11468 3080
rect 11790 3068 11796 3080
rect 11848 3068 11854 3120
rect 16316 3080 17356 3108
rect 16316 3052 16344 3080
rect 11425 3043 11483 3049
rect 11425 3040 11437 3043
rect 10744 3012 11437 3040
rect 10744 3000 10750 3012
rect 11425 3009 11437 3012
rect 11471 3009 11483 3043
rect 11425 3003 11483 3009
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 11664 3012 13001 3040
rect 11664 3000 11670 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3040 14427 3043
rect 14734 3040 14740 3052
rect 14415 3012 14740 3040
rect 14415 3009 14427 3012
rect 14369 3003 14427 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 15470 3040 15476 3052
rect 15427 3012 15476 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 16298 3040 16304 3052
rect 16259 3012 16304 3040
rect 16298 3000 16304 3012
rect 16356 3000 16362 3052
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 17328 3049 17356 3080
rect 17221 3043 17279 3049
rect 17221 3040 17233 3043
rect 17184 3012 17233 3040
rect 17184 3000 17190 3012
rect 17221 3009 17233 3012
rect 17267 3009 17279 3043
rect 17221 3003 17279 3009
rect 17313 3043 17371 3049
rect 17313 3009 17325 3043
rect 17359 3009 17371 3043
rect 17313 3003 17371 3009
rect 8478 2972 8484 2984
rect 7668 2944 8484 2972
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8573 2975 8631 2981
rect 8573 2941 8585 2975
rect 8619 2972 8631 2975
rect 8754 2972 8760 2984
rect 8619 2944 8760 2972
rect 8619 2941 8631 2944
rect 8573 2935 8631 2941
rect 8754 2932 8760 2944
rect 8812 2932 8818 2984
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9306 2972 9312 2984
rect 9263 2944 9312 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 11146 2972 11152 2984
rect 9416 2944 11152 2972
rect 2225 2907 2283 2913
rect 2225 2873 2237 2907
rect 2271 2904 2283 2907
rect 2958 2904 2964 2916
rect 2271 2876 2964 2904
rect 2271 2873 2283 2876
rect 2225 2867 2283 2873
rect 2958 2864 2964 2876
rect 3016 2864 3022 2916
rect 3237 2907 3295 2913
rect 3237 2873 3249 2907
rect 3283 2904 3295 2907
rect 3510 2904 3516 2916
rect 3283 2876 3516 2904
rect 3283 2873 3295 2876
rect 3237 2867 3295 2873
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 3786 2864 3792 2916
rect 3844 2904 3850 2916
rect 6273 2907 6331 2913
rect 6273 2904 6285 2907
rect 3844 2876 6285 2904
rect 3844 2864 3850 2876
rect 6273 2873 6285 2876
rect 6319 2873 6331 2907
rect 6273 2867 6331 2873
rect 6362 2864 6368 2916
rect 6420 2904 6426 2916
rect 7469 2907 7527 2913
rect 6420 2876 6776 2904
rect 6420 2864 6426 2876
rect 6748 2848 6776 2876
rect 7469 2873 7481 2907
rect 7515 2904 7527 2907
rect 9416 2904 9444 2944
rect 11146 2932 11152 2944
rect 11204 2972 11210 2984
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 11204 2944 11253 2972
rect 11204 2932 11210 2944
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 12434 2972 12440 2984
rect 11572 2944 12440 2972
rect 11572 2932 11578 2944
rect 12434 2932 12440 2944
rect 12492 2932 12498 2984
rect 12894 2972 12900 2984
rect 12855 2944 12900 2972
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2972 14243 2975
rect 15746 2972 15752 2984
rect 14231 2944 15752 2972
rect 14231 2941 14243 2944
rect 14185 2935 14243 2941
rect 15746 2932 15752 2944
rect 15804 2932 15810 2984
rect 16114 2972 16120 2984
rect 16075 2944 16120 2972
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 16209 2975 16267 2981
rect 16209 2941 16221 2975
rect 16255 2972 16267 2975
rect 16574 2972 16580 2984
rect 16255 2944 16580 2972
rect 16255 2941 16267 2944
rect 16209 2935 16267 2941
rect 16574 2932 16580 2944
rect 16632 2932 16638 2984
rect 9490 2913 9496 2916
rect 7515 2876 9444 2904
rect 7515 2873 7527 2876
rect 7469 2867 7527 2873
rect 9484 2867 9496 2913
rect 9548 2904 9554 2916
rect 9548 2876 9584 2904
rect 9490 2864 9496 2867
rect 9548 2864 9554 2876
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 12805 2907 12863 2913
rect 12805 2904 12817 2907
rect 9732 2876 12817 2904
rect 9732 2864 9738 2876
rect 12805 2873 12817 2876
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 14093 2907 14151 2913
rect 14093 2873 14105 2907
rect 14139 2904 14151 2907
rect 15105 2907 15163 2913
rect 14139 2876 14780 2904
rect 14139 2873 14151 2876
rect 14093 2867 14151 2873
rect 1854 2836 1860 2848
rect 1815 2808 1860 2836
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 2317 2839 2375 2845
rect 2317 2805 2329 2839
rect 2363 2836 2375 2839
rect 2869 2839 2927 2845
rect 2869 2836 2881 2839
rect 2363 2808 2881 2836
rect 2363 2805 2375 2808
rect 2317 2799 2375 2805
rect 2869 2805 2881 2808
rect 2915 2805 2927 2839
rect 2869 2799 2927 2805
rect 3881 2839 3939 2845
rect 3881 2805 3893 2839
rect 3927 2836 3939 2839
rect 4062 2836 4068 2848
rect 3927 2808 4068 2836
rect 3927 2805 3939 2808
rect 3881 2799 3939 2805
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 4246 2836 4252 2848
rect 4207 2808 4252 2836
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 4982 2836 4988 2848
rect 4943 2808 4988 2836
rect 4982 2796 4988 2808
rect 5040 2796 5046 2848
rect 5074 2796 5080 2848
rect 5132 2836 5138 2848
rect 5353 2839 5411 2845
rect 5353 2836 5365 2839
rect 5132 2808 5365 2836
rect 5132 2796 5138 2808
rect 5353 2805 5365 2808
rect 5399 2805 5411 2839
rect 5353 2799 5411 2805
rect 5445 2839 5503 2845
rect 5445 2805 5457 2839
rect 5491 2836 5503 2839
rect 5994 2836 6000 2848
rect 5491 2808 6000 2836
rect 5491 2805 5503 2808
rect 5445 2799 5503 2805
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 6730 2796 6736 2848
rect 6788 2796 6794 2848
rect 7101 2839 7159 2845
rect 7101 2805 7113 2839
rect 7147 2836 7159 2839
rect 7374 2836 7380 2848
rect 7147 2808 7380 2836
rect 7147 2805 7159 2808
rect 7101 2799 7159 2805
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 7561 2839 7619 2845
rect 7561 2805 7573 2839
rect 7607 2836 7619 2839
rect 8110 2836 8116 2848
rect 7607 2808 8116 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 8478 2836 8484 2848
rect 8439 2808 8484 2836
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 10870 2836 10876 2848
rect 10831 2808 10876 2836
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 11333 2839 11391 2845
rect 11333 2805 11345 2839
rect 11379 2836 11391 2839
rect 11882 2836 11888 2848
rect 11379 2808 11888 2836
rect 11379 2805 11391 2808
rect 11333 2799 11391 2805
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 12710 2796 12716 2848
rect 12768 2836 12774 2848
rect 13814 2836 13820 2848
rect 12768 2808 13820 2836
rect 12768 2796 12774 2808
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 13998 2796 14004 2848
rect 14056 2836 14062 2848
rect 14366 2836 14372 2848
rect 14056 2808 14372 2836
rect 14056 2796 14062 2808
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 14752 2845 14780 2876
rect 15105 2873 15117 2907
rect 15151 2904 15163 2907
rect 15654 2904 15660 2916
rect 15151 2876 15660 2904
rect 15151 2873 15163 2876
rect 15105 2867 15163 2873
rect 15654 2864 15660 2876
rect 15712 2864 15718 2916
rect 16942 2864 16948 2916
rect 17000 2904 17006 2916
rect 17129 2907 17187 2913
rect 17129 2904 17141 2907
rect 17000 2876 17141 2904
rect 17000 2864 17006 2876
rect 17129 2873 17141 2876
rect 17175 2873 17187 2907
rect 17129 2867 17187 2873
rect 14737 2839 14795 2845
rect 14737 2805 14749 2839
rect 14783 2805 14795 2839
rect 14737 2799 14795 2805
rect 15197 2839 15255 2845
rect 15197 2805 15209 2839
rect 15243 2836 15255 2839
rect 15749 2839 15807 2845
rect 15749 2836 15761 2839
rect 15243 2808 15761 2836
rect 15243 2805 15255 2808
rect 15197 2799 15255 2805
rect 15749 2805 15761 2808
rect 15795 2805 15807 2839
rect 16758 2836 16764 2848
rect 16719 2808 16764 2836
rect 15749 2799 15807 2805
rect 16758 2796 16764 2808
rect 16816 2796 16822 2848
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 2958 2632 2964 2644
rect 2919 2604 2964 2632
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 4246 2592 4252 2644
rect 4304 2632 4310 2644
rect 4525 2635 4583 2641
rect 4525 2632 4537 2635
rect 4304 2604 4537 2632
rect 4304 2592 4310 2604
rect 4525 2601 4537 2604
rect 4571 2601 4583 2635
rect 4982 2632 4988 2644
rect 4943 2604 4988 2632
rect 4525 2595 4583 2601
rect 4982 2592 4988 2604
rect 5040 2592 5046 2644
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 5813 2635 5871 2641
rect 5813 2632 5825 2635
rect 5776 2604 5825 2632
rect 5776 2592 5782 2604
rect 5813 2601 5825 2604
rect 5859 2601 5871 2635
rect 7374 2632 7380 2644
rect 7335 2604 7380 2632
rect 5813 2595 5871 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 9674 2632 9680 2644
rect 8711 2604 9680 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 9766 2592 9772 2644
rect 9824 2632 9830 2644
rect 9861 2635 9919 2641
rect 9861 2632 9873 2635
rect 9824 2604 9873 2632
rect 9824 2592 9830 2604
rect 9861 2601 9873 2604
rect 9907 2601 9919 2635
rect 9861 2595 9919 2601
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10321 2635 10379 2641
rect 10321 2632 10333 2635
rect 10284 2604 10333 2632
rect 10284 2592 10290 2604
rect 10321 2601 10333 2604
rect 10367 2601 10379 2635
rect 10321 2595 10379 2601
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 11241 2635 11299 2641
rect 11241 2632 11253 2635
rect 11020 2604 11253 2632
rect 11020 2592 11026 2604
rect 11241 2601 11253 2604
rect 11287 2601 11299 2635
rect 11241 2595 11299 2601
rect 11333 2635 11391 2641
rect 11333 2601 11345 2635
rect 11379 2632 11391 2635
rect 11422 2632 11428 2644
rect 11379 2604 11428 2632
rect 11379 2601 11391 2604
rect 11333 2595 11391 2601
rect 11422 2592 11428 2604
rect 11480 2632 11486 2644
rect 12250 2632 12256 2644
rect 11480 2604 12256 2632
rect 11480 2592 11486 2604
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 12989 2635 13047 2641
rect 12989 2601 13001 2635
rect 13035 2632 13047 2635
rect 13449 2635 13507 2641
rect 13449 2632 13461 2635
rect 13035 2604 13461 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 13449 2601 13461 2604
rect 13495 2601 13507 2635
rect 13630 2632 13636 2644
rect 13591 2604 13636 2632
rect 13449 2595 13507 2601
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 13722 2592 13728 2644
rect 13780 2632 13786 2644
rect 14001 2635 14059 2641
rect 14001 2632 14013 2635
rect 13780 2604 14013 2632
rect 13780 2592 13786 2604
rect 14001 2601 14013 2604
rect 14047 2601 14059 2635
rect 15654 2632 15660 2644
rect 15615 2604 15660 2632
rect 14001 2595 14059 2601
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 15746 2592 15752 2644
rect 15804 2632 15810 2644
rect 16669 2635 16727 2641
rect 16669 2632 16681 2635
rect 15804 2604 16681 2632
rect 15804 2592 15810 2604
rect 16669 2601 16681 2604
rect 16715 2601 16727 2635
rect 16669 2595 16727 2601
rect 16758 2592 16764 2644
rect 16816 2632 16822 2644
rect 17129 2635 17187 2641
rect 17129 2632 17141 2635
rect 16816 2604 17141 2632
rect 16816 2592 16822 2604
rect 17129 2601 17141 2604
rect 17175 2601 17187 2635
rect 17129 2595 17187 2601
rect 2682 2564 2688 2576
rect 1412 2536 2688 2564
rect 1412 2505 1440 2536
rect 2682 2524 2688 2536
rect 2740 2524 2746 2576
rect 2774 2524 2780 2576
rect 2832 2564 2838 2576
rect 3421 2567 3479 2573
rect 3421 2564 3433 2567
rect 2832 2536 3433 2564
rect 2832 2524 2838 2536
rect 3421 2533 3433 2536
rect 3467 2533 3479 2567
rect 4890 2564 4896 2576
rect 4851 2536 4896 2564
rect 3421 2527 3479 2533
rect 4890 2524 4896 2536
rect 4948 2524 4954 2576
rect 5074 2524 5080 2576
rect 5132 2564 5138 2576
rect 8205 2567 8263 2573
rect 8205 2564 8217 2567
rect 5132 2536 8217 2564
rect 5132 2524 5138 2536
rect 8205 2533 8217 2536
rect 8251 2533 8263 2567
rect 8205 2527 8263 2533
rect 9125 2567 9183 2573
rect 9125 2533 9137 2567
rect 9171 2564 9183 2567
rect 10870 2564 10876 2576
rect 9171 2536 10876 2564
rect 9171 2533 9183 2536
rect 9125 2527 9183 2533
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 13814 2524 13820 2576
rect 13872 2564 13878 2576
rect 14921 2567 14979 2573
rect 14921 2564 14933 2567
rect 13872 2536 14933 2564
rect 13872 2524 13878 2536
rect 14921 2533 14933 2536
rect 14967 2533 14979 2567
rect 14921 2527 14979 2533
rect 15562 2524 15568 2576
rect 15620 2564 15626 2576
rect 16025 2567 16083 2573
rect 16025 2564 16037 2567
rect 15620 2536 16037 2564
rect 15620 2524 15626 2536
rect 16025 2533 16037 2536
rect 16071 2533 16083 2567
rect 16025 2527 16083 2533
rect 16114 2524 16120 2576
rect 16172 2564 16178 2576
rect 16172 2536 16217 2564
rect 16172 2524 16178 2536
rect 16850 2524 16856 2576
rect 16908 2564 16914 2576
rect 17037 2567 17095 2573
rect 17037 2564 17049 2567
rect 16908 2536 17049 2564
rect 16908 2524 16914 2536
rect 17037 2533 17049 2536
rect 17083 2533 17095 2567
rect 17037 2527 17095 2533
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 3602 2496 3608 2508
rect 1995 2468 3608 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 3602 2456 3608 2468
rect 3660 2456 3666 2508
rect 5350 2456 5356 2508
rect 5408 2496 5414 2508
rect 6181 2499 6239 2505
rect 6181 2496 6193 2499
rect 5408 2468 6193 2496
rect 5408 2456 5414 2468
rect 6181 2465 6193 2468
rect 6227 2465 6239 2499
rect 6181 2459 6239 2465
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 7926 2496 7932 2508
rect 7331 2468 7696 2496
rect 7887 2468 7932 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 2130 2428 2136 2440
rect 2091 2400 2136 2428
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 3970 2428 3976 2440
rect 3559 2400 3976 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 5166 2428 5172 2440
rect 5127 2400 5172 2428
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 6273 2431 6331 2437
rect 6273 2397 6285 2431
rect 6319 2397 6331 2431
rect 6273 2391 6331 2397
rect 6288 2360 6316 2391
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 7466 2428 7472 2440
rect 6420 2400 6465 2428
rect 7427 2400 7472 2428
rect 6420 2388 6426 2400
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 7668 2428 7696 2468
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 9033 2499 9091 2505
rect 9033 2465 9045 2499
rect 9079 2496 9091 2499
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9079 2468 9781 2496
rect 9079 2465 9091 2468
rect 9033 2459 9091 2465
rect 9769 2465 9781 2468
rect 9815 2465 9827 2499
rect 9769 2459 9827 2465
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2496 10287 2499
rect 11698 2496 11704 2508
rect 10275 2468 11704 2496
rect 10275 2465 10287 2468
rect 10229 2459 10287 2465
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 13446 2456 13452 2508
rect 13504 2496 13510 2508
rect 14645 2499 14703 2505
rect 13504 2468 14228 2496
rect 13504 2456 13510 2468
rect 8294 2428 8300 2440
rect 7668 2400 8300 2428
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 10134 2428 10140 2440
rect 9355 2400 10140 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 10686 2428 10692 2440
rect 10551 2400 10692 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 10686 2388 10692 2400
rect 10744 2428 10750 2440
rect 11425 2431 11483 2437
rect 11425 2428 11437 2431
rect 10744 2400 11437 2428
rect 10744 2388 10750 2400
rect 11425 2397 11437 2400
rect 11471 2397 11483 2431
rect 11425 2391 11483 2397
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 13078 2428 13084 2440
rect 12400 2400 12756 2428
rect 13039 2400 13084 2428
rect 12400 2388 12406 2400
rect 12621 2363 12679 2369
rect 12621 2360 12633 2363
rect 6288 2332 12633 2360
rect 12621 2329 12633 2332
rect 12667 2329 12679 2363
rect 12728 2360 12756 2400
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 13262 2428 13268 2440
rect 13223 2400 13268 2428
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 14200 2437 14228 2468
rect 14645 2465 14657 2499
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 14185 2431 14243 2437
rect 14185 2397 14197 2431
rect 14231 2397 14243 2431
rect 14185 2391 14243 2397
rect 14660 2360 14688 2459
rect 15470 2456 15476 2508
rect 15528 2496 15534 2508
rect 15528 2468 17264 2496
rect 15528 2456 15534 2468
rect 16298 2428 16304 2440
rect 16259 2400 16304 2428
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 17236 2437 17264 2468
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2397 17279 2431
rect 17221 2391 17279 2397
rect 12728 2332 14688 2360
rect 12621 2323 12679 2329
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2292 1639 2295
rect 2774 2292 2780 2304
rect 1627 2264 2780 2292
rect 1627 2261 1639 2264
rect 1581 2255 1639 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 6917 2295 6975 2301
rect 6917 2261 6929 2295
rect 6963 2292 6975 2295
rect 8478 2292 8484 2304
rect 6963 2264 8484 2292
rect 6963 2261 6975 2264
rect 6917 2255 6975 2261
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 9769 2295 9827 2301
rect 9769 2261 9781 2295
rect 9815 2292 9827 2295
rect 10873 2295 10931 2301
rect 10873 2292 10885 2295
rect 9815 2264 10885 2292
rect 9815 2261 9827 2264
rect 9769 2255 9827 2261
rect 10873 2261 10885 2264
rect 10919 2261 10931 2295
rect 10873 2255 10931 2261
rect 13449 2295 13507 2301
rect 13449 2261 13461 2295
rect 13495 2292 13507 2295
rect 13998 2292 14004 2304
rect 13495 2264 14004 2292
rect 13495 2261 13507 2264
rect 13449 2255 13507 2261
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 13078 2048 13084 2100
rect 13136 2088 13142 2100
rect 14182 2088 14188 2100
rect 13136 2060 14188 2088
rect 13136 2048 13142 2060
rect 14182 2048 14188 2060
rect 14240 2048 14246 2100
rect 3234 1844 3240 1896
rect 3292 1884 3298 1896
rect 5902 1884 5908 1896
rect 3292 1856 5908 1884
rect 3292 1844 3298 1856
rect 5902 1844 5908 1856
rect 5960 1844 5966 1896
rect 2038 1300 2044 1352
rect 2096 1340 2102 1352
rect 15194 1340 15200 1352
rect 2096 1312 15200 1340
rect 2096 1300 2102 1312
rect 15194 1300 15200 1312
rect 15252 1300 15258 1352
<< via1 >>
rect 4068 15240 4120 15292
rect 10508 15240 10560 15292
rect 3976 15172 4028 15224
rect 15016 15172 15068 15224
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 1584 14560 1636 14612
rect 16948 14492 17000 14544
rect 2964 14424 3016 14476
rect 7748 14424 7800 14476
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 5908 14016 5960 14068
rect 1952 13948 2004 14000
rect 9772 13948 9824 14000
rect 1676 13880 1728 13932
rect 2780 13880 2832 13932
rect 10232 13880 10284 13932
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 2872 13812 2924 13864
rect 6092 13855 6144 13864
rect 6092 13821 6101 13855
rect 6101 13821 6135 13855
rect 6135 13821 6144 13855
rect 6092 13812 6144 13821
rect 3240 13744 3292 13796
rect 10508 13812 10560 13864
rect 16396 14016 16448 14068
rect 13912 13948 13964 14000
rect 17592 13948 17644 14000
rect 17868 13880 17920 13932
rect 9496 13676 9548 13728
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 9772 13676 9824 13685
rect 11520 13744 11572 13796
rect 16212 13676 16264 13728
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 1492 13472 1544 13524
rect 15568 13472 15620 13524
rect 2872 13404 2924 13456
rect 12440 13404 12492 13456
rect 2780 13336 2832 13388
rect 10324 13379 10376 13388
rect 10324 13345 10333 13379
rect 10333 13345 10367 13379
rect 10367 13345 10376 13379
rect 10324 13336 10376 13345
rect 11244 13336 11296 13388
rect 12624 13336 12676 13388
rect 16948 13379 17000 13388
rect 16948 13345 16957 13379
rect 16957 13345 16991 13379
rect 16991 13345 17000 13379
rect 16948 13336 17000 13345
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2044 13268 2096 13277
rect 10508 13311 10560 13320
rect 10508 13277 10517 13311
rect 10517 13277 10551 13311
rect 10551 13277 10560 13311
rect 10508 13268 10560 13277
rect 10784 13268 10836 13320
rect 17224 13311 17276 13320
rect 17224 13277 17233 13311
rect 17233 13277 17267 13311
rect 17267 13277 17276 13311
rect 17224 13268 17276 13277
rect 2780 13243 2832 13252
rect 2780 13209 2789 13243
rect 2789 13209 2823 13243
rect 2823 13209 2832 13243
rect 2780 13200 2832 13209
rect 7104 13200 7156 13252
rect 10416 13200 10468 13252
rect 10600 13200 10652 13252
rect 18512 13268 18564 13320
rect 3792 13132 3844 13184
rect 8852 13132 8904 13184
rect 8944 13132 8996 13184
rect 11612 13132 11664 13184
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 8392 12928 8444 12980
rect 10324 12928 10376 12980
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 3332 12792 3384 12844
rect 7196 12792 7248 12844
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 8760 12860 8812 12912
rect 8852 12860 8904 12912
rect 13268 12860 13320 12912
rect 1492 12724 1544 12776
rect 7932 12724 7984 12776
rect 8116 12792 8168 12844
rect 10600 12792 10652 12844
rect 10876 12792 10928 12844
rect 12256 12792 12308 12844
rect 8484 12724 8536 12776
rect 11428 12724 11480 12776
rect 17776 12928 17828 12980
rect 14924 12860 14976 12912
rect 16948 12792 17000 12844
rect 14280 12724 14332 12776
rect 7104 12656 7156 12708
rect 11060 12656 11112 12708
rect 15752 12656 15804 12708
rect 7840 12588 7892 12640
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 9036 12588 9088 12640
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 9680 12631 9732 12640
rect 9680 12597 9689 12631
rect 9689 12597 9723 12631
rect 9723 12597 9732 12631
rect 9680 12588 9732 12597
rect 10692 12631 10744 12640
rect 10692 12597 10701 12631
rect 10701 12597 10735 12631
rect 10735 12597 10744 12631
rect 10692 12588 10744 12597
rect 11152 12588 11204 12640
rect 11704 12631 11756 12640
rect 11704 12597 11713 12631
rect 11713 12597 11747 12631
rect 11747 12597 11756 12631
rect 11704 12588 11756 12597
rect 12532 12588 12584 12640
rect 15200 12588 15252 12640
rect 17040 12631 17092 12640
rect 17040 12597 17049 12631
rect 17049 12597 17083 12631
rect 17083 12597 17092 12631
rect 17040 12588 17092 12597
rect 17132 12631 17184 12640
rect 17132 12597 17141 12631
rect 17141 12597 17175 12631
rect 17175 12597 17184 12631
rect 18236 12631 18288 12640
rect 17132 12588 17184 12597
rect 18236 12597 18245 12631
rect 18245 12597 18279 12631
rect 18279 12597 18288 12631
rect 18236 12588 18288 12597
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 7288 12384 7340 12436
rect 8944 12427 8996 12436
rect 8944 12393 8953 12427
rect 8953 12393 8987 12427
rect 8987 12393 8996 12427
rect 8944 12384 8996 12393
rect 9312 12384 9364 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 11244 12384 11296 12436
rect 17040 12384 17092 12436
rect 17776 12427 17828 12436
rect 17776 12393 17785 12427
rect 17785 12393 17819 12427
rect 17819 12393 17828 12427
rect 17776 12384 17828 12393
rect 4068 12316 4120 12368
rect 2228 12291 2280 12300
rect 2228 12257 2237 12291
rect 2237 12257 2271 12291
rect 2271 12257 2280 12291
rect 2228 12248 2280 12257
rect 2136 12180 2188 12232
rect 2688 12180 2740 12232
rect 3148 12180 3200 12232
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 5816 12180 5868 12232
rect 7840 12180 7892 12232
rect 8576 12248 8628 12300
rect 9128 12248 9180 12300
rect 11060 12291 11112 12300
rect 11060 12257 11069 12291
rect 11069 12257 11103 12291
rect 11103 12257 11112 12291
rect 11060 12248 11112 12257
rect 11980 12248 12032 12300
rect 12164 12291 12216 12300
rect 12164 12257 12173 12291
rect 12173 12257 12207 12291
rect 12207 12257 12216 12291
rect 12164 12248 12216 12257
rect 13912 12291 13964 12300
rect 13912 12257 13921 12291
rect 13921 12257 13955 12291
rect 13955 12257 13964 12291
rect 13912 12248 13964 12257
rect 15568 12291 15620 12300
rect 15568 12257 15577 12291
rect 15577 12257 15611 12291
rect 15611 12257 15620 12291
rect 15568 12248 15620 12257
rect 16672 12291 16724 12300
rect 16672 12257 16681 12291
rect 16681 12257 16715 12291
rect 16715 12257 16724 12291
rect 16672 12248 16724 12257
rect 17316 12248 17368 12300
rect 17500 12248 17552 12300
rect 5632 12112 5684 12164
rect 6920 12112 6972 12164
rect 7380 12112 7432 12164
rect 8944 12180 8996 12232
rect 9404 12180 9456 12232
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 10876 12180 10928 12232
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 4620 12044 4672 12096
rect 14188 12112 14240 12164
rect 10416 12044 10468 12096
rect 10876 12044 10928 12096
rect 11888 12044 11940 12096
rect 15384 12180 15436 12232
rect 17040 12180 17092 12232
rect 17868 12223 17920 12232
rect 17868 12189 17877 12223
rect 17877 12189 17911 12223
rect 17911 12189 17920 12223
rect 17868 12180 17920 12189
rect 15568 12112 15620 12164
rect 17684 12112 17736 12164
rect 16304 12087 16356 12096
rect 16304 12053 16313 12087
rect 16313 12053 16347 12087
rect 16347 12053 16356 12087
rect 16304 12044 16356 12053
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 2136 11883 2188 11892
rect 2136 11849 2145 11883
rect 2145 11849 2179 11883
rect 2179 11849 2188 11883
rect 2136 11840 2188 11849
rect 3148 11883 3200 11892
rect 3148 11849 3157 11883
rect 3157 11849 3191 11883
rect 3191 11849 3200 11883
rect 3148 11840 3200 11849
rect 4620 11883 4672 11892
rect 4620 11849 4629 11883
rect 4629 11849 4663 11883
rect 4663 11849 4672 11883
rect 4620 11840 4672 11849
rect 8852 11883 8904 11892
rect 3240 11772 3292 11824
rect 3608 11772 3660 11824
rect 6000 11772 6052 11824
rect 2412 11568 2464 11620
rect 5264 11747 5316 11756
rect 5264 11713 5273 11747
rect 5273 11713 5307 11747
rect 5307 11713 5316 11747
rect 5264 11704 5316 11713
rect 7656 11772 7708 11824
rect 8852 11849 8861 11883
rect 8861 11849 8895 11883
rect 8895 11849 8904 11883
rect 8852 11840 8904 11849
rect 8944 11840 8996 11892
rect 10692 11883 10744 11892
rect 9680 11772 9732 11824
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 6920 11704 6972 11756
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 8024 11704 8076 11756
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 6276 11636 6328 11688
rect 7380 11636 7432 11688
rect 8208 11636 8260 11688
rect 8576 11704 8628 11756
rect 10692 11849 10701 11883
rect 10701 11849 10735 11883
rect 10735 11849 10744 11883
rect 10692 11840 10744 11849
rect 13912 11840 13964 11892
rect 15200 11840 15252 11892
rect 19432 11840 19484 11892
rect 12072 11772 12124 11824
rect 14464 11772 14516 11824
rect 8668 11636 8720 11688
rect 10968 11636 11020 11688
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 13176 11704 13228 11756
rect 15568 11772 15620 11824
rect 14740 11704 14792 11756
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 15016 11636 15068 11688
rect 16856 11636 16908 11688
rect 2688 11568 2740 11620
rect 5356 11568 5408 11620
rect 2596 11543 2648 11552
rect 2596 11509 2605 11543
rect 2605 11509 2639 11543
rect 2639 11509 2648 11543
rect 2596 11500 2648 11509
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 4068 11500 4120 11552
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 6644 11568 6696 11620
rect 7288 11611 7340 11620
rect 7288 11577 7297 11611
rect 7297 11577 7331 11611
rect 7331 11577 7340 11611
rect 7288 11568 7340 11577
rect 8024 11500 8076 11552
rect 8576 11568 8628 11620
rect 11428 11568 11480 11620
rect 12624 11568 12676 11620
rect 13636 11568 13688 11620
rect 15292 11568 15344 11620
rect 16580 11568 16632 11620
rect 16764 11568 16816 11620
rect 8944 11500 8996 11552
rect 9220 11543 9272 11552
rect 9220 11509 9229 11543
rect 9229 11509 9263 11543
rect 9263 11509 9272 11543
rect 9220 11500 9272 11509
rect 9588 11500 9640 11552
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 17040 11500 17092 11552
rect 17776 11500 17828 11552
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 2320 11296 2372 11348
rect 2688 11296 2740 11348
rect 5724 11296 5776 11348
rect 1400 11160 1452 11212
rect 2412 11203 2464 11212
rect 2412 11169 2446 11203
rect 2446 11169 2464 11203
rect 2412 11160 2464 11169
rect 6368 11228 6420 11280
rect 9220 11296 9272 11348
rect 10600 11296 10652 11348
rect 10324 11228 10376 11280
rect 4712 11160 4764 11212
rect 5816 11160 5868 11212
rect 7380 11160 7432 11212
rect 8024 11160 8076 11212
rect 10692 11160 10744 11212
rect 11704 11296 11756 11348
rect 17132 11296 17184 11348
rect 14004 11228 14056 11280
rect 14188 11228 14240 11280
rect 11336 11160 11388 11212
rect 13544 11203 13596 11212
rect 13544 11169 13578 11203
rect 13578 11169 13596 11203
rect 13544 11160 13596 11169
rect 15568 11203 15620 11212
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 6920 11092 6972 11144
rect 9220 11092 9272 11144
rect 9496 11092 9548 11144
rect 5448 11067 5500 11076
rect 5448 11033 5457 11067
rect 5457 11033 5491 11067
rect 5491 11033 5500 11067
rect 5448 11024 5500 11033
rect 7564 11024 7616 11076
rect 9404 11024 9456 11076
rect 3792 10956 3844 11008
rect 8576 10956 8628 11008
rect 13176 11092 13228 11144
rect 10968 11024 11020 11076
rect 11796 11024 11848 11076
rect 10692 10956 10744 11008
rect 11612 10956 11664 11008
rect 15568 11169 15602 11203
rect 15602 11169 15620 11203
rect 15568 11160 15620 11169
rect 17684 11135 17736 11144
rect 14740 10956 14792 11008
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 16580 11024 16632 11076
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 2228 10752 2280 10804
rect 3608 10752 3660 10804
rect 4252 10752 4304 10804
rect 5264 10752 5316 10804
rect 5356 10752 5408 10804
rect 9588 10752 9640 10804
rect 10324 10752 10376 10804
rect 11152 10795 11204 10804
rect 11152 10761 11161 10795
rect 11161 10761 11195 10795
rect 11195 10761 11204 10795
rect 11152 10752 11204 10761
rect 3792 10684 3844 10736
rect 2412 10616 2464 10668
rect 6276 10684 6328 10736
rect 6920 10684 6972 10736
rect 4712 10616 4764 10668
rect 5448 10616 5500 10668
rect 6368 10616 6420 10668
rect 1676 10548 1728 10600
rect 2872 10480 2924 10532
rect 5540 10548 5592 10600
rect 5908 10591 5960 10600
rect 5908 10557 5917 10591
rect 5917 10557 5951 10591
rect 5951 10557 5960 10591
rect 5908 10548 5960 10557
rect 3884 10455 3936 10464
rect 3884 10421 3893 10455
rect 3893 10421 3927 10455
rect 3927 10421 3936 10455
rect 3884 10412 3936 10421
rect 5356 10480 5408 10532
rect 5724 10480 5776 10532
rect 6552 10480 6604 10532
rect 7104 10616 7156 10668
rect 7564 10616 7616 10668
rect 9496 10684 9548 10736
rect 11244 10684 11296 10736
rect 7288 10548 7340 10600
rect 9680 10616 9732 10668
rect 9864 10616 9916 10668
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 10324 10548 10376 10600
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 11428 10616 11480 10668
rect 11244 10548 11296 10600
rect 13360 10752 13412 10804
rect 13728 10752 13780 10804
rect 16672 10752 16724 10804
rect 12164 10548 12216 10600
rect 13176 10548 13228 10600
rect 13452 10548 13504 10600
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 14740 10591 14792 10600
rect 14740 10557 14749 10591
rect 14749 10557 14783 10591
rect 14783 10557 14792 10591
rect 14740 10548 14792 10557
rect 16856 10616 16908 10668
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 17868 10616 17920 10668
rect 7748 10412 7800 10464
rect 8024 10412 8076 10464
rect 11796 10480 11848 10532
rect 15844 10548 15896 10600
rect 16488 10548 16540 10600
rect 17500 10548 17552 10600
rect 17040 10480 17092 10532
rect 8852 10412 8904 10464
rect 9496 10412 9548 10464
rect 9680 10412 9732 10464
rect 10508 10412 10560 10464
rect 11428 10412 11480 10464
rect 12716 10412 12768 10464
rect 13544 10412 13596 10464
rect 15200 10412 15252 10464
rect 15476 10412 15528 10464
rect 15844 10412 15896 10464
rect 16028 10412 16080 10464
rect 16580 10455 16632 10464
rect 16580 10421 16589 10455
rect 16589 10421 16623 10455
rect 16623 10421 16632 10455
rect 16580 10412 16632 10421
rect 16672 10412 16724 10464
rect 18420 10412 18472 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 2964 10208 3016 10260
rect 3424 10208 3476 10260
rect 3884 10208 3936 10260
rect 5540 10208 5592 10260
rect 6000 10208 6052 10260
rect 6184 10208 6236 10260
rect 6736 10208 6788 10260
rect 9680 10208 9732 10260
rect 2320 10140 2372 10192
rect 4068 10140 4120 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 1952 10072 2004 10124
rect 3056 10115 3108 10124
rect 3056 10081 3065 10115
rect 3065 10081 3099 10115
rect 3099 10081 3108 10115
rect 3056 10072 3108 10081
rect 5080 10072 5132 10124
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 5540 10072 5592 10124
rect 5816 10072 5868 10124
rect 6276 10072 6328 10124
rect 6920 10140 6972 10192
rect 7472 10140 7524 10192
rect 8484 10183 8536 10192
rect 8484 10149 8493 10183
rect 8493 10149 8527 10183
rect 8527 10149 8536 10183
rect 8484 10140 8536 10149
rect 8576 10140 8628 10192
rect 10324 10208 10376 10260
rect 11428 10208 11480 10260
rect 12716 10208 12768 10260
rect 13452 10208 13504 10260
rect 13820 10208 13872 10260
rect 14280 10251 14332 10260
rect 14280 10217 14289 10251
rect 14289 10217 14323 10251
rect 14323 10217 14332 10251
rect 14280 10208 14332 10217
rect 14372 10208 14424 10260
rect 15108 10208 15160 10260
rect 15292 10251 15344 10260
rect 15292 10217 15301 10251
rect 15301 10217 15335 10251
rect 15335 10217 15344 10251
rect 15292 10208 15344 10217
rect 4712 9936 4764 9988
rect 6184 10004 6236 10056
rect 3148 9868 3200 9920
rect 4528 9868 4580 9920
rect 6368 9936 6420 9988
rect 7472 9936 7524 9988
rect 9680 10072 9732 10124
rect 9864 10072 9916 10124
rect 11244 10140 11296 10192
rect 11612 10183 11664 10192
rect 11612 10149 11621 10183
rect 11621 10149 11655 10183
rect 11655 10149 11664 10183
rect 11612 10140 11664 10149
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 9128 9936 9180 9988
rect 8208 9868 8260 9920
rect 9496 9936 9548 9988
rect 9864 9936 9916 9988
rect 9956 9936 10008 9988
rect 10692 9936 10744 9988
rect 11060 9936 11112 9988
rect 13268 10072 13320 10124
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 14280 10004 14332 10056
rect 14556 10072 14608 10124
rect 15292 10072 15344 10124
rect 15568 10140 15620 10192
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 15752 10115 15804 10124
rect 15752 10081 15761 10115
rect 15761 10081 15795 10115
rect 15795 10081 15804 10115
rect 15752 10072 15804 10081
rect 15568 10004 15620 10056
rect 16948 10140 17000 10192
rect 17408 10072 17460 10124
rect 17868 10047 17920 10056
rect 11428 9868 11480 9920
rect 14004 9868 14056 9920
rect 14188 9868 14240 9920
rect 14740 9868 14792 9920
rect 15108 9868 15160 9920
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 16028 9936 16080 9988
rect 17316 9979 17368 9988
rect 17316 9945 17325 9979
rect 17325 9945 17359 9979
rect 17359 9945 17368 9979
rect 17316 9936 17368 9945
rect 16488 9868 16540 9920
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 4712 9664 4764 9716
rect 6920 9664 6972 9716
rect 8852 9707 8904 9716
rect 8852 9673 8861 9707
rect 8861 9673 8895 9707
rect 8895 9673 8904 9707
rect 8852 9664 8904 9673
rect 9128 9664 9180 9716
rect 10692 9664 10744 9716
rect 11612 9664 11664 9716
rect 13728 9664 13780 9716
rect 11060 9639 11112 9648
rect 6276 9528 6328 9580
rect 11060 9605 11069 9639
rect 11069 9605 11103 9639
rect 11103 9605 11112 9639
rect 11060 9596 11112 9605
rect 11336 9639 11388 9648
rect 11336 9605 11345 9639
rect 11345 9605 11379 9639
rect 11379 9605 11388 9639
rect 11336 9596 11388 9605
rect 15016 9664 15068 9716
rect 16488 9664 16540 9716
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 2964 9460 3016 9512
rect 3056 9460 3108 9512
rect 3516 9392 3568 9444
rect 4528 9460 4580 9512
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 7380 9460 7432 9512
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 3792 9324 3844 9376
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 4436 9367 4488 9376
rect 4436 9333 4445 9367
rect 4445 9333 4479 9367
rect 4479 9333 4488 9367
rect 4436 9324 4488 9333
rect 5448 9392 5500 9444
rect 8576 9460 8628 9512
rect 11244 9503 11296 9512
rect 7748 9435 7800 9444
rect 7748 9401 7782 9435
rect 7782 9401 7800 9435
rect 7748 9392 7800 9401
rect 5540 9324 5592 9376
rect 11244 9469 11253 9503
rect 11253 9469 11287 9503
rect 11287 9469 11296 9503
rect 11244 9460 11296 9469
rect 11612 9460 11664 9512
rect 13268 9528 13320 9580
rect 13728 9528 13780 9580
rect 14096 9596 14148 9648
rect 14188 9528 14240 9580
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 15108 9528 15160 9580
rect 12072 9460 12124 9512
rect 12164 9460 12216 9512
rect 12900 9460 12952 9512
rect 14832 9460 14884 9512
rect 15844 9503 15896 9512
rect 15844 9469 15878 9503
rect 15878 9469 15896 9503
rect 15844 9460 15896 9469
rect 16764 9460 16816 9512
rect 17316 9460 17368 9512
rect 9312 9392 9364 9444
rect 10600 9392 10652 9444
rect 10692 9392 10744 9444
rect 12716 9392 12768 9444
rect 9588 9324 9640 9376
rect 10324 9324 10376 9376
rect 10784 9324 10836 9376
rect 11796 9367 11848 9376
rect 11796 9333 11805 9367
rect 11805 9333 11839 9367
rect 11839 9333 11848 9367
rect 17500 9435 17552 9444
rect 17500 9401 17509 9435
rect 17509 9401 17543 9435
rect 17543 9401 17552 9435
rect 17500 9392 17552 9401
rect 11796 9324 11848 9333
rect 13176 9324 13228 9376
rect 13544 9324 13596 9376
rect 14372 9367 14424 9376
rect 14372 9333 14381 9367
rect 14381 9333 14415 9367
rect 14415 9333 14424 9367
rect 14372 9324 14424 9333
rect 16396 9324 16448 9376
rect 17224 9324 17276 9376
rect 17868 9324 17920 9376
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 2136 9120 2188 9172
rect 4620 9120 4672 9172
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 7288 9120 7340 9172
rect 7932 9163 7984 9172
rect 7932 9129 7941 9163
rect 7941 9129 7975 9163
rect 7975 9129 7984 9163
rect 7932 9120 7984 9129
rect 8024 9120 8076 9172
rect 3332 9052 3384 9104
rect 4436 9052 4488 9104
rect 1952 8984 2004 9036
rect 2688 8984 2740 9036
rect 2964 8984 3016 9036
rect 3700 8984 3752 9036
rect 4344 9027 4396 9036
rect 4344 8993 4378 9027
rect 4378 8993 4396 9027
rect 6276 9027 6328 9036
rect 4344 8984 4396 8993
rect 2412 8916 2464 8968
rect 3792 8916 3844 8968
rect 1124 8780 1176 8832
rect 5080 8780 5132 8832
rect 6276 8993 6285 9027
rect 6285 8993 6319 9027
rect 6319 8993 6328 9027
rect 6276 8984 6328 8993
rect 7564 8984 7616 9036
rect 8300 9027 8352 9036
rect 8300 8993 8309 9027
rect 8309 8993 8343 9027
rect 8343 8993 8352 9027
rect 8300 8984 8352 8993
rect 8944 9120 8996 9172
rect 9128 9120 9180 9172
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 10876 9120 10928 9172
rect 11796 9120 11848 9172
rect 14372 9120 14424 9172
rect 14556 9120 14608 9172
rect 14924 9120 14976 9172
rect 16304 9120 16356 9172
rect 16672 9120 16724 9172
rect 8576 9052 8628 9104
rect 9588 9052 9640 9104
rect 12348 9052 12400 9104
rect 12532 8984 12584 9036
rect 12624 8984 12676 9036
rect 8668 8916 8720 8968
rect 8852 8916 8904 8968
rect 8944 8916 8996 8968
rect 10048 8916 10100 8968
rect 8116 8780 8168 8832
rect 10140 8848 10192 8900
rect 11060 8916 11112 8968
rect 11980 8916 12032 8968
rect 12164 8916 12216 8968
rect 12440 8916 12492 8968
rect 13268 9052 13320 9104
rect 13728 9027 13780 9036
rect 13728 8993 13762 9027
rect 13762 8993 13780 9027
rect 13728 8984 13780 8993
rect 15108 8984 15160 9036
rect 17224 8984 17276 9036
rect 18052 9027 18104 9036
rect 18052 8993 18061 9027
rect 18061 8993 18095 9027
rect 18095 8993 18104 9027
rect 18052 8984 18104 8993
rect 10692 8780 10744 8832
rect 12348 8780 12400 8832
rect 15844 8916 15896 8968
rect 15108 8848 15160 8900
rect 15016 8780 15068 8832
rect 16764 8780 16816 8832
rect 18328 8780 18380 8832
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 3240 8576 3292 8628
rect 8300 8576 8352 8628
rect 9036 8576 9088 8628
rect 4344 8508 4396 8560
rect 6736 8508 6788 8560
rect 8576 8508 8628 8560
rect 11060 8576 11112 8628
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 3332 8440 3384 8492
rect 4620 8440 4672 8492
rect 6276 8440 6328 8492
rect 6644 8440 6696 8492
rect 8944 8440 8996 8492
rect 9312 8440 9364 8492
rect 6000 8415 6052 8424
rect 6000 8381 6009 8415
rect 6009 8381 6043 8415
rect 6043 8381 6052 8415
rect 6000 8372 6052 8381
rect 2596 8347 2648 8356
rect 2596 8313 2630 8347
rect 2630 8313 2648 8347
rect 2596 8304 2648 8313
rect 3240 8304 3292 8356
rect 4252 8304 4304 8356
rect 6460 8304 6512 8356
rect 8668 8372 8720 8424
rect 9036 8372 9088 8424
rect 10048 8415 10100 8424
rect 8116 8304 8168 8356
rect 8576 8304 8628 8356
rect 2412 8236 2464 8288
rect 2964 8236 3016 8288
rect 3056 8236 3108 8288
rect 3608 8236 3660 8288
rect 4344 8279 4396 8288
rect 4344 8245 4353 8279
rect 4353 8245 4387 8279
rect 4387 8245 4396 8279
rect 4344 8236 4396 8245
rect 4528 8236 4580 8288
rect 5264 8236 5316 8288
rect 5356 8279 5408 8288
rect 5356 8245 5365 8279
rect 5365 8245 5399 8279
rect 5399 8245 5408 8279
rect 6184 8279 6236 8288
rect 5356 8236 5408 8245
rect 6184 8245 6193 8279
rect 6193 8245 6227 8279
rect 6227 8245 6236 8279
rect 6184 8236 6236 8245
rect 6552 8236 6604 8288
rect 8944 8279 8996 8288
rect 8944 8245 8953 8279
rect 8953 8245 8987 8279
rect 8987 8245 8996 8279
rect 8944 8236 8996 8245
rect 10048 8381 10057 8415
rect 10057 8381 10091 8415
rect 10091 8381 10100 8415
rect 10048 8372 10100 8381
rect 10876 8372 10928 8424
rect 12164 8576 12216 8628
rect 12348 8576 12400 8628
rect 11336 8508 11388 8560
rect 9864 8304 9916 8356
rect 10692 8304 10744 8356
rect 10968 8304 11020 8356
rect 13912 8508 13964 8560
rect 14188 8508 14240 8560
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 12164 8440 12216 8492
rect 12716 8372 12768 8424
rect 12900 8440 12952 8492
rect 13268 8440 13320 8492
rect 13452 8440 13504 8492
rect 17224 8483 17276 8492
rect 14372 8372 14424 8424
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 14924 8304 14976 8356
rect 15660 8372 15712 8424
rect 16488 8372 16540 8424
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 18236 8551 18288 8560
rect 18236 8517 18245 8551
rect 18245 8517 18279 8551
rect 18279 8517 18288 8551
rect 18236 8508 18288 8517
rect 17132 8372 17184 8381
rect 15108 8304 15160 8356
rect 16764 8304 16816 8356
rect 17224 8304 17276 8356
rect 17684 8304 17736 8356
rect 11152 8236 11204 8288
rect 11888 8236 11940 8288
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 12440 8236 12492 8245
rect 12624 8236 12676 8288
rect 16212 8236 16264 8288
rect 16304 8236 16356 8288
rect 16672 8279 16724 8288
rect 16672 8245 16681 8279
rect 16681 8245 16715 8279
rect 16715 8245 16724 8279
rect 16672 8236 16724 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 3516 8032 3568 8084
rect 4436 8032 4488 8084
rect 7656 8032 7708 8084
rect 8392 8075 8444 8084
rect 8392 8041 8401 8075
rect 8401 8041 8435 8075
rect 8435 8041 8444 8075
rect 8392 8032 8444 8041
rect 8484 8032 8536 8084
rect 9864 8032 9916 8084
rect 12164 8032 12216 8084
rect 12348 8032 12400 8084
rect 12624 8032 12676 8084
rect 13728 8032 13780 8084
rect 16212 8032 16264 8084
rect 17960 8032 18012 8084
rect 6552 7964 6604 8016
rect 6736 7964 6788 8016
rect 5080 7939 5132 7948
rect 2504 7828 2556 7880
rect 3056 7828 3108 7880
rect 1952 7735 2004 7744
rect 1952 7701 1961 7735
rect 1961 7701 1995 7735
rect 1995 7701 2004 7735
rect 1952 7692 2004 7701
rect 2320 7760 2372 7812
rect 3424 7760 3476 7812
rect 3792 7828 3844 7880
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 3516 7692 3568 7744
rect 5080 7905 5089 7939
rect 5089 7905 5123 7939
rect 5123 7905 5132 7939
rect 5080 7896 5132 7905
rect 7380 7896 7432 7948
rect 8024 7896 8076 7948
rect 11888 7964 11940 8016
rect 12256 7964 12308 8016
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 6644 7828 6696 7880
rect 8852 7828 8904 7880
rect 9404 7828 9456 7880
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 12072 7896 12124 7948
rect 13268 7939 13320 7948
rect 13268 7905 13291 7939
rect 13291 7905 13320 7939
rect 13268 7896 13320 7905
rect 14372 7896 14424 7948
rect 16304 7896 16356 7948
rect 17316 7939 17368 7948
rect 8392 7760 8444 7812
rect 10048 7760 10100 7812
rect 10600 7760 10652 7812
rect 15108 7828 15160 7880
rect 7748 7692 7800 7744
rect 13360 7692 13412 7744
rect 14556 7692 14608 7744
rect 15200 7692 15252 7744
rect 15568 7692 15620 7744
rect 17316 7905 17325 7939
rect 17325 7905 17359 7939
rect 17359 7905 17368 7939
rect 17316 7896 17368 7905
rect 16764 7760 16816 7812
rect 17684 7760 17736 7812
rect 16580 7692 16632 7744
rect 16948 7735 17000 7744
rect 16948 7701 16957 7735
rect 16957 7701 16991 7735
rect 16991 7701 17000 7735
rect 16948 7692 17000 7701
rect 17776 7692 17828 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 2504 7488 2556 7540
rect 3700 7488 3752 7540
rect 4528 7488 4580 7540
rect 4712 7488 4764 7540
rect 10324 7488 10376 7540
rect 4344 7420 4396 7472
rect 7840 7420 7892 7472
rect 10600 7420 10652 7472
rect 10968 7420 11020 7472
rect 11244 7488 11296 7540
rect 11980 7488 12032 7540
rect 12716 7488 12768 7540
rect 13452 7488 13504 7540
rect 2320 7352 2372 7404
rect 3056 7352 3108 7404
rect 3424 7395 3476 7404
rect 3424 7361 3433 7395
rect 3433 7361 3467 7395
rect 3467 7361 3476 7395
rect 3424 7352 3476 7361
rect 4528 7327 4580 7336
rect 2872 7216 2924 7268
rect 4528 7293 4537 7327
rect 4537 7293 4571 7327
rect 4571 7293 4580 7327
rect 4528 7284 4580 7293
rect 6276 7352 6328 7404
rect 8024 7352 8076 7404
rect 7840 7327 7892 7336
rect 7840 7293 7849 7327
rect 7849 7293 7883 7327
rect 7883 7293 7892 7327
rect 7840 7284 7892 7293
rect 11152 7352 11204 7404
rect 12256 7420 12308 7472
rect 16396 7420 16448 7472
rect 9128 7284 9180 7336
rect 11244 7284 11296 7336
rect 12532 7352 12584 7404
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 13820 7352 13872 7404
rect 16764 7352 16816 7404
rect 15108 7284 15160 7336
rect 15200 7284 15252 7336
rect 16120 7284 16172 7336
rect 16212 7284 16264 7336
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 2320 7191 2372 7200
rect 2320 7157 2329 7191
rect 2329 7157 2363 7191
rect 2363 7157 2372 7191
rect 2320 7148 2372 7157
rect 2964 7148 3016 7200
rect 6736 7216 6788 7268
rect 7564 7216 7616 7268
rect 7656 7216 7708 7268
rect 9036 7216 9088 7268
rect 11060 7216 11112 7268
rect 12716 7216 12768 7268
rect 14464 7216 14516 7268
rect 14556 7216 14608 7268
rect 16672 7284 16724 7336
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 5632 7148 5684 7200
rect 6552 7148 6604 7200
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 10968 7148 11020 7200
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 14004 7148 14056 7200
rect 15568 7191 15620 7200
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 16120 7148 16172 7200
rect 16488 7148 16540 7200
rect 17868 7148 17920 7200
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 1952 6944 2004 6996
rect 4436 6944 4488 6996
rect 6276 6987 6328 6996
rect 6276 6953 6285 6987
rect 6285 6953 6319 6987
rect 6319 6953 6328 6987
rect 6276 6944 6328 6953
rect 6460 6944 6512 6996
rect 7564 6987 7616 6996
rect 3424 6876 3476 6928
rect 2964 6808 3016 6860
rect 3332 6808 3384 6860
rect 4068 6851 4120 6860
rect 3056 6672 3108 6724
rect 3700 6672 3752 6724
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 5540 6876 5592 6928
rect 4528 6740 4580 6792
rect 6644 6740 6696 6792
rect 7564 6953 7573 6987
rect 7573 6953 7607 6987
rect 7607 6953 7616 6987
rect 7564 6944 7616 6953
rect 8116 6944 8168 6996
rect 7932 6919 7984 6928
rect 7932 6885 7941 6919
rect 7941 6885 7975 6919
rect 7975 6885 7984 6919
rect 7932 6876 7984 6885
rect 8392 6944 8444 6996
rect 9036 6944 9088 6996
rect 10692 6944 10744 6996
rect 11244 6944 11296 6996
rect 9220 6876 9272 6928
rect 9588 6876 9640 6928
rect 8024 6783 8076 6792
rect 2504 6604 2556 6656
rect 3608 6647 3660 6656
rect 3608 6613 3617 6647
rect 3617 6613 3651 6647
rect 3651 6613 3660 6647
rect 3608 6604 3660 6613
rect 3792 6604 3844 6656
rect 7380 6672 7432 6724
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 8208 6672 8260 6724
rect 8576 6715 8628 6724
rect 8576 6681 8585 6715
rect 8585 6681 8619 6715
rect 8619 6681 8628 6715
rect 8576 6672 8628 6681
rect 8852 6740 8904 6792
rect 10416 6808 10468 6860
rect 13452 6944 13504 6996
rect 13820 6944 13872 6996
rect 14188 6944 14240 6996
rect 14372 6987 14424 6996
rect 14372 6953 14381 6987
rect 14381 6953 14415 6987
rect 14415 6953 14424 6987
rect 14372 6944 14424 6953
rect 13728 6876 13780 6928
rect 18052 6876 18104 6928
rect 9220 6740 9272 6792
rect 10324 6740 10376 6792
rect 12072 6808 12124 6860
rect 11060 6783 11112 6792
rect 10416 6672 10468 6724
rect 11060 6749 11069 6783
rect 11069 6749 11103 6783
rect 11103 6749 11112 6783
rect 11060 6740 11112 6749
rect 11152 6740 11204 6792
rect 13268 6808 13320 6860
rect 16580 6808 16632 6860
rect 17132 6808 17184 6860
rect 13084 6740 13136 6792
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 15108 6740 15160 6792
rect 17224 6740 17276 6792
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 18144 6783 18196 6792
rect 17684 6740 17736 6749
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 6000 6604 6052 6656
rect 7196 6604 7248 6656
rect 7564 6604 7616 6656
rect 11244 6604 11296 6656
rect 12992 6672 13044 6724
rect 14372 6672 14424 6724
rect 16764 6672 16816 6724
rect 16856 6647 16908 6656
rect 16856 6613 16865 6647
rect 16865 6613 16899 6647
rect 16899 6613 16908 6647
rect 16856 6604 16908 6613
rect 17224 6604 17276 6656
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 2228 6400 2280 6452
rect 3424 6400 3476 6452
rect 6184 6400 6236 6452
rect 6276 6400 6328 6452
rect 7472 6400 7524 6452
rect 8208 6443 8260 6452
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 8300 6400 8352 6452
rect 10416 6400 10468 6452
rect 14004 6443 14056 6452
rect 2504 6332 2556 6384
rect 2228 6264 2280 6316
rect 2596 6196 2648 6248
rect 5540 6264 5592 6316
rect 5816 6264 5868 6316
rect 8208 6264 8260 6316
rect 10140 6332 10192 6384
rect 12716 6332 12768 6384
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 14372 6400 14424 6452
rect 15384 6400 15436 6452
rect 3056 6239 3108 6248
rect 3056 6205 3090 6239
rect 3090 6205 3108 6239
rect 3056 6196 3108 6205
rect 3608 6196 3660 6248
rect 4528 6196 4580 6248
rect 6460 6196 6512 6248
rect 2964 6128 3016 6180
rect 2872 6060 2924 6112
rect 3056 6060 3108 6112
rect 4620 6128 4672 6180
rect 4528 6060 4580 6112
rect 5908 6060 5960 6112
rect 6736 6060 6788 6112
rect 8576 6196 8628 6248
rect 7472 6128 7524 6180
rect 12164 6264 12216 6316
rect 13728 6264 13780 6316
rect 14464 6264 14516 6316
rect 11336 6128 11388 6180
rect 11980 6128 12032 6180
rect 15108 6196 15160 6248
rect 13636 6128 13688 6180
rect 13820 6128 13872 6180
rect 15476 6171 15528 6180
rect 15476 6137 15485 6171
rect 15485 6137 15519 6171
rect 15519 6137 15528 6171
rect 15476 6128 15528 6137
rect 16856 6128 16908 6180
rect 17316 6128 17368 6180
rect 8484 6060 8536 6112
rect 11244 6060 11296 6112
rect 11612 6060 11664 6112
rect 12072 6103 12124 6112
rect 12072 6069 12081 6103
rect 12081 6069 12115 6103
rect 12115 6069 12124 6103
rect 12072 6060 12124 6069
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 13452 6060 13504 6069
rect 13912 6060 13964 6112
rect 14096 6060 14148 6112
rect 14556 6060 14608 6112
rect 14740 6060 14792 6112
rect 14924 6060 14976 6112
rect 15200 6060 15252 6112
rect 15384 6103 15436 6112
rect 15384 6069 15393 6103
rect 15393 6069 15427 6103
rect 15427 6069 15436 6103
rect 15384 6060 15436 6069
rect 15660 6060 15712 6112
rect 17776 6060 17828 6112
rect 18236 6103 18288 6112
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 2320 5856 2372 5908
rect 2872 5899 2924 5908
rect 2872 5865 2881 5899
rect 2881 5865 2915 5899
rect 2915 5865 2924 5899
rect 2872 5856 2924 5865
rect 3976 5856 4028 5908
rect 4436 5899 4488 5908
rect 4436 5865 4445 5899
rect 4445 5865 4479 5899
rect 4479 5865 4488 5899
rect 4436 5856 4488 5865
rect 4988 5856 5040 5908
rect 6644 5856 6696 5908
rect 8024 5856 8076 5908
rect 1768 5788 1820 5840
rect 4252 5788 4304 5840
rect 10784 5856 10836 5908
rect 11244 5856 11296 5908
rect 12624 5856 12676 5908
rect 13176 5856 13228 5908
rect 14464 5856 14516 5908
rect 16120 5856 16172 5908
rect 18144 5856 18196 5908
rect 8944 5788 8996 5840
rect 9036 5788 9088 5840
rect 10416 5788 10468 5840
rect 3148 5720 3200 5772
rect 2320 5695 2372 5704
rect 2320 5661 2329 5695
rect 2329 5661 2363 5695
rect 2363 5661 2372 5695
rect 2320 5652 2372 5661
rect 3056 5652 3108 5704
rect 2688 5584 2740 5636
rect 2872 5584 2924 5636
rect 2504 5516 2556 5568
rect 3332 5516 3384 5568
rect 3608 5584 3660 5636
rect 3976 5584 4028 5636
rect 4344 5720 4396 5772
rect 4896 5720 4948 5772
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 4804 5652 4856 5704
rect 5356 5652 5408 5704
rect 5908 5720 5960 5772
rect 6184 5720 6236 5772
rect 6368 5720 6420 5772
rect 9128 5763 9180 5772
rect 5816 5652 5868 5704
rect 4712 5584 4764 5636
rect 7472 5695 7524 5704
rect 7472 5661 7481 5695
rect 7481 5661 7515 5695
rect 7515 5661 7524 5695
rect 7472 5652 7524 5661
rect 8484 5652 8536 5704
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 10324 5720 10376 5772
rect 12532 5788 12584 5840
rect 11152 5763 11204 5772
rect 9312 5652 9364 5661
rect 10416 5652 10468 5704
rect 11152 5729 11161 5763
rect 11161 5729 11195 5763
rect 11195 5729 11204 5763
rect 11152 5720 11204 5729
rect 12164 5720 12216 5772
rect 15108 5788 15160 5840
rect 16948 5788 17000 5840
rect 17408 5788 17460 5840
rect 15016 5720 15068 5772
rect 15476 5720 15528 5772
rect 8944 5584 8996 5636
rect 4804 5516 4856 5568
rect 5080 5559 5132 5568
rect 5080 5525 5089 5559
rect 5089 5525 5123 5559
rect 5123 5525 5132 5559
rect 5080 5516 5132 5525
rect 6000 5516 6052 5568
rect 7196 5516 7248 5568
rect 7564 5516 7616 5568
rect 8024 5516 8076 5568
rect 8208 5516 8260 5568
rect 11060 5652 11112 5704
rect 13912 5652 13964 5704
rect 14740 5652 14792 5704
rect 12532 5627 12584 5636
rect 12532 5593 12541 5627
rect 12541 5593 12575 5627
rect 12575 5593 12584 5627
rect 12532 5584 12584 5593
rect 14188 5584 14240 5636
rect 14924 5584 14976 5636
rect 11060 5516 11112 5568
rect 15384 5559 15436 5568
rect 15384 5525 15393 5559
rect 15393 5525 15427 5559
rect 15427 5525 15436 5559
rect 15384 5516 15436 5525
rect 16304 5652 16356 5704
rect 17316 5652 17368 5704
rect 17684 5652 17736 5704
rect 16580 5559 16632 5568
rect 16580 5525 16589 5559
rect 16589 5525 16623 5559
rect 16623 5525 16632 5559
rect 16580 5516 16632 5525
rect 16948 5559 17000 5568
rect 16948 5525 16957 5559
rect 16957 5525 16991 5559
rect 16991 5525 17000 5559
rect 16948 5516 17000 5525
rect 17868 5516 17920 5568
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 3056 5312 3108 5364
rect 4988 5312 5040 5364
rect 5356 5312 5408 5364
rect 7380 5312 7432 5364
rect 7932 5312 7984 5364
rect 11796 5312 11848 5364
rect 13452 5312 13504 5364
rect 14188 5312 14240 5364
rect 14556 5312 14608 5364
rect 17960 5312 18012 5364
rect 3884 5244 3936 5296
rect 4436 5176 4488 5228
rect 4620 5219 4672 5228
rect 4620 5185 4629 5219
rect 4629 5185 4663 5219
rect 4663 5185 4672 5219
rect 4620 5176 4672 5185
rect 1400 5040 1452 5092
rect 2228 5040 2280 5092
rect 5908 5176 5960 5228
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 8392 5219 8444 5228
rect 7472 5176 7524 5185
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 9036 5244 9088 5296
rect 10416 5287 10468 5296
rect 10416 5253 10425 5287
rect 10425 5253 10459 5287
rect 10459 5253 10468 5287
rect 10416 5244 10468 5253
rect 8576 5108 8628 5160
rect 9036 5151 9088 5160
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9036 5108 9088 5117
rect 12164 5244 12216 5296
rect 13728 5244 13780 5296
rect 16488 5244 16540 5296
rect 12900 5219 12952 5228
rect 12900 5185 12909 5219
rect 12909 5185 12943 5219
rect 12943 5185 12952 5219
rect 12900 5176 12952 5185
rect 14280 5176 14332 5228
rect 15108 5219 15160 5228
rect 15108 5185 15117 5219
rect 15117 5185 15151 5219
rect 15151 5185 15160 5219
rect 15108 5176 15160 5185
rect 13268 5108 13320 5160
rect 13452 5108 13504 5160
rect 2504 5040 2556 5092
rect 4804 5040 4856 5092
rect 11612 5040 11664 5092
rect 3056 4972 3108 5024
rect 4344 4972 4396 5024
rect 4436 4972 4488 5024
rect 4620 4972 4672 5024
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 7288 5015 7340 5024
rect 7288 4981 7297 5015
rect 7297 4981 7331 5015
rect 7331 4981 7340 5015
rect 7288 4972 7340 4981
rect 8208 4972 8260 5024
rect 8576 4972 8628 5024
rect 9128 4972 9180 5024
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 13544 5040 13596 5092
rect 14372 5108 14424 5160
rect 15660 5108 15712 5160
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 17316 5219 17368 5228
rect 17316 5185 17325 5219
rect 17325 5185 17359 5219
rect 17359 5185 17368 5219
rect 17316 5176 17368 5185
rect 16580 5108 16632 5160
rect 16764 5108 16816 5160
rect 16948 5108 17000 5160
rect 13176 4972 13228 5024
rect 14556 5015 14608 5024
rect 14556 4981 14565 5015
rect 14565 4981 14599 5015
rect 14599 4981 14608 5015
rect 14556 4972 14608 4981
rect 16488 5015 16540 5024
rect 16488 4981 16497 5015
rect 16497 4981 16531 5015
rect 16531 4981 16540 5015
rect 16488 4972 16540 4981
rect 16764 5015 16816 5024
rect 16764 4981 16773 5015
rect 16773 4981 16807 5015
rect 16807 4981 16816 5015
rect 16764 4972 16816 4981
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 2320 4768 2372 4820
rect 3148 4768 3200 4820
rect 4436 4811 4488 4820
rect 4436 4777 4445 4811
rect 4445 4777 4479 4811
rect 4479 4777 4488 4811
rect 4436 4768 4488 4777
rect 4712 4768 4764 4820
rect 5080 4768 5132 4820
rect 8392 4768 8444 4820
rect 8576 4768 8628 4820
rect 12164 4768 12216 4820
rect 13452 4768 13504 4820
rect 13728 4768 13780 4820
rect 1492 4675 1544 4684
rect 1492 4641 1501 4675
rect 1501 4641 1535 4675
rect 1535 4641 1544 4675
rect 1492 4632 1544 4641
rect 3884 4700 3936 4752
rect 3976 4700 4028 4752
rect 5632 4700 5684 4752
rect 6368 4700 6420 4752
rect 10416 4700 10468 4752
rect 11428 4700 11480 4752
rect 13544 4700 13596 4752
rect 14096 4700 14148 4752
rect 14372 4700 14424 4752
rect 2596 4632 2648 4684
rect 2688 4632 2740 4684
rect 5172 4632 5224 4684
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 5448 4632 5500 4641
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 6460 4632 6512 4641
rect 6920 4632 6972 4684
rect 8208 4632 8260 4684
rect 10508 4632 10560 4684
rect 12440 4632 12492 4684
rect 1952 4564 2004 4616
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 2964 4496 3016 4548
rect 3332 4496 3384 4548
rect 6000 4564 6052 4616
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 2596 4428 2648 4480
rect 3424 4428 3476 4480
rect 5632 4428 5684 4480
rect 9036 4428 9088 4480
rect 9312 4428 9364 4480
rect 12164 4564 12216 4616
rect 12808 4607 12860 4616
rect 12808 4573 12817 4607
rect 12817 4573 12851 4607
rect 12851 4573 12860 4607
rect 12808 4564 12860 4573
rect 14280 4632 14332 4684
rect 15384 4768 15436 4820
rect 15844 4768 15896 4820
rect 17960 4768 18012 4820
rect 16764 4700 16816 4752
rect 10784 4496 10836 4548
rect 11060 4428 11112 4480
rect 11796 4496 11848 4548
rect 13452 4496 13504 4548
rect 12716 4428 12768 4480
rect 15844 4564 15896 4616
rect 16672 4632 16724 4684
rect 15016 4496 15068 4548
rect 16856 4496 16908 4548
rect 17408 4496 17460 4548
rect 15108 4428 15160 4480
rect 17132 4471 17184 4480
rect 17132 4437 17141 4471
rect 17141 4437 17175 4471
rect 17175 4437 17184 4471
rect 17132 4428 17184 4437
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 6184 4224 6236 4276
rect 7012 4224 7064 4276
rect 7564 4224 7616 4276
rect 8208 4267 8260 4276
rect 2228 4088 2280 4140
rect 4712 4156 4764 4208
rect 1860 4063 1912 4072
rect 1860 4029 1869 4063
rect 1869 4029 1903 4063
rect 1903 4029 1912 4063
rect 1860 4020 1912 4029
rect 5448 4156 5500 4208
rect 6000 4156 6052 4208
rect 6644 4156 6696 4208
rect 8208 4233 8217 4267
rect 8217 4233 8251 4267
rect 8251 4233 8260 4267
rect 8208 4224 8260 4233
rect 8852 4224 8904 4276
rect 1400 3952 1452 4004
rect 4804 4020 4856 4072
rect 5448 4020 5500 4072
rect 6000 4020 6052 4072
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 10324 4199 10376 4208
rect 10324 4165 10333 4199
rect 10333 4165 10367 4199
rect 10367 4165 10376 4199
rect 10324 4156 10376 4165
rect 10232 4088 10284 4140
rect 10784 4020 10836 4072
rect 10876 4020 10928 4072
rect 1768 3884 1820 3936
rect 2412 3884 2464 3936
rect 2780 3884 2832 3936
rect 4712 3884 4764 3936
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 6460 3952 6512 4004
rect 6644 3952 6696 4004
rect 10508 3952 10560 4004
rect 11704 4156 11756 4208
rect 11796 4088 11848 4140
rect 12808 4224 12860 4276
rect 14004 4156 14056 4208
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 14280 4131 14332 4140
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 15108 4088 15160 4140
rect 17408 4088 17460 4140
rect 14556 4020 14608 4072
rect 15476 4063 15528 4072
rect 15476 4029 15510 4063
rect 15510 4029 15528 4063
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 5908 3884 5960 3936
rect 8392 3884 8444 3936
rect 9220 3884 9272 3936
rect 9496 3884 9548 3936
rect 10232 3884 10284 3936
rect 11520 3884 11572 3936
rect 12256 3952 12308 4004
rect 12532 3952 12584 4004
rect 15476 4020 15528 4029
rect 16488 4020 16540 4072
rect 17316 4020 17368 4072
rect 14924 3952 14976 4004
rect 17960 4020 18012 4072
rect 13636 3927 13688 3936
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 13636 3884 13688 3893
rect 14648 3884 14700 3936
rect 14740 3884 14792 3936
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 2504 3680 2556 3732
rect 6276 3680 6328 3732
rect 6460 3680 6512 3732
rect 7288 3723 7340 3732
rect 2412 3612 2464 3664
rect 4896 3612 4948 3664
rect 5172 3612 5224 3664
rect 6736 3612 6788 3664
rect 7288 3689 7297 3723
rect 7297 3689 7331 3723
rect 7331 3689 7340 3723
rect 7288 3680 7340 3689
rect 7932 3680 7984 3732
rect 8668 3723 8720 3732
rect 8668 3689 8677 3723
rect 8677 3689 8711 3723
rect 8711 3689 8720 3723
rect 8668 3680 8720 3689
rect 11428 3680 11480 3732
rect 7564 3612 7616 3664
rect 12072 3680 12124 3732
rect 12532 3680 12584 3732
rect 14280 3723 14332 3732
rect 388 3544 440 3596
rect 4160 3544 4212 3596
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 3056 3476 3108 3528
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 3240 3408 3292 3460
rect 5080 3476 5132 3528
rect 7380 3544 7432 3596
rect 6460 3476 6512 3528
rect 8300 3544 8352 3596
rect 11704 3612 11756 3664
rect 13176 3655 13228 3664
rect 13176 3621 13210 3655
rect 13210 3621 13228 3655
rect 13176 3612 13228 3621
rect 14280 3689 14289 3723
rect 14289 3689 14323 3723
rect 14323 3689 14332 3723
rect 14280 3680 14332 3689
rect 14832 3680 14884 3732
rect 17776 3680 17828 3732
rect 18052 3680 18104 3732
rect 18236 3723 18288 3732
rect 18236 3689 18245 3723
rect 18245 3689 18279 3723
rect 18279 3689 18288 3723
rect 18236 3680 18288 3689
rect 16672 3612 16724 3664
rect 8208 3476 8260 3528
rect 8484 3476 8536 3528
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 10784 3544 10836 3596
rect 11152 3544 11204 3596
rect 11336 3544 11388 3596
rect 13544 3544 13596 3596
rect 10508 3476 10560 3528
rect 10876 3519 10928 3528
rect 10876 3485 10885 3519
rect 10885 3485 10919 3519
rect 10919 3485 10928 3519
rect 10876 3476 10928 3485
rect 12716 3476 12768 3528
rect 14004 3476 14056 3528
rect 10232 3451 10284 3460
rect 10232 3417 10241 3451
rect 10241 3417 10275 3451
rect 10275 3417 10284 3451
rect 10232 3408 10284 3417
rect 14096 3408 14148 3460
rect 14924 3408 14976 3460
rect 1768 3340 1820 3392
rect 3332 3340 3384 3392
rect 4896 3340 4948 3392
rect 5448 3340 5500 3392
rect 6644 3383 6696 3392
rect 6644 3349 6653 3383
rect 6653 3349 6687 3383
rect 6687 3349 6696 3383
rect 6644 3340 6696 3349
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 9588 3340 9640 3392
rect 12900 3340 12952 3392
rect 13176 3340 13228 3392
rect 15660 3476 15712 3528
rect 16304 3476 16356 3528
rect 17408 3408 17460 3460
rect 16856 3340 16908 3392
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 5724 3068 5776 3120
rect 7840 3136 7892 3188
rect 11336 3136 11388 3188
rect 11980 3136 12032 3188
rect 16396 3136 16448 3188
rect 3976 3000 4028 3052
rect 4436 3000 4488 3052
rect 5448 3000 5500 3052
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 1216 2932 1268 2984
rect 4068 2932 4120 2984
rect 5632 2932 5684 2984
rect 6552 2932 6604 2984
rect 7748 3000 7800 3052
rect 10692 3000 10744 3052
rect 11796 3068 11848 3120
rect 11612 3000 11664 3052
rect 14740 3000 14792 3052
rect 15476 3000 15528 3052
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 17132 3000 17184 3052
rect 8484 2932 8536 2984
rect 8760 2932 8812 2984
rect 9312 2932 9364 2984
rect 2964 2864 3016 2916
rect 3516 2864 3568 2916
rect 3792 2864 3844 2916
rect 6368 2864 6420 2916
rect 11152 2932 11204 2984
rect 11520 2932 11572 2984
rect 12440 2932 12492 2984
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 15752 2932 15804 2984
rect 16120 2975 16172 2984
rect 16120 2941 16129 2975
rect 16129 2941 16163 2975
rect 16163 2941 16172 2975
rect 16120 2932 16172 2941
rect 16580 2932 16632 2984
rect 9496 2907 9548 2916
rect 9496 2873 9530 2907
rect 9530 2873 9548 2907
rect 9496 2864 9548 2873
rect 9680 2864 9732 2916
rect 1860 2839 1912 2848
rect 1860 2805 1869 2839
rect 1869 2805 1903 2839
rect 1903 2805 1912 2839
rect 1860 2796 1912 2805
rect 4068 2796 4120 2848
rect 4252 2839 4304 2848
rect 4252 2805 4261 2839
rect 4261 2805 4295 2839
rect 4295 2805 4304 2839
rect 4252 2796 4304 2805
rect 4988 2839 5040 2848
rect 4988 2805 4997 2839
rect 4997 2805 5031 2839
rect 5031 2805 5040 2839
rect 4988 2796 5040 2805
rect 5080 2796 5132 2848
rect 6000 2796 6052 2848
rect 6736 2796 6788 2848
rect 7380 2796 7432 2848
rect 8116 2796 8168 2848
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 11888 2796 11940 2848
rect 12716 2796 12768 2848
rect 13820 2796 13872 2848
rect 14004 2796 14056 2848
rect 14372 2796 14424 2848
rect 15660 2864 15712 2916
rect 16948 2864 17000 2916
rect 16764 2839 16816 2848
rect 16764 2805 16773 2839
rect 16773 2805 16807 2839
rect 16807 2805 16816 2839
rect 16764 2796 16816 2805
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 2964 2635 3016 2644
rect 2964 2601 2973 2635
rect 2973 2601 3007 2635
rect 3007 2601 3016 2635
rect 2964 2592 3016 2601
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 4252 2592 4304 2644
rect 4988 2635 5040 2644
rect 4988 2601 4997 2635
rect 4997 2601 5031 2635
rect 5031 2601 5040 2635
rect 4988 2592 5040 2601
rect 5724 2592 5776 2644
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 9680 2592 9732 2644
rect 9772 2592 9824 2644
rect 10232 2592 10284 2644
rect 10968 2592 11020 2644
rect 11428 2592 11480 2644
rect 12256 2592 12308 2644
rect 13636 2635 13688 2644
rect 13636 2601 13645 2635
rect 13645 2601 13679 2635
rect 13679 2601 13688 2635
rect 13636 2592 13688 2601
rect 13728 2592 13780 2644
rect 15660 2635 15712 2644
rect 15660 2601 15669 2635
rect 15669 2601 15703 2635
rect 15703 2601 15712 2635
rect 15660 2592 15712 2601
rect 15752 2592 15804 2644
rect 16764 2592 16816 2644
rect 2688 2524 2740 2576
rect 2780 2524 2832 2576
rect 4896 2567 4948 2576
rect 4896 2533 4905 2567
rect 4905 2533 4939 2567
rect 4939 2533 4948 2567
rect 4896 2524 4948 2533
rect 5080 2524 5132 2576
rect 10876 2524 10928 2576
rect 13820 2524 13872 2576
rect 15568 2524 15620 2576
rect 16120 2567 16172 2576
rect 16120 2533 16129 2567
rect 16129 2533 16163 2567
rect 16163 2533 16172 2567
rect 16120 2524 16172 2533
rect 16856 2524 16908 2576
rect 3608 2456 3660 2508
rect 5356 2456 5408 2508
rect 7932 2499 7984 2508
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 3976 2388 4028 2440
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 7472 2431 7524 2440
rect 6368 2388 6420 2397
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 7932 2465 7941 2499
rect 7941 2465 7975 2499
rect 7975 2465 7984 2499
rect 7932 2456 7984 2465
rect 11704 2456 11756 2508
rect 13452 2456 13504 2508
rect 8300 2388 8352 2440
rect 10140 2388 10192 2440
rect 10692 2388 10744 2440
rect 12348 2388 12400 2440
rect 13084 2431 13136 2440
rect 13084 2397 13093 2431
rect 13093 2397 13127 2431
rect 13127 2397 13136 2431
rect 13084 2388 13136 2397
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 15476 2456 15528 2508
rect 16304 2431 16356 2440
rect 16304 2397 16313 2431
rect 16313 2397 16347 2431
rect 16347 2397 16356 2431
rect 16304 2388 16356 2397
rect 2780 2252 2832 2304
rect 8484 2252 8536 2304
rect 14004 2252 14056 2304
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 13084 2048 13136 2100
rect 14188 2048 14240 2100
rect 3240 1844 3292 1896
rect 5908 1844 5960 1896
rect 2044 1300 2096 1352
rect 15200 1300 15252 1352
<< metal2 >>
rect 1582 16552 1638 16561
rect 1582 16487 1638 16496
rect 1490 15192 1546 15201
rect 1490 15127 1546 15136
rect 1504 13530 1532 15127
rect 1596 14618 1624 16487
rect 1950 16200 2006 17000
rect 4066 16824 4122 16833
rect 4066 16759 4122 16768
rect 1674 14920 1730 14929
rect 1674 14855 1730 14864
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1596 13870 1624 14554
rect 1688 13938 1716 14855
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1780 14249 1808 14350
rect 1766 14240 1822 14249
rect 1766 14175 1822 14184
rect 1964 14006 1992 16200
rect 2870 16144 2926 16153
rect 2870 16079 2926 16088
rect 2778 14512 2834 14521
rect 2778 14447 2834 14456
rect 1952 14000 2004 14006
rect 1952 13942 2004 13948
rect 2792 13938 2820 14447
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2884 13870 2912 16079
rect 3974 15872 4030 15881
rect 3974 15807 4030 15816
rect 2962 15464 3018 15473
rect 2962 15399 3018 15408
rect 2976 14482 3004 15399
rect 3988 15230 4016 15807
rect 4080 15298 4108 16759
rect 5906 16200 5962 17000
rect 9862 16200 9918 17000
rect 13910 16200 13966 17000
rect 15474 16552 15530 16561
rect 15474 16487 15530 16496
rect 4068 15292 4120 15298
rect 4068 15234 4120 15240
rect 3976 15224 4028 15230
rect 3976 15166 4028 15172
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 5920 14074 5948 16200
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 1584 13864 1636 13870
rect 2872 13864 2924 13870
rect 1584 13806 1636 13812
rect 1766 13832 1822 13841
rect 2872 13806 2924 13812
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 1766 13767 1822 13776
rect 1492 13524 1544 13530
rect 1492 13466 1544 13472
rect 1504 12782 1532 13466
rect 1780 12850 1808 13767
rect 2778 13560 2834 13569
rect 2778 13495 2834 13504
rect 2792 13394 2820 13495
rect 2884 13462 2912 13806
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2778 13288 2834 13297
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10130 1440 11154
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1688 10606 1716 11086
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1964 9518 1992 10066
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1124 8832 1176 8838
rect 1124 8774 1176 8780
rect 1136 4457 1164 8774
rect 1596 5409 1624 9318
rect 1674 9072 1730 9081
rect 1964 9042 1992 9454
rect 1674 9007 1730 9016
rect 1952 9036 2004 9042
rect 1688 8430 1716 9007
rect 1952 8978 2004 8984
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1766 7984 1822 7993
rect 1766 7919 1822 7928
rect 1780 5846 1808 7919
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1964 7002 1992 7686
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1950 6760 2006 6769
rect 1950 6695 2006 6704
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1582 5400 1638 5409
rect 1582 5335 1638 5344
rect 1400 5092 1452 5098
rect 1400 5034 1452 5040
rect 1122 4448 1178 4457
rect 1122 4383 1178 4392
rect 1412 4010 1440 5034
rect 1490 4856 1546 4865
rect 1490 4791 1546 4800
rect 1504 4690 1532 4791
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1964 4622 1992 6695
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1858 4176 1914 4185
rect 1858 4111 1914 4120
rect 1872 4078 1900 4111
rect 1860 4072 1912 4078
rect 1490 4040 1546 4049
rect 1400 4004 1452 4010
rect 1860 4014 1912 4020
rect 1490 3975 1546 3984
rect 1400 3946 1452 3952
rect 388 3596 440 3602
rect 388 3538 440 3544
rect 400 800 428 3538
rect 1412 3534 1440 3946
rect 1504 3777 1532 3975
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1490 3768 1546 3777
rect 1490 3703 1546 3712
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1780 3398 1808 3878
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1216 2984 1268 2990
rect 1216 2926 1268 2932
rect 1858 2952 1914 2961
rect 1228 800 1256 2926
rect 1858 2887 1914 2896
rect 1872 2854 1900 2887
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 2056 1358 2084 13262
rect 2778 13223 2780 13232
rect 2832 13223 2834 13232
rect 2780 13194 2832 13200
rect 3252 12889 3280 13738
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3238 12880 3294 12889
rect 3238 12815 3294 12824
rect 3332 12844 3384 12850
rect 2594 12336 2650 12345
rect 2228 12300 2280 12306
rect 2594 12271 2650 12280
rect 2228 12242 2280 12248
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2148 11898 2176 12174
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2240 10810 2268 12242
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2332 10198 2360 11290
rect 2424 11218 2452 11562
rect 2608 11558 2636 12271
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2700 11626 2728 12174
rect 3160 11898 3188 12174
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3252 11830 3280 12815
rect 3332 12786 3384 12792
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2700 11354 2728 11562
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2424 10674 2452 11154
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2778 10024 2834 10033
rect 2778 9959 2834 9968
rect 2686 9208 2742 9217
rect 2136 9172 2188 9178
rect 2686 9143 2742 9152
rect 2136 9114 2188 9120
rect 2148 4128 2176 9114
rect 2700 9042 2728 9143
rect 2688 9036 2740 9042
rect 2608 8996 2688 9024
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2320 8424 2372 8430
rect 2424 8412 2452 8910
rect 2372 8384 2452 8412
rect 2320 8366 2372 8372
rect 2608 8362 2636 8996
rect 2688 8978 2740 8984
rect 2596 8356 2648 8362
rect 2596 8298 2648 8304
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2332 7410 2360 7754
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2240 6458 2268 7142
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2240 5098 2268 6258
rect 2332 5914 2360 7142
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2228 5092 2280 5098
rect 2228 5034 2280 5040
rect 2332 4826 2360 5646
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2228 4140 2280 4146
rect 2148 4100 2228 4128
rect 2228 4082 2280 4088
rect 2240 3641 2268 4082
rect 2424 3942 2452 8230
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2516 7546 2544 7822
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2792 7460 2820 9959
rect 2608 7432 2820 7460
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 6390 2544 6598
rect 2608 6497 2636 7432
rect 2884 7392 2912 10474
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2976 9518 3004 10202
rect 3054 10160 3110 10169
rect 3054 10095 3056 10104
rect 3108 10095 3110 10104
rect 3056 10066 3108 10072
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2976 8294 3004 8978
rect 3068 8945 3096 9454
rect 3054 8936 3110 8945
rect 3054 8871 3110 8880
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 3068 7970 3096 8230
rect 2792 7364 2912 7392
rect 2976 7942 3096 7970
rect 2686 6760 2742 6769
rect 2686 6695 2742 6704
rect 2594 6488 2650 6497
rect 2594 6423 2650 6432
rect 2504 6384 2556 6390
rect 2504 6326 2556 6332
rect 2608 6254 2636 6423
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2700 5642 2728 6695
rect 2792 5681 2820 7364
rect 2872 7268 2924 7274
rect 2872 7210 2924 7216
rect 2884 6769 2912 7210
rect 2976 7206 3004 7942
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3068 7410 3096 7822
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2870 6760 2926 6769
rect 2870 6695 2926 6704
rect 2976 6186 3004 6802
rect 3068 6730 3096 7346
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3068 6254 3096 6666
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 3056 6112 3108 6118
rect 3160 6089 3188 9862
rect 3344 9738 3372 12786
rect 3804 12617 3832 13126
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 3790 12608 3846 12617
rect 3790 12543 3846 12552
rect 4068 12368 4120 12374
rect 3698 12336 3754 12345
rect 4068 12310 4120 12316
rect 3698 12271 3754 12280
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3436 10266 3464 12174
rect 3606 11928 3662 11937
rect 3606 11863 3662 11872
rect 3620 11830 3648 11863
rect 3608 11824 3660 11830
rect 3608 11766 3660 11772
rect 3620 11642 3648 11766
rect 3528 11614 3648 11642
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3252 9710 3372 9738
rect 3252 8634 3280 9710
rect 3528 9602 3556 11614
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 10810 3648 11494
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3528 9574 3648 9602
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 9110 3372 9318
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3344 8498 3372 9046
rect 3528 8945 3556 9386
rect 3514 8936 3570 8945
rect 3514 8871 3570 8880
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3056 6054 3108 6060
rect 3146 6080 3202 6089
rect 2884 5914 2912 6054
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 3068 5710 3096 6054
rect 3146 6015 3202 6024
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3056 5704 3108 5710
rect 2778 5672 2834 5681
rect 2688 5636 2740 5642
rect 3056 5646 3108 5652
rect 2778 5607 2834 5616
rect 2872 5636 2924 5642
rect 2688 5578 2740 5584
rect 2872 5578 2924 5584
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2516 5098 2544 5510
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2424 3670 2452 3878
rect 2516 3738 2544 5034
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2608 4486 2636 4626
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2412 3664 2464 3670
rect 2226 3632 2282 3641
rect 2412 3606 2464 3612
rect 2226 3567 2282 3576
rect 2700 2689 2728 4626
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2686 2680 2742 2689
rect 2686 2615 2742 2624
rect 2700 2582 2728 2615
rect 2792 2582 2820 3878
rect 2884 3505 2912 5578
rect 3068 5370 3096 5646
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 3068 4706 3096 4966
rect 3160 4826 3188 5714
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3068 4678 3188 4706
rect 3056 4616 3108 4622
rect 3054 4584 3056 4593
rect 3108 4584 3110 4593
rect 2964 4548 3016 4554
rect 3054 4519 3110 4528
rect 2964 4490 3016 4496
rect 2870 3496 2926 3505
rect 2870 3431 2926 3440
rect 2976 3346 3004 4490
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2884 3318 3004 3346
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 2044 1352 2096 1358
rect 2044 1294 2096 1300
rect 2148 800 2176 2382
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 386 0 442 800
rect 1214 0 1270 800
rect 2134 0 2190 800
rect 2792 241 2820 2246
rect 2884 785 2912 3318
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2976 2650 3004 2858
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3068 800 3096 3470
rect 3160 1193 3188 4678
rect 3252 4049 3280 8298
rect 3528 8090 3556 8871
rect 3620 8294 3648 9574
rect 3712 9042 3740 12271
rect 4080 12209 4108 12310
rect 5816 12232 5868 12238
rect 4066 12200 4122 12209
rect 5816 12174 5868 12180
rect 4066 12135 4122 12144
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 4632 11898 4660 12038
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4802 11792 4858 11801
rect 4802 11727 4858 11736
rect 5264 11756 5316 11762
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4080 11257 4108 11494
rect 4066 11248 4122 11257
rect 4066 11183 4122 11192
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10742 3832 10950
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3896 10266 3924 10406
rect 4066 10296 4122 10305
rect 3884 10260 3936 10266
rect 4066 10231 4122 10240
rect 3884 10202 3936 10208
rect 4080 10198 4108 10231
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 4066 9480 4122 9489
rect 4066 9415 4122 9424
rect 4080 9382 4108 9415
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3804 8974 3832 9318
rect 4264 9217 4292 10746
rect 4618 10704 4674 10713
rect 4724 10674 4752 11154
rect 4618 10639 4674 10648
rect 4712 10668 4764 10674
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4540 9518 4568 9862
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4436 9376 4488 9382
rect 4488 9336 4568 9364
rect 4436 9318 4488 9324
rect 4250 9208 4306 9217
rect 4250 9143 4306 9152
rect 4436 9104 4488 9110
rect 4436 9046 4488 9052
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 4356 8566 4384 8978
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 4264 7993 4292 8298
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4250 7984 4306 7993
rect 4250 7919 4306 7928
rect 4356 7936 4384 8230
rect 4448 8090 4476 9046
rect 4540 8809 4568 9336
rect 4632 9178 4660 10639
rect 4712 10610 4764 10616
rect 4724 9994 4752 10610
rect 4816 10470 4844 11727
rect 5264 11698 5316 11704
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 5092 11257 5120 11630
rect 5078 11248 5134 11257
rect 5078 11183 5134 11192
rect 4894 11112 4950 11121
rect 4894 11047 4950 11056
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4724 9722 4752 9930
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4526 8800 4582 8809
rect 4526 8735 4582 8744
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4356 7908 4476 7936
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3436 7410 3464 7754
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3436 6934 3464 7346
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3344 6225 3372 6802
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3436 6361 3464 6394
rect 3422 6352 3478 6361
rect 3422 6287 3478 6296
rect 3330 6216 3386 6225
rect 3330 6151 3386 6160
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3344 4554 3372 5510
rect 3332 4548 3384 4554
rect 3332 4490 3384 4496
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3238 4040 3294 4049
rect 3238 3975 3294 3984
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 3252 2825 3280 3402
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3238 2816 3294 2825
rect 3238 2751 3294 2760
rect 3344 2650 3372 3334
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3240 1896 3292 1902
rect 3238 1864 3240 1873
rect 3292 1864 3294 1873
rect 3238 1799 3294 1808
rect 3146 1184 3202 1193
rect 3146 1119 3202 1128
rect 2870 776 2926 785
rect 2870 711 2926 720
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 3054 0 3110 800
rect 3436 513 3464 4422
rect 3528 3233 3556 7686
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3712 7313 3740 7482
rect 3698 7304 3754 7313
rect 3698 7239 3754 7248
rect 3804 6905 3832 7822
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4448 7426 4476 7908
rect 4540 7546 4568 8230
rect 4632 7886 4660 8434
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4724 7546 4752 9658
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 3790 6896 3846 6905
rect 3790 6831 3846 6840
rect 4066 6896 4122 6905
rect 4066 6831 4068 6840
rect 4120 6831 4122 6840
rect 4068 6802 4120 6808
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 6254 3648 6598
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 3514 3224 3570 3233
rect 3514 3159 3570 3168
rect 3514 3088 3570 3097
rect 3514 3023 3570 3032
rect 3528 2922 3556 3023
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3620 2514 3648 5578
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 3712 2145 3740 6666
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 3108 3832 6598
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3988 5642 4016 5850
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3896 4758 3924 5238
rect 4264 5137 4292 5782
rect 4356 5778 4384 7414
rect 4448 7398 4752 7426
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4448 5914 4476 6938
rect 4540 6798 4568 7278
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6254 4568 6734
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4434 5808 4490 5817
rect 4344 5772 4396 5778
rect 4434 5743 4490 5752
rect 4344 5714 4396 5720
rect 4448 5234 4476 5743
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4250 5128 4306 5137
rect 4250 5063 4306 5072
rect 4448 5030 4476 5170
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 3884 4752 3936 4758
rect 3976 4752 4028 4758
rect 3884 4694 3936 4700
rect 3974 4720 3976 4729
rect 4028 4720 4030 4729
rect 3974 4655 4030 4664
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4172 3380 4200 3538
rect 4172 3352 4292 3380
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 3804 3080 3924 3108
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 3698 2136 3754 2145
rect 3698 2071 3754 2080
rect 3804 1442 3832 2858
rect 3896 2417 3924 3080
rect 4066 3088 4122 3097
rect 3976 3052 4028 3058
rect 4066 3023 4122 3032
rect 3976 2994 4028 3000
rect 3988 2446 4016 2994
rect 4080 2990 4108 3023
rect 4068 2984 4120 2990
rect 4264 2938 4292 3352
rect 4068 2926 4120 2932
rect 4172 2910 4292 2938
rect 4068 2848 4120 2854
rect 4172 2836 4200 2910
rect 4120 2808 4200 2836
rect 4252 2848 4304 2854
rect 4068 2790 4120 2796
rect 4252 2790 4304 2796
rect 4264 2650 4292 2790
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 3976 2440 4028 2446
rect 3882 2408 3938 2417
rect 3976 2382 4028 2388
rect 3882 2343 3938 2352
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 4356 1578 4384 4966
rect 4434 4856 4490 4865
rect 4434 4791 4436 4800
rect 4488 4791 4490 4800
rect 4436 4762 4488 4768
rect 4540 3913 4568 6054
rect 4632 5710 4660 6122
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4724 5642 4752 7398
rect 4816 5817 4844 10406
rect 4908 10062 4936 11047
rect 5276 10849 5304 11698
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5262 10840 5318 10849
rect 5368 10810 5396 11562
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5262 10775 5264 10784
rect 5316 10775 5318 10784
rect 5356 10804 5408 10810
rect 5264 10746 5316 10752
rect 5356 10746 5408 10752
rect 5276 10715 5304 10746
rect 5460 10674 5488 11018
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5080 10124 5132 10130
rect 5000 10084 5080 10112
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4908 7041 4936 9998
rect 4894 7032 4950 7041
rect 5000 7018 5028 10084
rect 5080 10066 5132 10072
rect 5368 9897 5396 10474
rect 5552 10266 5580 10542
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5354 9888 5410 9897
rect 5354 9823 5410 9832
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5092 8838 5120 9454
rect 5368 8888 5396 9823
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5460 9178 5488 9386
rect 5552 9382 5580 10066
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5368 8860 5488 8888
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5354 8800 5410 8809
rect 5092 7954 5120 8774
rect 5354 8735 5410 8744
rect 5368 8294 5396 8735
rect 5264 8288 5316 8294
rect 5262 8256 5264 8265
rect 5356 8288 5408 8294
rect 5316 8256 5318 8265
rect 5184 8214 5262 8242
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5000 6990 5120 7018
rect 4894 6967 4950 6976
rect 4802 5808 4858 5817
rect 4908 5778 4936 6967
rect 4988 5908 5040 5914
rect 5092 5896 5120 6990
rect 5040 5868 5120 5896
rect 4988 5850 5040 5856
rect 4802 5743 4858 5752
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4632 5137 4660 5170
rect 4618 5128 4674 5137
rect 4618 5063 4674 5072
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4632 4298 4660 4966
rect 4724 4826 4752 5578
rect 4816 5574 4844 5646
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4816 5098 4844 5510
rect 5000 5370 5028 5850
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 5092 4826 5120 5510
rect 5184 5250 5212 8214
rect 5356 8230 5408 8236
rect 5262 8191 5318 8200
rect 5368 5710 5396 8230
rect 5460 7857 5488 8860
rect 5446 7848 5502 7857
rect 5446 7783 5502 7792
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5368 5250 5396 5306
rect 5184 5222 5396 5250
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5184 4690 5212 5222
rect 5262 5128 5318 5137
rect 5262 5063 5318 5072
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5276 4570 5304 5063
rect 5460 4690 5488 7783
rect 5552 6934 5580 9318
rect 5644 7290 5672 12106
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5736 11354 5764 11494
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5828 11218 5856 12174
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 6012 11665 6040 11766
rect 5998 11656 6054 11665
rect 5998 11591 6054 11600
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5722 10704 5778 10713
rect 5722 10639 5778 10648
rect 5736 10538 5764 10639
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5736 10441 5764 10474
rect 5722 10432 5778 10441
rect 5722 10367 5778 10376
rect 5828 10130 5856 11154
rect 5998 10704 6054 10713
rect 5998 10639 6054 10648
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5920 9489 5948 10542
rect 6012 10266 6040 10639
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5906 9480 5962 9489
rect 5906 9415 5962 9424
rect 6012 8430 6040 10202
rect 6000 8424 6052 8430
rect 5814 8392 5870 8401
rect 6000 8366 6052 8372
rect 5814 8327 5870 8336
rect 5644 7262 5764 7290
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5448 4684 5500 4690
rect 5092 4542 5304 4570
rect 5368 4644 5448 4672
rect 4632 4270 4752 4298
rect 4724 4214 4752 4270
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4712 3936 4764 3942
rect 4526 3904 4582 3913
rect 4526 3839 4582 3848
rect 4710 3904 4712 3913
rect 4764 3904 4766 3913
rect 4710 3839 4766 3848
rect 4816 3534 4844 4014
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3670 4936 3878
rect 5092 3777 5120 4542
rect 5078 3768 5134 3777
rect 5078 3703 5134 3712
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4986 3632 5042 3641
rect 4986 3567 5042 3576
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4434 3224 4490 3233
rect 4434 3159 4490 3168
rect 4448 3058 4476 3159
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4908 2582 4936 3334
rect 5000 2938 5028 3567
rect 5092 3534 5120 3703
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5000 2910 5120 2938
rect 5092 2854 5120 2910
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5000 2650 5028 2790
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 4080 1550 4384 1578
rect 4080 1465 4108 1550
rect 4066 1456 4122 1465
rect 3804 1414 4016 1442
rect 3988 800 4016 1414
rect 4066 1391 4122 1400
rect 5092 1306 5120 2518
rect 5184 2446 5212 3606
rect 5368 2514 5396 4644
rect 5448 4626 5500 4632
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5460 4078 5488 4150
rect 5448 4072 5500 4078
rect 5552 4049 5580 6258
rect 5644 4758 5672 7142
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5448 4014 5500 4020
rect 5538 4040 5594 4049
rect 5460 3754 5488 4014
rect 5538 3975 5594 3984
rect 5552 3942 5580 3975
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5460 3726 5580 3754
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 3058 5488 3334
rect 5552 3058 5580 3726
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5644 2990 5672 4422
rect 5736 3369 5764 7262
rect 5828 6322 5856 8327
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5920 5778 5948 6054
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5722 3360 5778 3369
rect 5722 3295 5778 3304
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5736 2650 5764 3062
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 4908 1278 5120 1306
rect 4908 800 4936 1278
rect 5828 800 5856 5646
rect 5920 5234 5948 5714
rect 6012 5574 6040 6598
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4622 6040 4966
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6012 4214 6040 4558
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5908 3936 5960 3942
rect 6012 3913 6040 4014
rect 5908 3878 5960 3884
rect 5998 3904 6054 3913
rect 5920 1902 5948 3878
rect 5998 3839 6054 3848
rect 6012 2854 6040 3839
rect 6104 3641 6132 13806
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7116 12714 7144 13194
rect 7392 12850 7512 12866
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7392 12844 7524 12850
rect 7392 12838 7472 12844
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7208 12628 7236 12786
rect 7208 12600 7328 12628
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 7300 12442 7328 12600
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7392 12170 7420 12838
rect 7472 12786 7524 12792
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 6274 12064 6330 12073
rect 6274 11999 6330 12008
rect 6288 11694 6316 11999
rect 6932 11762 6960 12106
rect 7378 12064 7434 12073
rect 7378 11999 7434 12008
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6380 11286 6408 11698
rect 7392 11694 7420 11999
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6196 10062 6224 10202
rect 6288 10130 6316 10678
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6288 9586 6316 10066
rect 6380 9994 6408 10610
rect 6458 10568 6514 10577
rect 6458 10503 6514 10512
rect 6552 10532 6604 10538
rect 6472 10033 6500 10503
rect 6552 10474 6604 10480
rect 6458 10024 6514 10033
rect 6368 9988 6420 9994
rect 6458 9959 6514 9968
rect 6368 9930 6420 9936
rect 6564 9761 6592 10474
rect 6656 10248 6684 11562
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 6920 11144 6972 11150
rect 7300 11121 7328 11562
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 6920 11086 6972 11092
rect 7286 11112 7342 11121
rect 6932 10742 6960 11086
rect 7286 11047 7342 11056
rect 7102 10840 7158 10849
rect 7102 10775 7158 10784
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 7116 10674 7144 10775
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 6736 10260 6788 10266
rect 6656 10220 6736 10248
rect 6736 10202 6788 10208
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 6550 9752 6606 9761
rect 6932 9722 6960 10134
rect 6550 9687 6606 9696
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 9042 6316 9522
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 7300 9178 7328 10542
rect 7392 9625 7420 11154
rect 7484 10198 7512 11698
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7576 10674 7604 11018
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7378 9616 7434 9625
rect 7378 9551 7434 9560
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7392 9353 7420 9454
rect 7378 9344 7434 9353
rect 7378 9279 7434 9288
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6288 8498 6316 8978
rect 6736 8560 6788 8566
rect 6366 8528 6422 8537
rect 6276 8492 6328 8498
rect 6736 8502 6788 8508
rect 6366 8463 6422 8472
rect 6644 8492 6696 8498
rect 6276 8434 6328 8440
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6196 6458 6224 8230
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6288 7002 6316 7346
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6184 5772 6236 5778
rect 6288 5760 6316 6394
rect 6380 5778 6408 8463
rect 6644 8434 6696 8440
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6472 7002 6500 8298
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 8022 6592 8230
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6656 7886 6684 8434
rect 6748 8022 6776 8502
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6472 5817 6500 6190
rect 6458 5808 6514 5817
rect 6236 5732 6316 5760
rect 6368 5772 6420 5778
rect 6184 5714 6236 5720
rect 6458 5743 6514 5752
rect 6368 5714 6420 5720
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6090 3632 6146 3641
rect 6090 3567 6146 3576
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6196 2428 6224 4218
rect 6288 3738 6316 4966
rect 6368 4752 6420 4758
rect 6368 4694 6420 4700
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6380 2922 6408 4694
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6472 4010 6500 4626
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6458 3768 6514 3777
rect 6458 3703 6460 3712
rect 6512 3703 6514 3712
rect 6460 3674 6512 3680
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6368 2916 6420 2922
rect 6368 2858 6420 2864
rect 6472 2689 6500 3470
rect 6564 2990 6592 7142
rect 6748 6905 6776 7210
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 7300 6984 7328 7142
rect 7208 6956 7328 6984
rect 6734 6896 6790 6905
rect 6734 6831 6790 6840
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6656 5914 6684 6734
rect 7208 6662 7236 6956
rect 7392 6916 7420 7890
rect 7300 6888 7420 6916
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6642 5672 6698 5681
rect 6642 5607 6698 5616
rect 6656 4214 6684 5607
rect 6748 4808 6776 6054
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7208 5250 7236 5510
rect 7300 5409 7328 6888
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7286 5400 7342 5409
rect 7392 5370 7420 6666
rect 7484 6458 7512 9930
rect 7576 9042 7604 10610
rect 7668 10441 7696 11766
rect 7760 10470 7788 14418
rect 9876 14362 9904 16200
rect 10508 15292 10560 15298
rect 10508 15234 10560 15240
rect 9784 14334 9904 14362
rect 9784 14006 9812 14334
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 12481 7880 12582
rect 7838 12472 7894 12481
rect 7838 12407 7894 12416
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7748 10464 7800 10470
rect 7654 10432 7710 10441
rect 7748 10406 7800 10412
rect 7654 10367 7710 10376
rect 7852 10282 7880 12174
rect 7760 10254 7880 10282
rect 7760 9874 7788 10254
rect 7668 9846 7788 9874
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7668 8090 7696 9846
rect 7838 9752 7894 9761
rect 7838 9687 7894 9696
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7760 7750 7788 9386
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7576 7002 7604 7210
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7562 6896 7618 6905
rect 7562 6831 7618 6840
rect 7576 6662 7604 6831
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7484 5710 7512 6122
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7286 5335 7342 5344
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7208 5222 7420 5250
rect 7484 5234 7512 5646
rect 7576 5574 7604 6598
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7562 5400 7618 5409
rect 7562 5335 7618 5344
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 6748 4780 6960 4808
rect 6932 4690 6960 4780
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6656 3398 6684 3946
rect 6748 3670 6776 4558
rect 6932 4298 6960 4626
rect 6932 4282 7052 4298
rect 6932 4276 7064 4282
rect 6932 4270 7012 4276
rect 6828 4072 6880 4078
rect 6932 4026 6960 4270
rect 7012 4218 7064 4224
rect 6880 4020 6960 4026
rect 6828 4014 6960 4020
rect 6840 3998 6960 4014
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 7300 3738 7328 4966
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 7392 3602 7420 5222
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7576 5114 7604 5335
rect 7484 5086 7604 5114
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 6458 2680 6514 2689
rect 6458 2615 6514 2624
rect 6368 2440 6420 2446
rect 6196 2400 6368 2428
rect 6368 2382 6420 2388
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 6748 800 6776 2790
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 7392 2650 7420 2790
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7484 2446 7512 5086
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7576 3670 7604 4218
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7668 3516 7696 7210
rect 7576 3488 7696 3516
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7576 800 7604 3488
rect 7760 3058 7788 7686
rect 7852 7478 7880 9687
rect 7944 9178 7972 12718
rect 8022 11792 8078 11801
rect 8022 11727 8024 11736
rect 8076 11727 8078 11736
rect 8024 11698 8076 11704
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 11218 8064 11494
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 9178 8064 10406
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8128 8956 8156 12786
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8220 12073 8248 12582
rect 8206 12064 8262 12073
rect 8206 11999 8262 12008
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8220 9926 8248 11630
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8206 9752 8262 9761
rect 8206 9687 8262 9696
rect 8036 8928 8156 8956
rect 8036 7954 8064 8928
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8128 8362 8156 8774
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7852 3194 7880 7278
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 8036 6882 8064 7346
rect 8128 7002 8156 8298
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8220 6882 8248 9687
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8312 8634 8340 8978
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8404 8090 8432 12922
rect 8864 12918 8892 13126
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8496 10198 8524 12718
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 11762 8616 12242
rect 8666 11928 8722 11937
rect 8666 11863 8722 11872
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8680 11694 8708 11863
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8588 11014 8616 11562
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8666 10840 8722 10849
rect 8666 10775 8722 10784
rect 8574 10432 8630 10441
rect 8574 10367 8630 10376
rect 8588 10198 8616 10367
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9518 8616 9998
rect 8576 9512 8628 9518
rect 8482 9480 8538 9489
rect 8576 9454 8628 9460
rect 8482 9415 8538 9424
rect 8496 8090 8524 9415
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8588 8673 8616 9046
rect 8680 8974 8708 10775
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8574 8664 8630 8673
rect 8574 8599 8630 8608
rect 8576 8560 8628 8566
rect 8574 8528 8576 8537
rect 8628 8528 8630 8537
rect 8574 8463 8630 8472
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 7002 8432 7754
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 7944 5370 7972 6870
rect 8036 6854 8156 6882
rect 8220 6854 8340 6882
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8036 5914 8064 6734
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 8036 4672 8064 5510
rect 8128 5386 8156 6854
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8220 6458 8248 6666
rect 8312 6458 8340 6854
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8404 6338 8432 6938
rect 8588 6730 8616 8298
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8312 6310 8432 6338
rect 8220 5574 8248 6258
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8128 5358 8248 5386
rect 8220 5030 8248 5358
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8208 4684 8260 4690
rect 8036 4644 8156 4672
rect 7930 4584 7986 4593
rect 7930 4519 7986 4528
rect 7944 3738 7972 4519
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7930 3360 7986 3369
rect 7930 3295 7986 3304
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7944 2514 7972 3295
rect 8128 2854 8156 4644
rect 8208 4626 8260 4632
rect 8220 4282 8248 4626
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8220 3534 8248 4218
rect 8312 3602 8340 6310
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8496 6118 8524 6149
rect 8484 6112 8536 6118
rect 8482 6080 8484 6089
rect 8536 6080 8538 6089
rect 8482 6015 8538 6024
rect 8496 5710 8524 6015
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8404 4826 8432 5170
rect 8588 5166 8616 6190
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8588 4826 8616 4966
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8312 2446 8340 3334
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8404 2122 8432 3878
rect 8680 3738 8708 8366
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8496 2990 8524 3470
rect 8772 2990 8800 12854
rect 8850 12472 8906 12481
rect 8956 12442 8984 13126
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 8850 12407 8906 12416
rect 8944 12436 8996 12442
rect 8864 11898 8892 12407
rect 8944 12378 8996 12384
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8956 11898 8984 12174
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 9722 8892 10406
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8956 9178 8984 11494
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8864 7886 8892 8910
rect 8956 8809 8984 8910
rect 8942 8800 8998 8809
rect 8942 8735 8998 8744
rect 9048 8634 9076 12582
rect 9324 12442 9352 12582
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9140 9994 9168 12242
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11354 9260 11494
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 9140 9722 9168 9930
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 8294 8984 8434
rect 9036 8424 9088 8430
rect 9034 8392 9036 8401
rect 9088 8392 9090 8401
rect 9034 8327 9090 8336
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 9140 8106 9168 9114
rect 8956 8078 9168 8106
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8852 6792 8904 6798
rect 8956 6769 8984 8078
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9048 7002 9076 7210
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8852 6734 8904 6740
rect 8942 6760 8998 6769
rect 8864 4593 8892 6734
rect 8942 6695 8998 6704
rect 8956 5846 8984 6695
rect 9140 6361 9168 7278
rect 9232 6934 9260 11086
rect 9416 11082 9444 12174
rect 9508 11150 9536 13670
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12442 9720 12582
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9680 11824 9732 11830
rect 9586 11792 9642 11801
rect 9680 11766 9732 11772
rect 9586 11727 9642 11736
rect 9600 11558 9628 11727
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 9568 9444 11018
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9508 10470 9536 10678
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9508 9897 9536 9930
rect 9494 9888 9550 9897
rect 9494 9823 9550 9832
rect 9600 9568 9628 10746
rect 9692 10674 9720 11766
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9692 10266 9720 10406
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9315 9540 9444 9568
rect 9499 9540 9628 9568
rect 9315 9450 9343 9540
rect 9312 9444 9364 9450
rect 9499 9432 9527 9540
rect 9499 9404 9536 9432
rect 9312 9386 9364 9392
rect 9508 9092 9536 9404
rect 9588 9376 9640 9382
rect 9586 9344 9588 9353
rect 9640 9344 9642 9353
rect 9586 9279 9642 9288
rect 9692 9178 9720 10066
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 9104 9640 9110
rect 9508 9064 9588 9092
rect 9588 9046 9640 9052
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9126 6352 9182 6361
rect 9126 6287 9182 6296
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 8850 4584 8906 4593
rect 8850 4519 8906 4528
rect 8864 4282 8892 4519
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8956 3534 8984 5578
rect 9048 5302 9076 5782
rect 9140 5778 9168 6287
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9048 4486 9076 5102
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9140 4185 9168 4966
rect 9126 4176 9182 4185
rect 9126 4111 9182 4120
rect 9232 3942 9260 6734
rect 9324 5710 9352 8434
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9324 3398 9352 4422
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 2990 9352 3334
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8496 2310 8524 2790
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8404 2094 8524 2122
rect 8496 800 8524 2094
rect 9416 800 9444 7822
rect 9678 7440 9734 7449
rect 9678 7375 9734 7384
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9508 3233 9536 3878
rect 9600 3398 9628 6870
rect 9692 3602 9720 7375
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9494 3224 9550 3233
rect 9494 3159 9550 3168
rect 9508 2922 9536 3159
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9692 2650 9720 2858
rect 9784 2650 9812 13670
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 9864 10668 9916 10674
rect 9916 10628 9996 10656
rect 9864 10610 9916 10616
rect 9862 10432 9918 10441
rect 9862 10367 9918 10376
rect 9876 10130 9904 10367
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9876 9994 9904 10066
rect 9968 9994 9996 10628
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 10046 9480 10102 9489
rect 10046 9415 10102 9424
rect 10060 8974 10088 9415
rect 10138 9344 10194 9353
rect 10138 9279 10194 9288
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10152 8906 10180 9279
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9876 8090 9904 8298
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 10060 7818 10088 8366
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 10140 6384 10192 6390
rect 10244 6372 10272 13874
rect 10520 13870 10548 15234
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 12070 14512 12126 14521
rect 12070 14447 12126 14456
rect 10508 13864 10560 13870
rect 10560 13824 10640 13852
rect 10508 13806 10560 13812
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10336 12986 10364 13330
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10428 12594 10456 13194
rect 10520 12832 10548 13262
rect 10612 13258 10640 13824
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10600 12844 10652 12850
rect 10520 12804 10600 12832
rect 10600 12786 10652 12792
rect 10428 12566 10548 12594
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10336 11286 10364 12174
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10324 11280 10376 11286
rect 10324 11222 10376 11228
rect 10336 10810 10364 11222
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10336 10266 10364 10542
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10336 7546 10364 9318
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10428 6866 10456 12038
rect 10520 10606 10548 12566
rect 10612 11778 10640 12786
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10704 11898 10732 12582
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10612 11750 10732 11778
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10612 10674 10640 11290
rect 10704 11218 10732 11750
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10192 6344 10272 6372
rect 10140 6326 10192 6332
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 10244 4570 10272 6344
rect 10336 5778 10364 6734
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10428 6458 10456 6666
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10414 6352 10470 6361
rect 10414 6287 10470 6296
rect 10428 5846 10456 6287
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10428 5409 10456 5646
rect 10414 5400 10470 5409
rect 10414 5335 10470 5344
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10428 4758 10456 5238
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10520 4690 10548 10406
rect 10704 10169 10732 10950
rect 10690 10160 10746 10169
rect 10690 10095 10746 10104
rect 10704 9994 10732 10095
rect 10692 9988 10744 9994
rect 10612 9948 10692 9976
rect 10612 9450 10640 9948
rect 10692 9930 10744 9936
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10704 9450 10732 9658
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10612 7818 10640 9386
rect 10796 9382 10824 13262
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10888 12238 10916 12786
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 11072 12306 11100 12650
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8362 10732 8774
rect 10796 8412 10824 9318
rect 10888 9178 10916 12038
rect 10968 11688 11020 11694
rect 10966 11656 10968 11665
rect 11020 11656 11022 11665
rect 10966 11591 11022 11600
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10980 9489 11008 11018
rect 11072 10282 11100 12242
rect 11164 10810 11192 12582
rect 11256 12442 11284 13330
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11256 11744 11284 12174
rect 11336 11756 11388 11762
rect 11256 11716 11336 11744
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11256 10742 11284 11716
rect 11336 11698 11388 11704
rect 11440 11626 11468 12718
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11072 10254 11192 10282
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9654 11100 9930
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10966 9480 11022 9489
rect 10966 9415 11022 9424
rect 11164 9353 11192 10254
rect 11256 10198 11284 10542
rect 11244 10192 11296 10198
rect 11244 10134 11296 10140
rect 11348 9654 11376 11154
rect 11426 11112 11482 11121
rect 11426 11047 11482 11056
rect 11440 10674 11468 11047
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11440 10266 11468 10406
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11440 10033 11468 10202
rect 11426 10024 11482 10033
rect 11426 9959 11482 9968
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11150 9344 11206 9353
rect 11150 9279 11206 9288
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8634 11100 8910
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11058 8528 11114 8537
rect 11058 8463 11114 8472
rect 10876 8424 10928 8430
rect 10796 8384 10876 8412
rect 10876 8366 10928 8372
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10612 6882 10640 7414
rect 10704 7002 10732 7890
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10612 6854 10732 6882
rect 10598 6352 10654 6361
rect 10598 6287 10654 6296
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10244 4542 10456 4570
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 10324 4208 10376 4214
rect 10322 4176 10324 4185
rect 10376 4176 10378 4185
rect 10232 4140 10284 4146
rect 10322 4111 10378 4120
rect 10232 4082 10284 4088
rect 10244 3942 10272 4082
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10232 3460 10284 3466
rect 10232 3402 10284 3408
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 10244 2650 10272 3402
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10428 2530 10456 4542
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10520 3534 10548 3946
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10152 2502 10456 2530
rect 10152 2446 10180 2502
rect 10140 2440 10192 2446
rect 10612 2428 10640 6287
rect 10704 3584 10732 6854
rect 10796 5914 10824 7822
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10796 4078 10824 4490
rect 10888 4078 10916 8366
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10980 7478 11008 8298
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 11072 7274 11100 8463
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 7410 11192 8230
rect 11256 7546 11284 9454
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11242 7440 11298 7449
rect 11152 7404 11204 7410
rect 11242 7375 11298 7384
rect 11152 7346 11204 7352
rect 11256 7342 11284 7375
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10784 3596 10836 3602
rect 10704 3556 10784 3584
rect 10784 3538 10836 3544
rect 10888 3534 10916 4014
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10704 2446 10732 2994
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10888 2582 10916 2790
rect 10980 2650 11008 7142
rect 11242 7032 11298 7041
rect 11242 6967 11244 6976
rect 11296 6967 11298 6976
rect 11244 6938 11296 6944
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11072 5710 11100 6734
rect 11164 5778 11192 6734
rect 11244 6656 11296 6662
rect 11242 6624 11244 6633
rect 11296 6624 11298 6633
rect 11242 6559 11298 6568
rect 11348 6186 11376 8502
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11256 5914 11284 6054
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11060 5568 11112 5574
rect 11058 5536 11060 5545
rect 11112 5536 11114 5545
rect 11058 5471 11114 5480
rect 11060 4480 11112 4486
rect 11164 4468 11192 5714
rect 11112 4440 11192 4468
rect 11060 4422 11112 4428
rect 11164 3602 11192 4440
rect 11348 4321 11376 6122
rect 11440 4758 11468 9862
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11334 4312 11390 4321
rect 11334 4247 11390 4256
rect 11532 3942 11560 13738
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11624 11234 11652 13126
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11716 11354 11744 12582
rect 12084 12345 12112 14447
rect 13924 14006 13952 16200
rect 15016 15224 15068 15230
rect 14646 15192 14702 15201
rect 15016 15166 15068 15172
rect 14646 15127 14702 15136
rect 13912 14000 13964 14006
rect 12162 13968 12218 13977
rect 13912 13942 13964 13948
rect 12162 13903 12218 13912
rect 12070 12336 12126 12345
rect 11980 12300 12032 12306
rect 12176 12306 12204 13903
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12070 12271 12126 12280
rect 12164 12300 12216 12306
rect 11980 12242 12032 12248
rect 12164 12242 12216 12248
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11794 11792 11850 11801
rect 11794 11727 11850 11736
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11624 11206 11744 11234
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10198 11652 10950
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11610 9888 11666 9897
rect 11610 9823 11666 9832
rect 11624 9722 11652 9823
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11624 9518 11652 9658
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11624 6225 11652 9454
rect 11610 6216 11666 6225
rect 11610 6151 11666 6160
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11624 5098 11652 6054
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11150 3224 11206 3233
rect 11348 3194 11376 3538
rect 11150 3159 11206 3168
rect 11336 3188 11388 3194
rect 11164 2990 11192 3159
rect 11336 3130 11388 3136
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11440 2650 11468 3674
rect 11624 3058 11652 5034
rect 11716 4214 11744 11206
rect 11808 11082 11836 11727
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11794 10568 11850 10577
rect 11794 10503 11796 10512
rect 11848 10503 11850 10512
rect 11796 10474 11848 10480
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11808 9178 11836 9318
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11900 8294 11928 12038
rect 11992 9500 12020 12242
rect 12176 12050 12204 12242
rect 12268 12238 12296 12786
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12176 12022 12296 12050
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12084 10441 12112 11766
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12070 10432 12126 10441
rect 12070 10367 12126 10376
rect 12176 10169 12204 10542
rect 12162 10160 12218 10169
rect 12162 10095 12218 10104
rect 12176 10062 12204 10095
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12072 9512 12124 9518
rect 11992 9472 12072 9500
rect 11992 9058 12020 9472
rect 12164 9512 12216 9518
rect 12072 9454 12124 9460
rect 12162 9480 12164 9489
rect 12216 9480 12218 9489
rect 12162 9415 12218 9424
rect 12268 9217 12296 12022
rect 12452 10418 12480 13398
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12360 10390 12480 10418
rect 12360 9500 12388 10390
rect 12360 9472 12480 9500
rect 12254 9208 12310 9217
rect 12254 9143 12310 9152
rect 12348 9104 12400 9110
rect 12346 9072 12348 9081
rect 12400 9072 12402 9081
rect 11992 9030 12296 9058
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11888 8016 11940 8022
rect 11888 7958 11940 7964
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11808 5370 11836 7142
rect 11900 5896 11928 7958
rect 11992 7857 12020 8910
rect 12176 8634 12204 8910
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12084 7954 12112 8434
rect 12176 8090 12204 8434
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12268 8022 12296 9030
rect 12346 9007 12402 9016
rect 12452 8974 12480 9472
rect 12544 9042 12572 12582
rect 12636 11626 12664 13330
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 13188 11150 13216 11698
rect 13176 11144 13228 11150
rect 12622 11112 12678 11121
rect 13176 11086 13228 11092
rect 12622 11047 12678 11056
rect 12636 9761 12664 11047
rect 13188 10606 13216 11086
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10266 12756 10406
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 12716 10260 12768 10266
rect 13280 10248 13308 12854
rect 13924 12306 13952 13942
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 10810 13400 11494
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 10266 13492 10542
rect 13556 10470 13584 11154
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 12716 10202 12768 10208
rect 12912 10220 13308 10248
rect 13452 10260 13504 10266
rect 12622 9752 12678 9761
rect 12622 9687 12678 9696
rect 12912 9518 12940 10220
rect 13452 10202 13504 10208
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13280 9586 13308 10066
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 12900 9512 12952 9518
rect 12622 9480 12678 9489
rect 13648 9489 13676 11562
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13740 9722 13768 10746
rect 13832 10266 13860 11494
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13818 10024 13874 10033
rect 13818 9959 13874 9968
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 12900 9454 12952 9460
rect 13634 9480 13690 9489
rect 12622 9415 12678 9424
rect 12716 9444 12768 9450
rect 12636 9042 12664 9415
rect 13634 9415 13690 9424
rect 12716 9386 12768 9392
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12360 8634 12388 8774
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11978 7848 12034 7857
rect 11978 7783 12034 7792
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11992 6186 12020 7482
rect 12084 6866 12112 7890
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12162 7032 12218 7041
rect 12162 6967 12218 6976
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12176 6322 12204 6967
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 11900 5868 12020 5896
rect 11886 5808 11942 5817
rect 11886 5743 11942 5752
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11808 4554 11836 4966
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11794 4312 11850 4321
rect 11794 4247 11850 4256
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 11808 4146 11836 4247
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11704 3664 11756 3670
rect 11702 3632 11704 3641
rect 11756 3632 11758 3641
rect 11702 3567 11758 3576
rect 11702 3360 11758 3369
rect 11702 3295 11758 3304
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 10140 2382 10192 2388
rect 10336 2400 10640 2428
rect 10692 2440 10744 2446
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 10336 800 10364 2400
rect 10692 2382 10744 2388
rect 11532 1306 11560 2926
rect 11716 2514 11744 3295
rect 11808 3126 11836 4082
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11900 2854 11928 5743
rect 11992 3194 12020 5868
rect 12084 3738 12112 6054
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12176 5302 12204 5714
rect 12164 5296 12216 5302
rect 12164 5238 12216 5244
rect 12268 4978 12296 7414
rect 12360 5409 12388 8026
rect 12346 5400 12402 5409
rect 12346 5335 12402 5344
rect 12268 4950 12388 4978
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12176 4729 12204 4762
rect 12162 4720 12218 4729
rect 12162 4655 12218 4664
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11256 1278 11560 1306
rect 11256 800 11284 1278
rect 12176 800 12204 4558
rect 12254 4176 12310 4185
rect 12254 4111 12310 4120
rect 12268 4010 12296 4111
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 12254 3904 12310 3913
rect 12254 3839 12310 3848
rect 12268 2650 12296 3839
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12360 2446 12388 4950
rect 12452 4690 12480 8230
rect 12544 7698 12572 8978
rect 12636 8294 12664 8978
rect 12728 8514 12756 9386
rect 13176 9376 13228 9382
rect 13544 9376 13596 9382
rect 13266 9344 13322 9353
rect 13228 9324 13266 9330
rect 13176 9318 13266 9324
rect 13188 9302 13266 9318
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13188 8537 13216 9302
rect 13544 9318 13596 9324
rect 13266 9279 13322 9288
rect 13556 9217 13584 9318
rect 13542 9208 13598 9217
rect 13542 9143 13598 9152
rect 13268 9104 13320 9110
rect 13320 9052 13400 9058
rect 13268 9046 13400 9052
rect 13280 9030 13400 9046
rect 13740 9042 13768 9522
rect 13174 8528 13230 8537
rect 12728 8498 12940 8514
rect 12728 8492 12952 8498
rect 12728 8486 12900 8492
rect 13174 8463 13230 8472
rect 13268 8492 13320 8498
rect 12900 8434 12952 8440
rect 13268 8434 13320 8440
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 8090 12664 8230
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12544 7670 12664 7698
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12544 5846 12572 7346
rect 12636 5914 12664 7670
rect 12728 7546 12756 8366
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 13280 7954 13308 8434
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13372 7750 13400 9030
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13464 7546 13492 8434
rect 13740 8090 13768 8978
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13726 7848 13782 7857
rect 13832 7834 13860 9959
rect 13924 8566 13952 11834
rect 14094 11656 14150 11665
rect 14094 11591 14150 11600
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 14016 9926 14044 11222
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 14108 9654 14136 11591
rect 14200 11286 14228 12106
rect 14292 11937 14320 12718
rect 14278 11928 14334 11937
rect 14278 11863 14334 11872
rect 14188 11280 14240 11286
rect 14188 11222 14240 11228
rect 14200 10606 14228 11222
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14292 10266 14320 11863
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14476 10305 14504 11766
rect 14462 10296 14518 10305
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14372 10260 14424 10266
rect 14462 10231 14518 10240
rect 14372 10202 14424 10208
rect 14280 10056 14332 10062
rect 14384 10044 14412 10202
rect 14332 10016 14412 10044
rect 14280 9998 14332 10004
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14200 9586 14228 9862
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14094 9208 14150 9217
rect 14094 9143 14150 9152
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13832 7806 14044 7834
rect 13726 7783 13782 7792
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13464 7410 13492 7482
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12728 6390 12756 7210
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 13464 7002 13492 7346
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13740 6934 13768 7783
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13832 7002 13860 7346
rect 14016 7290 14044 7806
rect 13924 7262 14044 7290
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13728 6928 13780 6934
rect 13556 6888 13728 6916
rect 13268 6860 13320 6866
rect 13320 6820 13400 6848
rect 13268 6802 13320 6808
rect 13084 6792 13136 6798
rect 12990 6760 13046 6769
rect 13084 6734 13136 6740
rect 12990 6695 12992 6704
rect 13044 6695 13046 6704
rect 12992 6666 13044 6672
rect 12716 6384 12768 6390
rect 13096 6361 13124 6734
rect 12716 6326 12768 6332
rect 13082 6352 13138 6361
rect 13082 6287 13138 6296
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12544 5642 12572 5782
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12898 5400 12954 5409
rect 12898 5335 12954 5344
rect 12912 5234 12940 5335
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 13188 5030 13216 5850
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12544 3738 12572 3946
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12728 3534 12756 4422
rect 12820 4282 12848 4558
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 13188 3670 13216 4082
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 12912 2990 12940 3334
rect 12440 2984 12492 2990
rect 12900 2984 12952 2990
rect 12492 2932 12756 2938
rect 12440 2926 12756 2932
rect 12900 2926 12952 2932
rect 12452 2910 12756 2926
rect 12728 2854 12756 2910
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13096 2106 13124 2382
rect 13084 2100 13136 2106
rect 13084 2042 13136 2048
rect 13188 1850 13216 3334
rect 13280 2446 13308 5102
rect 13372 2961 13400 6820
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13464 5370 13492 6054
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13464 4826 13492 5102
rect 13556 5098 13584 6888
rect 13728 6870 13780 6876
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13358 2952 13414 2961
rect 13358 2887 13414 2896
rect 13464 2514 13492 4490
rect 13556 3602 13584 4694
rect 13648 3942 13676 6122
rect 13740 5302 13768 6258
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13740 4826 13768 5238
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13726 4040 13782 4049
rect 13832 4026 13860 6122
rect 13924 6118 13952 7262
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 6458 14044 7142
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14108 6202 14136 9143
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14200 7002 14228 8502
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14016 6174 14136 6202
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13782 3998 13860 4026
rect 13726 3975 13782 3984
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13634 3496 13690 3505
rect 13634 3431 13690 3440
rect 13648 2650 13676 3431
rect 13740 2650 13768 3975
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13832 2582 13860 2790
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13096 1822 13216 1850
rect 13096 800 13124 1822
rect 13924 800 13952 5646
rect 14016 4214 14044 6174
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14108 4758 14136 6054
rect 14200 5642 14228 6938
rect 14292 6225 14320 9998
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 9178 14412 9318
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14384 7954 14412 8366
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14476 7528 14504 10231
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14568 9586 14596 10066
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14568 9178 14596 9522
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14384 7500 14504 7528
rect 14384 7002 14412 7500
rect 14568 7274 14596 7686
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14476 6798 14504 7210
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14384 6458 14412 6666
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14278 6216 14334 6225
rect 14278 6151 14334 6160
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14096 4752 14148 4758
rect 14096 4694 14148 4700
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 14016 3534 14044 4150
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 14016 2310 14044 2790
rect 14108 2446 14136 3402
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 14200 2106 14228 5306
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14292 4690 14320 5170
rect 14384 5166 14412 6394
rect 14476 6322 14504 6734
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14476 5914 14504 6258
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14568 5370 14596 6054
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14292 4146 14320 4626
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14292 3738 14320 4082
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14384 2854 14412 4694
rect 14568 4078 14596 4966
rect 14660 4729 14688 15127
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14752 11014 14780 11698
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10606 14780 10950
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14752 9926 14780 10542
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14738 9752 14794 9761
rect 14738 9687 14794 9696
rect 14752 6118 14780 9687
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14738 5808 14794 5817
rect 14738 5743 14794 5752
rect 14752 5710 14780 5743
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14844 5545 14872 9454
rect 14936 9178 14964 12854
rect 15028 11694 15056 15166
rect 15106 14512 15162 14521
rect 15106 14447 15162 14456
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15014 10432 15070 10441
rect 15014 10367 15070 10376
rect 15028 9722 15056 10367
rect 15120 10266 15148 14447
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15212 12481 15240 12582
rect 15198 12472 15254 12481
rect 15198 12407 15254 12416
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15212 11529 15240 11834
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15198 11520 15254 11529
rect 15198 11455 15254 11464
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 15120 9586 15148 9862
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 15120 9042 15148 9522
rect 15212 9489 15240 10406
rect 15304 10266 15332 11562
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15304 9761 15332 10066
rect 15290 9752 15346 9761
rect 15290 9687 15346 9696
rect 15198 9480 15254 9489
rect 15198 9415 15254 9424
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15120 8906 15148 8978
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14936 6118 14964 8298
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 15028 5778 15056 8774
rect 15120 8362 15148 8842
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 15120 7886 15148 8298
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15120 7342 15148 7822
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15212 7449 15240 7686
rect 15396 7562 15424 12174
rect 15488 10577 15516 16487
rect 17866 16200 17922 17000
rect 17774 16144 17830 16153
rect 17774 16079 17830 16088
rect 15658 15872 15714 15881
rect 15658 15807 15714 15816
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15580 12306 15608 13466
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15580 11830 15608 12106
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15474 10568 15530 10577
rect 15474 10503 15530 10512
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15304 7534 15424 7562
rect 15198 7440 15254 7449
rect 15198 7375 15254 7384
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15120 6254 15148 6734
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15120 5846 15148 6190
rect 15212 6118 15240 7278
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 14830 5536 14886 5545
rect 14830 5471 14886 5480
rect 14646 4720 14702 4729
rect 14646 4655 14702 4664
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14660 3942 14688 4655
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14752 3097 14780 3878
rect 14844 3738 14872 5471
rect 14936 4010 14964 5578
rect 15120 5234 15148 5782
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14936 3466 14964 3946
rect 14924 3460 14976 3466
rect 14924 3402 14976 3408
rect 14738 3088 14794 3097
rect 14738 3023 14740 3032
rect 14792 3023 14794 3032
rect 14740 2994 14792 3000
rect 14752 2963 14780 2994
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 15028 2394 15056 4490
rect 15120 4486 15148 5170
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15120 4146 15148 4422
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 14844 2366 15056 2394
rect 14188 2100 14240 2106
rect 14188 2042 14240 2048
rect 14844 800 14872 2366
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 15212 1193 15240 1294
rect 15198 1184 15254 1193
rect 15198 1119 15254 1128
rect 3422 504 3478 513
rect 3422 439 3478 448
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15304 241 15332 7534
rect 15488 6610 15516 10406
rect 15580 10198 15608 11154
rect 15672 10248 15700 15807
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 15782 14172 16078 14192
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 13297 16252 13670
rect 16210 13288 16266 13297
rect 16210 13223 16266 13232
rect 16210 13152 16266 13161
rect 15782 13084 16078 13104
rect 16210 13087 16266 13096
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15750 12880 15806 12889
rect 15750 12815 15806 12824
rect 15764 12714 15792 12815
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 16224 11257 16252 13087
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16210 11248 16266 11257
rect 16210 11183 16266 11192
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15856 10470 15884 10542
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15672 10220 15792 10248
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15764 10130 15792 10220
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15580 8945 15608 9998
rect 15566 8936 15622 8945
rect 15566 8871 15622 8880
rect 15672 8430 15700 10066
rect 16040 9994 16068 10406
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15856 8974 15884 9454
rect 16316 9178 16344 12038
rect 16408 10169 16436 14010
rect 16960 13394 16988 14486
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 16592 11082 16620 11562
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16684 10810 16712 12242
rect 16960 12220 16988 12786
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17052 12442 17080 12582
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17040 12232 17092 12238
rect 16960 12192 17040 12220
rect 17040 12174 17092 12180
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16764 11620 16816 11626
rect 16764 11562 16816 11568
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16394 10160 16450 10169
rect 16394 10095 16450 10104
rect 16500 10044 16528 10542
rect 16580 10464 16632 10470
rect 16578 10432 16580 10441
rect 16672 10464 16724 10470
rect 16632 10432 16634 10441
rect 16672 10406 16724 10412
rect 16578 10367 16634 10376
rect 16408 10016 16528 10044
rect 16408 9466 16436 10016
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9722 16528 9862
rect 16578 9752 16634 9761
rect 16488 9716 16540 9722
rect 16578 9687 16634 9696
rect 16488 9658 16540 9664
rect 16408 9438 16528 9466
rect 16396 9376 16448 9382
rect 16500 9353 16528 9438
rect 16396 9318 16448 9324
rect 16486 9344 16542 9353
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 16408 8809 16436 9318
rect 16486 9279 16542 9288
rect 16394 8800 16450 8809
rect 15782 8732 16078 8752
rect 16394 8735 16450 8744
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 16500 8430 16528 9279
rect 16592 8537 16620 9687
rect 16684 9625 16712 10406
rect 16670 9616 16726 9625
rect 16670 9551 16726 9560
rect 16684 9178 16712 9551
rect 16776 9518 16804 11562
rect 16868 10674 16896 11630
rect 17052 11558 17080 12174
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16946 10840 17002 10849
rect 16946 10775 17002 10784
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16854 10568 16910 10577
rect 16854 10503 16910 10512
rect 16868 9897 16896 10503
rect 16960 10198 16988 10775
rect 17052 10538 17080 11494
rect 17144 11354 17172 12582
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17040 10532 17092 10538
rect 17040 10474 17092 10480
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16960 10033 16988 10134
rect 16946 10024 17002 10033
rect 16946 9959 17002 9968
rect 16854 9888 16910 9897
rect 16854 9823 16910 9832
rect 16854 9752 16910 9761
rect 16854 9687 16910 9696
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16578 8528 16634 8537
rect 16578 8463 16634 8472
rect 15660 8424 15712 8430
rect 16488 8424 16540 8430
rect 15660 8366 15712 8372
rect 16118 8392 16174 8401
rect 16488 8366 16540 8372
rect 16776 8362 16804 8774
rect 16118 8327 16174 8336
rect 16764 8356 16816 8362
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15580 7585 15608 7686
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15566 7576 15622 7585
rect 15782 7568 16078 7588
rect 15566 7511 15622 7520
rect 16132 7342 16160 8327
rect 16764 8298 16816 8304
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16224 8090 16252 8230
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16316 7954 16344 8230
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15396 6582 15516 6610
rect 15396 6458 15424 6582
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15396 5681 15424 6054
rect 15488 5778 15516 6122
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15382 5672 15438 5681
rect 15382 5607 15438 5616
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15396 4826 15424 5510
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15488 3058 15516 4014
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15488 2514 15516 2994
rect 15580 2582 15608 7142
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15672 5166 15700 6054
rect 16132 5914 16160 7142
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15672 3534 15700 5102
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15856 4622 15884 4762
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 16118 3088 16174 3097
rect 16118 3023 16174 3032
rect 16132 2990 16160 3023
rect 15752 2984 15804 2990
rect 15752 2926 15804 2932
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15672 2650 15700 2858
rect 15764 2650 15792 2926
rect 16118 2680 16174 2689
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15752 2644 15804 2650
rect 16118 2615 16174 2624
rect 15752 2586 15804 2592
rect 16132 2582 16160 2615
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16224 1986 16252 7278
rect 16316 5710 16344 7890
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16316 3058 16344 3470
rect 16408 3194 16436 7414
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16500 5302 16528 7142
rect 16592 6866 16620 7686
rect 16684 7342 16712 8230
rect 16776 7818 16804 8298
rect 16764 7812 16816 7818
rect 16764 7754 16816 7760
rect 16776 7410 16804 7754
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16580 6860 16632 6866
rect 16632 6820 16712 6848
rect 16580 6802 16632 6808
rect 16580 5568 16632 5574
rect 16578 5536 16580 5545
rect 16632 5536 16634 5545
rect 16578 5471 16634 5480
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16500 4078 16528 4966
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16316 2446 16344 2994
rect 16592 2990 16620 5102
rect 16684 4690 16712 6820
rect 16868 6746 16896 9687
rect 17236 9466 17264 13262
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17328 9994 17356 12242
rect 17512 11762 17540 12242
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17406 11520 17462 11529
rect 17406 11455 17462 11464
rect 17420 10674 17448 11455
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17512 10441 17540 10542
rect 17498 10432 17554 10441
rect 17498 10367 17554 10376
rect 17406 10296 17462 10305
rect 17406 10231 17462 10240
rect 17420 10130 17448 10231
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17052 9438 17264 9466
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16776 6730 16896 6746
rect 16764 6724 16896 6730
rect 16816 6718 16896 6724
rect 16764 6666 16816 6672
rect 16776 5166 16804 6666
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16868 6186 16896 6598
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16776 4758 16804 4966
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16868 4554 16896 6122
rect 16960 5846 16988 7686
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16960 5166 16988 5510
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 15764 1958 16252 1986
rect 15764 800 15792 1958
rect 16684 800 16712 3606
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16776 2650 16804 2790
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 16868 2582 16896 3334
rect 16960 2922 16988 3878
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 17052 1465 17080 9438
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17130 9208 17186 9217
rect 17130 9143 17186 9152
rect 17144 8430 17172 9143
rect 17236 9042 17264 9318
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 17236 8498 17264 8978
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17236 7834 17264 8298
rect 17328 7954 17356 9454
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17236 7806 17356 7834
rect 17130 6896 17186 6905
rect 17130 6831 17132 6840
rect 17184 6831 17186 6840
rect 17132 6802 17184 6808
rect 17224 6792 17276 6798
rect 17222 6760 17224 6769
rect 17276 6760 17278 6769
rect 17222 6695 17278 6704
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 5234 17264 6598
rect 17328 6186 17356 7806
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17420 5846 17448 10066
rect 17500 9444 17552 9450
rect 17500 9386 17552 9392
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17328 5234 17356 5646
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17420 4740 17448 5782
rect 17328 4712 17448 4740
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17144 3058 17172 4422
rect 17328 4078 17356 4712
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17420 4146 17448 4490
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17420 3466 17448 4082
rect 17408 3460 17460 3466
rect 17408 3402 17460 3408
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17038 1456 17094 1465
rect 17038 1391 17094 1400
rect 15290 232 15346 241
rect 15290 167 15346 176
rect 15750 0 15806 800
rect 16670 0 16726 800
rect 17512 785 17540 9386
rect 17604 800 17632 13942
rect 17682 13560 17738 13569
rect 17682 13495 17738 13504
rect 17696 12170 17724 13495
rect 17788 12986 17816 16079
rect 17880 13938 17908 16200
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17788 12442 17816 12922
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17696 11150 17724 12106
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17696 8362 17724 11086
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17788 8129 17816 11494
rect 17880 11150 17908 12174
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17958 11112 18014 11121
rect 17880 10674 17908 11086
rect 17958 11047 18014 11056
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17880 10062 17908 10610
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17774 8120 17830 8129
rect 17774 8055 17830 8064
rect 17684 7812 17736 7818
rect 17684 7754 17736 7760
rect 17696 6798 17724 7754
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17696 5710 17724 6734
rect 17788 6225 17816 7686
rect 17880 7313 17908 9318
rect 17972 8090 18000 11047
rect 18248 9217 18276 12582
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18234 9208 18290 9217
rect 18234 9143 18290 9152
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18064 7426 18092 8978
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 17972 7398 18092 7426
rect 17866 7304 17922 7313
rect 17866 7239 17922 7248
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17774 6216 17830 6225
rect 17774 6151 17830 6160
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17788 3738 17816 6054
rect 17880 5817 17908 7142
rect 17866 5808 17922 5817
rect 17866 5743 17922 5752
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17972 5522 18000 7398
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 6934 18092 7278
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18156 5914 18184 6734
rect 18248 6497 18276 8502
rect 18340 6905 18368 8774
rect 18432 7857 18460 10406
rect 18418 7848 18474 7857
rect 18418 7783 18474 7792
rect 18326 6896 18382 6905
rect 18326 6831 18382 6840
rect 18234 6488 18290 6497
rect 18234 6423 18290 6432
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 17880 4865 17908 5510
rect 17972 5494 18092 5522
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17866 4856 17922 4865
rect 17972 4826 18000 5306
rect 17866 4791 17922 4800
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17972 4078 18000 4762
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 18064 3738 18092 5494
rect 18248 5137 18276 6054
rect 18234 5128 18290 5137
rect 18234 5063 18290 5072
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4457 18276 4966
rect 18234 4448 18290 4457
rect 18234 4383 18290 4392
rect 18234 4176 18290 4185
rect 18234 4111 18290 4120
rect 18248 3942 18276 4111
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18234 3768 18290 3777
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 18052 3732 18104 3738
rect 18234 3703 18236 3712
rect 18052 3674 18104 3680
rect 18288 3703 18290 3712
rect 18236 3674 18288 3680
rect 18524 800 18552 13262
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 18602 9072 18658 9081
rect 18602 9007 18658 9016
rect 17498 776 17554 785
rect 17498 711 17554 720
rect 17590 0 17646 800
rect 18510 0 18566 800
rect 18616 513 18644 9007
rect 19444 800 19472 11834
rect 18602 504 18658 513
rect 18602 439 18658 448
rect 19430 0 19486 800
<< via2 >>
rect 1582 16496 1638 16552
rect 1490 15136 1546 15192
rect 4066 16768 4122 16824
rect 1674 14864 1730 14920
rect 1766 14184 1822 14240
rect 2870 16088 2926 16144
rect 2778 14456 2834 14512
rect 3974 15816 4030 15872
rect 2962 15408 3018 15464
rect 15474 16496 15530 16552
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 1766 13776 1822 13832
rect 2778 13504 2834 13560
rect 1674 9016 1730 9072
rect 1766 7928 1822 7984
rect 1950 6704 2006 6760
rect 1582 5344 1638 5400
rect 1122 4392 1178 4448
rect 1490 4800 1546 4856
rect 1858 4120 1914 4176
rect 1490 3984 1546 4040
rect 1490 3712 1546 3768
rect 1858 2896 1914 2952
rect 2778 13252 2834 13288
rect 2778 13232 2780 13252
rect 2780 13232 2832 13252
rect 2832 13232 2834 13252
rect 3238 12824 3294 12880
rect 2594 12280 2650 12336
rect 2778 9968 2834 10024
rect 2686 9152 2742 9208
rect 3054 10124 3110 10160
rect 3054 10104 3056 10124
rect 3056 10104 3108 10124
rect 3108 10104 3110 10124
rect 3054 8880 3110 8936
rect 2686 6704 2742 6760
rect 2594 6432 2650 6488
rect 2870 6704 2926 6760
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3790 12552 3846 12608
rect 3698 12280 3754 12336
rect 3606 11872 3662 11928
rect 3514 8880 3570 8936
rect 3146 6024 3202 6080
rect 2778 5616 2834 5672
rect 2226 3576 2282 3632
rect 2686 2624 2742 2680
rect 3054 4564 3056 4584
rect 3056 4564 3108 4584
rect 3108 4564 3110 4584
rect 3054 4528 3110 4564
rect 2870 3440 2926 3496
rect 4066 12144 4122 12200
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 4802 11736 4858 11792
rect 4066 11192 4122 11248
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 4066 10240 4122 10296
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 4066 9424 4122 9480
rect 4618 10648 4674 10704
rect 4250 9152 4306 9208
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 4250 7928 4306 7984
rect 5078 11192 5134 11248
rect 4894 11056 4950 11112
rect 4526 8744 4582 8800
rect 3422 6296 3478 6352
rect 3330 6160 3386 6216
rect 3238 3984 3294 4040
rect 3238 2760 3294 2816
rect 3238 1844 3240 1864
rect 3240 1844 3292 1864
rect 3292 1844 3294 1864
rect 3238 1808 3294 1844
rect 3146 1128 3202 1184
rect 2870 720 2926 776
rect 2778 176 2834 232
rect 3698 7248 3754 7304
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 3790 6840 3846 6896
rect 4066 6860 4122 6896
rect 4066 6840 4068 6860
rect 4068 6840 4120 6860
rect 4120 6840 4122 6860
rect 3514 3168 3570 3224
rect 3514 3032 3570 3088
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 4434 5752 4490 5808
rect 4250 5072 4306 5128
rect 3974 4700 3976 4720
rect 3976 4700 4028 4720
rect 4028 4700 4030 4720
rect 3974 4664 4030 4700
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 3698 2080 3754 2136
rect 4066 3032 4122 3088
rect 3882 2352 3938 2408
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 4434 4820 4490 4856
rect 4434 4800 4436 4820
rect 4436 4800 4488 4820
rect 4488 4800 4490 4820
rect 5262 10804 5318 10840
rect 5262 10784 5264 10804
rect 5264 10784 5316 10804
rect 5316 10784 5318 10804
rect 4894 6976 4950 7032
rect 5354 9832 5410 9888
rect 5354 8744 5410 8800
rect 5262 8236 5264 8256
rect 5264 8236 5316 8256
rect 5316 8236 5318 8256
rect 4802 5752 4858 5808
rect 4618 5072 4674 5128
rect 5262 8200 5318 8236
rect 5446 7792 5502 7848
rect 5262 5072 5318 5128
rect 5998 11600 6054 11656
rect 5722 10648 5778 10704
rect 5722 10376 5778 10432
rect 5998 10648 6054 10704
rect 5906 9424 5962 9480
rect 5814 8336 5870 8392
rect 4526 3848 4582 3904
rect 4710 3884 4712 3904
rect 4712 3884 4764 3904
rect 4764 3884 4766 3904
rect 4710 3848 4766 3884
rect 5078 3712 5134 3768
rect 4986 3576 5042 3632
rect 4434 3168 4490 3224
rect 4066 1400 4122 1456
rect 5538 3984 5594 4040
rect 5722 3304 5778 3360
rect 5998 3848 6054 3904
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6274 12008 6330 12064
rect 7378 12008 7434 12064
rect 6458 10512 6514 10568
rect 6458 9968 6514 10024
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 7286 11056 7342 11112
rect 7102 10784 7158 10840
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 6550 9696 6606 9752
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 7378 9560 7434 9616
rect 7378 9288 7434 9344
rect 6366 8472 6422 8528
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6458 5752 6514 5808
rect 6090 3576 6146 3632
rect 6458 3732 6514 3768
rect 6458 3712 6460 3732
rect 6460 3712 6512 3732
rect 6512 3712 6514 3732
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6734 6840 6790 6896
rect 6642 5616 6698 5672
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 7286 5344 7342 5400
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 7838 12416 7894 12472
rect 7654 10376 7710 10432
rect 7838 9696 7894 9752
rect 7562 6840 7618 6896
rect 7562 5344 7618 5400
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 6458 2624 6514 2680
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 8022 11756 8078 11792
rect 8022 11736 8024 11756
rect 8024 11736 8076 11756
rect 8076 11736 8078 11756
rect 8206 12008 8262 12064
rect 8206 9696 8262 9752
rect 8666 11872 8722 11928
rect 8666 10784 8722 10840
rect 8574 10376 8630 10432
rect 8482 9424 8538 9480
rect 8574 8608 8630 8664
rect 8574 8508 8576 8528
rect 8576 8508 8628 8528
rect 8628 8508 8630 8528
rect 8574 8472 8630 8508
rect 7930 4528 7986 4584
rect 7930 3304 7986 3360
rect 8482 6060 8484 6080
rect 8484 6060 8536 6080
rect 8536 6060 8538 6080
rect 8482 6024 8538 6060
rect 8850 12416 8906 12472
rect 8942 8744 8998 8800
rect 9034 8372 9036 8392
rect 9036 8372 9088 8392
rect 9088 8372 9090 8392
rect 9034 8336 9090 8372
rect 8942 6704 8998 6760
rect 9586 11736 9642 11792
rect 9494 9832 9550 9888
rect 9586 9324 9588 9344
rect 9588 9324 9640 9344
rect 9640 9324 9642 9344
rect 9586 9288 9642 9324
rect 9126 6296 9182 6352
rect 8850 4528 8906 4584
rect 9126 4120 9182 4176
rect 9678 7384 9734 7440
rect 9494 3168 9550 3224
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9862 10376 9918 10432
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 10046 9424 10102 9480
rect 10138 9288 10194 9344
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 12070 14456 12126 14512
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 10414 6296 10470 6352
rect 10414 5344 10470 5400
rect 10690 10104 10746 10160
rect 10966 11636 10968 11656
rect 10968 11636 11020 11656
rect 11020 11636 11022 11656
rect 10966 11600 11022 11636
rect 10966 9424 11022 9480
rect 11426 11056 11482 11112
rect 11426 9968 11482 10024
rect 11150 9288 11206 9344
rect 11058 8472 11114 8528
rect 10598 6296 10654 6352
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10322 4156 10324 4176
rect 10324 4156 10376 4176
rect 10376 4156 10378 4176
rect 10322 4120 10378 4156
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 11242 7384 11298 7440
rect 11242 6996 11298 7032
rect 11242 6976 11244 6996
rect 11244 6976 11296 6996
rect 11296 6976 11298 6996
rect 11242 6604 11244 6624
rect 11244 6604 11296 6624
rect 11296 6604 11298 6624
rect 11242 6568 11298 6604
rect 11058 5516 11060 5536
rect 11060 5516 11112 5536
rect 11112 5516 11114 5536
rect 11058 5480 11114 5516
rect 11334 4256 11390 4312
rect 14646 15136 14702 15192
rect 12162 13912 12218 13968
rect 12070 12280 12126 12336
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 11794 11736 11850 11792
rect 11610 9832 11666 9888
rect 11610 6160 11666 6216
rect 11150 3168 11206 3224
rect 11794 10532 11850 10568
rect 11794 10512 11796 10532
rect 11796 10512 11848 10532
rect 11848 10512 11850 10532
rect 12070 10376 12126 10432
rect 12162 10104 12218 10160
rect 12162 9460 12164 9480
rect 12164 9460 12216 9480
rect 12216 9460 12218 9480
rect 12162 9424 12218 9460
rect 12254 9152 12310 9208
rect 12346 9052 12348 9072
rect 12348 9052 12400 9072
rect 12400 9052 12402 9072
rect 12346 9016 12402 9052
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12622 11056 12678 11112
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12622 9696 12678 9752
rect 12622 9424 12678 9480
rect 13818 9968 13874 10024
rect 13634 9424 13690 9480
rect 11978 7792 12034 7848
rect 12162 6976 12218 7032
rect 11886 5752 11942 5808
rect 11794 4256 11850 4312
rect 11702 3612 11704 3632
rect 11704 3612 11756 3632
rect 11756 3612 11758 3632
rect 11702 3576 11758 3612
rect 11702 3304 11758 3360
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 12346 5344 12402 5400
rect 12162 4664 12218 4720
rect 12254 4120 12310 4176
rect 12254 3848 12310 3904
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 13266 9288 13322 9344
rect 13542 9152 13598 9208
rect 13174 8472 13230 8528
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 13726 7792 13782 7848
rect 14094 11600 14150 11656
rect 14278 11872 14334 11928
rect 14462 10240 14518 10296
rect 14094 9152 14150 9208
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 12990 6724 13046 6760
rect 12990 6704 12992 6724
rect 12992 6704 13044 6724
rect 13044 6704 13046 6724
rect 13082 6296 13138 6352
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12898 5344 12954 5400
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 13358 2896 13414 2952
rect 13726 3984 13782 4040
rect 13634 3440 13690 3496
rect 14278 6160 14334 6216
rect 14738 9696 14794 9752
rect 14738 5752 14794 5808
rect 15106 14456 15162 14512
rect 15014 10376 15070 10432
rect 15198 12416 15254 12472
rect 15198 11464 15254 11520
rect 15290 9696 15346 9752
rect 15198 9424 15254 9480
rect 17774 16088 17830 16144
rect 15658 15816 15714 15872
rect 15474 10512 15530 10568
rect 15198 7384 15254 7440
rect 14830 5480 14886 5536
rect 14646 4664 14702 4720
rect 14738 3052 14794 3088
rect 14738 3032 14740 3052
rect 14740 3032 14792 3052
rect 14792 3032 14794 3052
rect 15198 1128 15254 1184
rect 3422 448 3478 504
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 16210 13232 16266 13288
rect 16210 13096 16266 13152
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15750 12824 15806 12880
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 16210 11192 16266 11248
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15566 8880 15622 8936
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 16394 10104 16450 10160
rect 16578 10412 16580 10432
rect 16580 10412 16632 10432
rect 16632 10412 16634 10432
rect 16578 10376 16634 10412
rect 16578 9696 16634 9752
rect 16486 9288 16542 9344
rect 16394 8744 16450 8800
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 16670 9560 16726 9616
rect 16946 10784 17002 10840
rect 16854 10512 16910 10568
rect 16946 9968 17002 10024
rect 16854 9832 16910 9888
rect 16854 9696 16910 9752
rect 16578 8472 16634 8528
rect 16118 8336 16174 8392
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 15566 7520 15622 7576
rect 15382 5616 15438 5672
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 16118 3032 16174 3088
rect 16118 2624 16174 2680
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 16578 5516 16580 5536
rect 16580 5516 16632 5536
rect 16632 5516 16634 5536
rect 16578 5480 16634 5516
rect 17406 11464 17462 11520
rect 17498 10376 17554 10432
rect 17406 10240 17462 10296
rect 17130 9152 17186 9208
rect 17130 6860 17186 6896
rect 17130 6840 17132 6860
rect 17132 6840 17184 6860
rect 17184 6840 17186 6860
rect 17222 6740 17224 6760
rect 17224 6740 17276 6760
rect 17276 6740 17278 6760
rect 17222 6704 17278 6740
rect 17038 1400 17094 1456
rect 15290 176 15346 232
rect 17682 13504 17738 13560
rect 17958 11056 18014 11112
rect 17774 8064 17830 8120
rect 18234 9152 18290 9208
rect 17866 7248 17922 7304
rect 17774 6160 17830 6216
rect 17866 5752 17922 5808
rect 18418 7792 18474 7848
rect 18326 6840 18382 6896
rect 18234 6432 18290 6488
rect 17866 4800 17922 4856
rect 18234 5072 18290 5128
rect 18234 4392 18290 4448
rect 18234 4120 18290 4176
rect 18234 3732 18290 3768
rect 18234 3712 18236 3732
rect 18236 3712 18288 3732
rect 18288 3712 18290 3732
rect 18602 9016 18658 9072
rect 17498 720 17554 776
rect 18602 448 18658 504
<< metal3 >>
rect 0 16826 800 16856
rect 4061 16826 4127 16829
rect 0 16824 4127 16826
rect 0 16768 4066 16824
rect 4122 16768 4127 16824
rect 0 16766 4127 16768
rect 0 16736 800 16766
rect 4061 16763 4127 16766
rect 15510 16764 15516 16828
rect 15580 16826 15586 16828
rect 19200 16826 20000 16856
rect 15580 16766 20000 16826
rect 15580 16764 15586 16766
rect 19200 16736 20000 16766
rect 0 16554 800 16584
rect 1577 16554 1643 16557
rect 0 16552 1643 16554
rect 0 16496 1582 16552
rect 1638 16496 1643 16552
rect 0 16494 1643 16496
rect 0 16464 800 16494
rect 1577 16491 1643 16494
rect 15469 16554 15535 16557
rect 19200 16554 20000 16584
rect 15469 16552 20000 16554
rect 15469 16496 15474 16552
rect 15530 16496 20000 16552
rect 15469 16494 20000 16496
rect 15469 16491 15535 16494
rect 19200 16464 20000 16494
rect 0 16146 800 16176
rect 2865 16146 2931 16149
rect 0 16144 2931 16146
rect 0 16088 2870 16144
rect 2926 16088 2931 16144
rect 0 16086 2931 16088
rect 0 16056 800 16086
rect 2865 16083 2931 16086
rect 17769 16146 17835 16149
rect 19200 16146 20000 16176
rect 17769 16144 20000 16146
rect 17769 16088 17774 16144
rect 17830 16088 20000 16144
rect 17769 16086 20000 16088
rect 17769 16083 17835 16086
rect 19200 16056 20000 16086
rect 0 15874 800 15904
rect 3969 15874 4035 15877
rect 0 15872 4035 15874
rect 0 15816 3974 15872
rect 4030 15816 4035 15872
rect 0 15814 4035 15816
rect 0 15784 800 15814
rect 3969 15811 4035 15814
rect 15653 15874 15719 15877
rect 19200 15874 20000 15904
rect 15653 15872 20000 15874
rect 15653 15816 15658 15872
rect 15714 15816 20000 15872
rect 15653 15814 20000 15816
rect 15653 15811 15719 15814
rect 19200 15784 20000 15814
rect 0 15466 800 15496
rect 2957 15466 3023 15469
rect 0 15464 3023 15466
rect 0 15408 2962 15464
rect 3018 15408 3023 15464
rect 0 15406 3023 15408
rect 0 15376 800 15406
rect 2957 15403 3023 15406
rect 17166 15404 17172 15468
rect 17236 15466 17242 15468
rect 19200 15466 20000 15496
rect 17236 15406 20000 15466
rect 17236 15404 17242 15406
rect 19200 15376 20000 15406
rect 0 15194 800 15224
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 14641 15194 14707 15197
rect 19200 15194 20000 15224
rect 14641 15192 20000 15194
rect 14641 15136 14646 15192
rect 14702 15136 20000 15192
rect 14641 15134 20000 15136
rect 14641 15131 14707 15134
rect 19200 15104 20000 15134
rect 0 14922 800 14952
rect 1669 14922 1735 14925
rect 0 14920 1735 14922
rect 0 14864 1674 14920
rect 1730 14864 1735 14920
rect 0 14862 1735 14864
rect 0 14832 800 14862
rect 1669 14859 1735 14862
rect 19200 14786 20000 14816
rect 14230 14726 20000 14786
rect 6874 14720 7194 14721
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 14655 13125 14656
rect 0 14514 800 14544
rect 2773 14514 2839 14517
rect 0 14512 2839 14514
rect 0 14456 2778 14512
rect 2834 14456 2839 14512
rect 0 14454 2839 14456
rect 0 14424 800 14454
rect 2773 14451 2839 14454
rect 12065 14514 12131 14517
rect 14230 14514 14290 14726
rect 19200 14696 20000 14726
rect 12065 14512 14290 14514
rect 12065 14456 12070 14512
rect 12126 14456 14290 14512
rect 12065 14454 14290 14456
rect 15101 14514 15167 14517
rect 19200 14514 20000 14544
rect 15101 14512 20000 14514
rect 15101 14456 15106 14512
rect 15162 14456 20000 14512
rect 15101 14454 20000 14456
rect 12065 14451 12131 14454
rect 15101 14451 15167 14454
rect 19200 14424 20000 14454
rect 0 14242 800 14272
rect 1761 14242 1827 14245
rect 0 14240 1827 14242
rect 0 14184 1766 14240
rect 1822 14184 1827 14240
rect 0 14182 1827 14184
rect 0 14152 800 14182
rect 1761 14179 1827 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 15770 14111 16090 14112
rect 19200 14106 20000 14136
rect 16208 14046 20000 14106
rect 12157 13970 12223 13973
rect 16208 13970 16268 14046
rect 19200 14016 20000 14046
rect 12157 13968 16268 13970
rect 12157 13912 12162 13968
rect 12218 13912 16268 13968
rect 12157 13910 16268 13912
rect 12157 13907 12223 13910
rect 0 13834 800 13864
rect 1761 13834 1827 13837
rect 0 13832 1827 13834
rect 0 13776 1766 13832
rect 1822 13776 1827 13832
rect 0 13774 1827 13776
rect 0 13744 800 13774
rect 1761 13771 1827 13774
rect 15326 13772 15332 13836
rect 15396 13834 15402 13836
rect 19200 13834 20000 13864
rect 15396 13774 20000 13834
rect 15396 13772 15402 13774
rect 19200 13744 20000 13774
rect 6874 13632 7194 13633
rect 0 13562 800 13592
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 2773 13562 2839 13565
rect 0 13560 2839 13562
rect 0 13504 2778 13560
rect 2834 13504 2839 13560
rect 0 13502 2839 13504
rect 0 13472 800 13502
rect 2773 13499 2839 13502
rect 17677 13562 17743 13565
rect 19200 13562 20000 13592
rect 17677 13560 20000 13562
rect 17677 13504 17682 13560
rect 17738 13504 20000 13560
rect 17677 13502 20000 13504
rect 17677 13499 17743 13502
rect 19200 13472 20000 13502
rect 0 13290 800 13320
rect 2773 13290 2839 13293
rect 0 13288 2839 13290
rect 0 13232 2778 13288
rect 2834 13232 2839 13288
rect 0 13230 2839 13232
rect 0 13200 800 13230
rect 2773 13227 2839 13230
rect 16205 13292 16271 13293
rect 16205 13288 16252 13292
rect 16316 13290 16322 13292
rect 16205 13232 16210 13288
rect 16205 13228 16252 13232
rect 16316 13230 16362 13290
rect 16316 13228 16322 13230
rect 16205 13227 16271 13228
rect 16205 13154 16271 13157
rect 19200 13154 20000 13184
rect 16205 13152 20000 13154
rect 16205 13096 16210 13152
rect 16266 13096 20000 13152
rect 16205 13094 20000 13096
rect 16205 13091 16271 13094
rect 3909 13088 4229 13089
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 19200 13064 20000 13094
rect 15770 13023 16090 13024
rect 0 12882 800 12912
rect 3233 12882 3299 12885
rect 0 12880 3299 12882
rect 0 12824 3238 12880
rect 3294 12824 3299 12880
rect 0 12822 3299 12824
rect 0 12792 800 12822
rect 3233 12819 3299 12822
rect 15745 12882 15811 12885
rect 19200 12882 20000 12912
rect 15745 12880 20000 12882
rect 15745 12824 15750 12880
rect 15806 12824 20000 12880
rect 15745 12822 20000 12824
rect 15745 12819 15811 12822
rect 19200 12792 20000 12822
rect 0 12610 800 12640
rect 3785 12610 3851 12613
rect 0 12608 3851 12610
rect 0 12552 3790 12608
rect 3846 12552 3851 12608
rect 0 12550 3851 12552
rect 0 12520 800 12550
rect 3785 12547 3851 12550
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 12479 13125 12480
rect 7833 12474 7899 12477
rect 8845 12474 8911 12477
rect 7833 12472 8911 12474
rect 7833 12416 7838 12472
rect 7894 12416 8850 12472
rect 8906 12416 8911 12472
rect 7833 12414 8911 12416
rect 7833 12411 7899 12414
rect 8845 12411 8911 12414
rect 15193 12474 15259 12477
rect 19200 12474 20000 12504
rect 15193 12472 20000 12474
rect 15193 12416 15198 12472
rect 15254 12416 20000 12472
rect 15193 12414 20000 12416
rect 15193 12411 15259 12414
rect 19200 12384 20000 12414
rect 2589 12338 2655 12341
rect 3693 12338 3759 12341
rect 12065 12338 12131 12341
rect 2589 12336 12131 12338
rect 2589 12280 2594 12336
rect 2650 12280 3698 12336
rect 3754 12280 12070 12336
rect 12126 12280 12131 12336
rect 2589 12278 12131 12280
rect 2589 12275 2655 12278
rect 3693 12275 3759 12278
rect 12065 12275 12131 12278
rect 0 12202 800 12232
rect 4061 12202 4127 12205
rect 0 12200 4127 12202
rect 0 12144 4066 12200
rect 4122 12144 4127 12200
rect 0 12142 4127 12144
rect 0 12112 800 12142
rect 4061 12139 4127 12142
rect 16982 12140 16988 12204
rect 17052 12202 17058 12204
rect 19200 12202 20000 12232
rect 17052 12142 20000 12202
rect 17052 12140 17058 12142
rect 19200 12112 20000 12142
rect 6269 12066 6335 12069
rect 7373 12066 7439 12069
rect 8201 12068 8267 12069
rect 8150 12066 8156 12068
rect 6269 12064 7439 12066
rect 6269 12008 6274 12064
rect 6330 12008 7378 12064
rect 7434 12008 7439 12064
rect 6269 12006 7439 12008
rect 8110 12006 8156 12066
rect 8220 12064 8267 12068
rect 8262 12008 8267 12064
rect 6269 12003 6335 12006
rect 7373 12003 7439 12006
rect 8150 12004 8156 12006
rect 8220 12004 8267 12008
rect 8201 12003 8267 12004
rect 3909 12000 4229 12001
rect 0 11930 800 11960
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 3601 11930 3667 11933
rect 8661 11930 8727 11933
rect 14273 11930 14339 11933
rect 0 11928 3667 11930
rect 0 11872 3606 11928
rect 3662 11872 3667 11928
rect 0 11870 3667 11872
rect 0 11840 800 11870
rect 3601 11867 3667 11870
rect 4662 11928 8727 11930
rect 4662 11872 8666 11928
rect 8722 11872 8727 11928
rect 4662 11870 8727 11872
rect 0 11658 800 11688
rect 4662 11658 4722 11870
rect 8661 11867 8727 11870
rect 10734 11928 14339 11930
rect 10734 11872 14278 11928
rect 14334 11872 14339 11928
rect 10734 11870 14339 11872
rect 4797 11794 4863 11797
rect 8017 11794 8083 11797
rect 9581 11794 9647 11797
rect 4797 11792 9647 11794
rect 4797 11736 4802 11792
rect 4858 11736 8022 11792
rect 8078 11736 9586 11792
rect 9642 11736 9647 11792
rect 4797 11734 9647 11736
rect 4797 11731 4863 11734
rect 8017 11731 8083 11734
rect 9581 11731 9647 11734
rect 0 11598 4722 11658
rect 5993 11658 6059 11661
rect 10734 11658 10794 11870
rect 14273 11867 14339 11870
rect 11789 11794 11855 11797
rect 19200 11794 20000 11824
rect 11789 11792 20000 11794
rect 11789 11736 11794 11792
rect 11850 11736 20000 11792
rect 11789 11734 20000 11736
rect 11789 11731 11855 11734
rect 19200 11704 20000 11734
rect 5993 11656 10794 11658
rect 5993 11600 5998 11656
rect 6054 11600 10794 11656
rect 5993 11598 10794 11600
rect 10961 11658 11027 11661
rect 14089 11658 14155 11661
rect 10961 11656 14155 11658
rect 10961 11600 10966 11656
rect 11022 11600 14094 11656
rect 14150 11600 14155 11656
rect 10961 11598 14155 11600
rect 0 11568 800 11598
rect 5993 11595 6059 11598
rect 10961 11595 11027 11598
rect 14089 11595 14155 11598
rect 15193 11522 15259 11525
rect 17401 11522 17467 11525
rect 19200 11522 20000 11552
rect 15193 11520 20000 11522
rect 15193 11464 15198 11520
rect 15254 11464 17406 11520
rect 17462 11464 20000 11520
rect 15193 11462 20000 11464
rect 15193 11459 15259 11462
rect 17401 11459 17467 11462
rect 6874 11456 7194 11457
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 19200 11432 20000 11462
rect 12805 11391 13125 11392
rect 0 11250 800 11280
rect 4061 11250 4127 11253
rect 0 11248 4127 11250
rect 0 11192 4066 11248
rect 4122 11192 4127 11248
rect 0 11190 4127 11192
rect 0 11160 800 11190
rect 4061 11187 4127 11190
rect 5073 11250 5139 11253
rect 9622 11250 9628 11252
rect 5073 11248 9628 11250
rect 5073 11192 5078 11248
rect 5134 11192 9628 11248
rect 5073 11190 9628 11192
rect 5073 11187 5139 11190
rect 9622 11188 9628 11190
rect 9692 11250 9698 11252
rect 16205 11250 16271 11253
rect 9692 11248 16271 11250
rect 9692 11192 16210 11248
rect 16266 11192 16271 11248
rect 9692 11190 16271 11192
rect 9692 11188 9698 11190
rect 16205 11187 16271 11190
rect 4889 11114 4955 11117
rect 7281 11114 7347 11117
rect 11421 11114 11487 11117
rect 12617 11114 12683 11117
rect 4889 11112 12683 11114
rect 4889 11056 4894 11112
rect 4950 11056 7286 11112
rect 7342 11056 11426 11112
rect 11482 11056 12622 11112
rect 12678 11056 12683 11112
rect 4889 11054 12683 11056
rect 4889 11051 4955 11054
rect 7281 11051 7347 11054
rect 11421 11051 11487 11054
rect 12617 11051 12683 11054
rect 17953 11114 18019 11117
rect 19200 11114 20000 11144
rect 17953 11112 20000 11114
rect 17953 11056 17958 11112
rect 18014 11056 20000 11112
rect 17953 11054 20000 11056
rect 17953 11051 18019 11054
rect 19200 11024 20000 11054
rect 0 10978 800 11008
rect 0 10918 3848 10978
rect 0 10888 800 10918
rect 3788 10706 3848 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 5257 10842 5323 10845
rect 7097 10842 7163 10845
rect 8661 10842 8727 10845
rect 5257 10840 8727 10842
rect 5257 10784 5262 10840
rect 5318 10784 7102 10840
rect 7158 10784 8666 10840
rect 8722 10784 8727 10840
rect 5257 10782 8727 10784
rect 5257 10779 5323 10782
rect 7097 10779 7163 10782
rect 8661 10779 8727 10782
rect 16941 10842 17007 10845
rect 19200 10842 20000 10872
rect 16941 10840 20000 10842
rect 16941 10784 16946 10840
rect 17002 10784 20000 10840
rect 16941 10782 20000 10784
rect 16941 10779 17007 10782
rect 19200 10752 20000 10782
rect 4613 10706 4679 10709
rect 5717 10706 5783 10709
rect 3788 10704 5783 10706
rect 3788 10648 4618 10704
rect 4674 10648 5722 10704
rect 5778 10648 5783 10704
rect 3788 10646 5783 10648
rect 4613 10643 4679 10646
rect 5717 10643 5783 10646
rect 5993 10706 6059 10709
rect 15510 10706 15516 10708
rect 5993 10704 15516 10706
rect 5993 10648 5998 10704
rect 6054 10648 15516 10704
rect 5993 10646 15516 10648
rect 5993 10643 6059 10646
rect 15510 10644 15516 10646
rect 15580 10644 15586 10708
rect 0 10570 800 10600
rect 6453 10570 6519 10573
rect 11789 10570 11855 10573
rect 15469 10570 15535 10573
rect 16849 10570 16915 10573
rect 0 10568 6519 10570
rect 0 10512 6458 10568
rect 6514 10512 6519 10568
rect 0 10510 6519 10512
rect 0 10480 800 10510
rect 6453 10507 6519 10510
rect 6686 10568 11855 10570
rect 6686 10512 11794 10568
rect 11850 10512 11855 10568
rect 6686 10510 11855 10512
rect 5717 10434 5783 10437
rect 6686 10434 6746 10510
rect 11789 10507 11855 10510
rect 12390 10568 15535 10570
rect 12390 10512 15474 10568
rect 15530 10512 15535 10568
rect 12390 10510 15535 10512
rect 5717 10432 6746 10434
rect 5717 10376 5722 10432
rect 5778 10376 6746 10432
rect 5717 10374 6746 10376
rect 7649 10434 7715 10437
rect 8569 10434 8635 10437
rect 7649 10432 8635 10434
rect 7649 10376 7654 10432
rect 7710 10376 8574 10432
rect 8630 10376 8635 10432
rect 7649 10374 8635 10376
rect 5717 10371 5783 10374
rect 7649 10371 7715 10374
rect 8569 10371 8635 10374
rect 9857 10434 9923 10437
rect 12065 10434 12131 10437
rect 9857 10432 12131 10434
rect 9857 10376 9862 10432
rect 9918 10376 12070 10432
rect 12126 10376 12131 10432
rect 9857 10374 12131 10376
rect 9857 10371 9923 10374
rect 12065 10371 12131 10374
rect 6874 10368 7194 10369
rect 0 10298 800 10328
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 4061 10298 4127 10301
rect 12390 10300 12450 10510
rect 15469 10507 15535 10510
rect 15702 10568 16915 10570
rect 15702 10512 16854 10568
rect 16910 10512 16915 10568
rect 15702 10510 16915 10512
rect 15009 10434 15075 10437
rect 15702 10434 15762 10510
rect 16849 10507 16915 10510
rect 15009 10432 15762 10434
rect 15009 10376 15014 10432
rect 15070 10376 15762 10432
rect 15009 10374 15762 10376
rect 16573 10436 16639 10437
rect 16573 10432 16620 10436
rect 16684 10434 16690 10436
rect 17493 10434 17559 10437
rect 19200 10434 20000 10464
rect 16573 10376 16578 10432
rect 15009 10371 15075 10374
rect 16573 10372 16620 10376
rect 16684 10374 16730 10434
rect 17493 10432 20000 10434
rect 17493 10376 17498 10432
rect 17554 10376 20000 10432
rect 17493 10374 20000 10376
rect 16684 10372 16690 10374
rect 16573 10371 16639 10372
rect 17493 10371 17559 10374
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19200 10344 20000 10374
rect 12805 10303 13125 10304
rect 12382 10298 12388 10300
rect 0 10296 4127 10298
rect 0 10240 4066 10296
rect 4122 10240 4127 10296
rect 0 10238 4127 10240
rect 0 10208 800 10238
rect 4061 10235 4127 10238
rect 7790 10238 12388 10298
rect 3049 10162 3115 10165
rect 7790 10162 7850 10238
rect 12382 10236 12388 10238
rect 12452 10236 12458 10300
rect 14457 10298 14523 10301
rect 17401 10298 17467 10301
rect 14457 10296 17467 10298
rect 14457 10240 14462 10296
rect 14518 10240 17406 10296
rect 17462 10240 17467 10296
rect 14457 10238 17467 10240
rect 14457 10235 14523 10238
rect 17401 10235 17467 10238
rect 3049 10160 7850 10162
rect 3049 10104 3054 10160
rect 3110 10104 7850 10160
rect 3049 10102 7850 10104
rect 10685 10162 10751 10165
rect 12157 10162 12223 10165
rect 10685 10160 12223 10162
rect 10685 10104 10690 10160
rect 10746 10104 12162 10160
rect 12218 10104 12223 10160
rect 10685 10102 12223 10104
rect 3049 10099 3115 10102
rect 10685 10099 10751 10102
rect 12157 10099 12223 10102
rect 16389 10162 16455 10165
rect 19200 10162 20000 10192
rect 16389 10160 20000 10162
rect 16389 10104 16394 10160
rect 16450 10104 20000 10160
rect 16389 10102 20000 10104
rect 16389 10099 16455 10102
rect 19200 10072 20000 10102
rect 0 10026 800 10056
rect 2773 10026 2839 10029
rect 0 10024 2839 10026
rect 0 9968 2778 10024
rect 2834 9968 2839 10024
rect 0 9966 2839 9968
rect 0 9936 800 9966
rect 2773 9963 2839 9966
rect 6453 10026 6519 10029
rect 11421 10026 11487 10029
rect 13813 10026 13879 10029
rect 16941 10026 17007 10029
rect 6453 10024 11346 10026
rect 6453 9968 6458 10024
rect 6514 9968 11346 10024
rect 6453 9966 11346 9968
rect 6453 9963 6519 9966
rect 5349 9890 5415 9893
rect 9489 9890 9555 9893
rect 5349 9888 9555 9890
rect 5349 9832 5354 9888
rect 5410 9832 9494 9888
rect 9550 9832 9555 9888
rect 5349 9830 9555 9832
rect 11286 9890 11346 9966
rect 11421 10024 17007 10026
rect 11421 9968 11426 10024
rect 11482 9968 13818 10024
rect 13874 9968 16946 10024
rect 17002 9968 17007 10024
rect 11421 9966 17007 9968
rect 11421 9963 11487 9966
rect 13813 9963 13879 9966
rect 16941 9963 17007 9966
rect 11605 9890 11671 9893
rect 11286 9888 11671 9890
rect 11286 9832 11610 9888
rect 11666 9832 11671 9888
rect 11286 9830 11671 9832
rect 5349 9827 5415 9830
rect 9489 9827 9555 9830
rect 11605 9827 11671 9830
rect 16849 9890 16915 9893
rect 19200 9890 20000 9920
rect 16849 9888 20000 9890
rect 16849 9832 16854 9888
rect 16910 9832 20000 9888
rect 16849 9830 20000 9832
rect 16849 9827 16915 9830
rect 3909 9824 4229 9825
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 19200 9800 20000 9830
rect 15770 9759 16090 9760
rect 6545 9754 6611 9757
rect 7833 9754 7899 9757
rect 8201 9756 8267 9757
rect 6545 9752 7899 9754
rect 6545 9696 6550 9752
rect 6606 9696 7838 9752
rect 7894 9696 7899 9752
rect 6545 9694 7899 9696
rect 6545 9691 6611 9694
rect 7833 9691 7899 9694
rect 8150 9692 8156 9756
rect 8220 9754 8267 9756
rect 12617 9754 12683 9757
rect 14733 9754 14799 9757
rect 15285 9754 15351 9757
rect 16573 9756 16639 9757
rect 16573 9754 16620 9756
rect 8220 9752 8312 9754
rect 8262 9696 8312 9752
rect 8220 9694 8312 9696
rect 12617 9752 15351 9754
rect 12617 9696 12622 9752
rect 12678 9696 14738 9752
rect 14794 9696 15290 9752
rect 15346 9696 15351 9752
rect 12617 9694 15351 9696
rect 16528 9752 16620 9754
rect 16528 9696 16578 9752
rect 16528 9694 16620 9696
rect 8220 9692 8267 9694
rect 8201 9691 8267 9692
rect 12617 9691 12683 9694
rect 14733 9691 14799 9694
rect 15285 9691 15351 9694
rect 16573 9692 16620 9694
rect 16684 9692 16690 9756
rect 16849 9754 16915 9757
rect 17166 9754 17172 9756
rect 16849 9752 17172 9754
rect 16849 9696 16854 9752
rect 16910 9696 17172 9752
rect 16849 9694 17172 9696
rect 16573 9691 16639 9692
rect 16849 9691 16915 9694
rect 17166 9692 17172 9694
rect 17236 9692 17242 9756
rect 0 9618 800 9648
rect 7373 9618 7439 9621
rect 16665 9618 16731 9621
rect 0 9616 16731 9618
rect 0 9560 7378 9616
rect 7434 9560 16670 9616
rect 16726 9560 16731 9616
rect 0 9558 16731 9560
rect 0 9528 800 9558
rect 7373 9555 7439 9558
rect 16665 9555 16731 9558
rect 4061 9482 4127 9485
rect 5901 9482 5967 9485
rect 8477 9482 8543 9485
rect 4061 9480 5967 9482
rect 4061 9424 4066 9480
rect 4122 9424 5906 9480
rect 5962 9424 5967 9480
rect 4061 9422 5967 9424
rect 4061 9419 4127 9422
rect 5901 9419 5967 9422
rect 6732 9480 8543 9482
rect 6732 9424 8482 9480
rect 8538 9424 8543 9480
rect 6732 9422 8543 9424
rect 0 9346 800 9376
rect 6732 9346 6792 9422
rect 8477 9419 8543 9422
rect 10041 9482 10107 9485
rect 10961 9482 11027 9485
rect 10041 9480 11027 9482
rect 10041 9424 10046 9480
rect 10102 9424 10966 9480
rect 11022 9424 11027 9480
rect 10041 9422 11027 9424
rect 10041 9419 10107 9422
rect 10961 9419 11027 9422
rect 12014 9420 12020 9484
rect 12084 9482 12090 9484
rect 12157 9482 12223 9485
rect 12084 9480 12223 9482
rect 12084 9424 12162 9480
rect 12218 9424 12223 9480
rect 12084 9422 12223 9424
rect 12084 9420 12090 9422
rect 12157 9419 12223 9422
rect 12617 9482 12683 9485
rect 13629 9482 13695 9485
rect 12617 9480 13695 9482
rect 12617 9424 12622 9480
rect 12678 9424 13634 9480
rect 13690 9424 13695 9480
rect 12617 9422 13695 9424
rect 12617 9419 12683 9422
rect 13629 9419 13695 9422
rect 15193 9482 15259 9485
rect 19200 9482 20000 9512
rect 15193 9480 20000 9482
rect 15193 9424 15198 9480
rect 15254 9424 20000 9480
rect 15193 9422 20000 9424
rect 15193 9419 15259 9422
rect 19200 9392 20000 9422
rect 0 9286 6792 9346
rect 7373 9346 7439 9349
rect 9581 9346 9647 9349
rect 7373 9344 9647 9346
rect 7373 9288 7378 9344
rect 7434 9288 9586 9344
rect 9642 9288 9647 9344
rect 7373 9286 9647 9288
rect 0 9256 800 9286
rect 7373 9283 7439 9286
rect 9581 9283 9647 9286
rect 10133 9346 10199 9349
rect 11145 9346 11211 9349
rect 10133 9344 11211 9346
rect 10133 9288 10138 9344
rect 10194 9288 11150 9344
rect 11206 9288 11211 9344
rect 10133 9286 11211 9288
rect 10133 9283 10199 9286
rect 11145 9283 11211 9286
rect 13261 9346 13327 9349
rect 16481 9346 16547 9349
rect 13261 9344 16547 9346
rect 13261 9288 13266 9344
rect 13322 9288 16486 9344
rect 16542 9288 16547 9344
rect 13261 9286 16547 9288
rect 13261 9283 13327 9286
rect 16481 9283 16547 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 2681 9210 2747 9213
rect 4245 9210 4311 9213
rect 12249 9210 12315 9213
rect 2681 9208 4311 9210
rect 2681 9152 2686 9208
rect 2742 9152 4250 9208
rect 4306 9152 4311 9208
rect 2681 9150 4311 9152
rect 2681 9147 2747 9150
rect 4245 9147 4311 9150
rect 10366 9208 12315 9210
rect 10366 9152 12254 9208
rect 12310 9152 12315 9208
rect 10366 9150 12315 9152
rect 1669 9074 1735 9077
rect 10366 9076 10426 9150
rect 12249 9147 12315 9150
rect 13537 9210 13603 9213
rect 14089 9210 14155 9213
rect 17125 9210 17191 9213
rect 13537 9208 17191 9210
rect 13537 9152 13542 9208
rect 13598 9152 14094 9208
rect 14150 9152 17130 9208
rect 17186 9152 17191 9208
rect 13537 9150 17191 9152
rect 13537 9147 13603 9150
rect 14089 9147 14155 9150
rect 17125 9147 17191 9150
rect 18229 9210 18295 9213
rect 19200 9210 20000 9240
rect 18229 9208 20000 9210
rect 18229 9152 18234 9208
rect 18290 9152 20000 9208
rect 18229 9150 20000 9152
rect 18229 9147 18295 9150
rect 19200 9120 20000 9150
rect 10358 9074 10364 9076
rect 1669 9072 10364 9074
rect 1669 9016 1674 9072
rect 1730 9016 10364 9072
rect 1669 9014 10364 9016
rect 1669 9011 1735 9014
rect 10358 9012 10364 9014
rect 10428 9012 10434 9076
rect 12341 9074 12407 9077
rect 18597 9074 18663 9077
rect 12341 9072 18663 9074
rect 12341 9016 12346 9072
rect 12402 9016 18602 9072
rect 18658 9016 18663 9072
rect 12341 9014 18663 9016
rect 12341 9011 12407 9014
rect 18597 9011 18663 9014
rect 0 8938 800 8968
rect 3049 8938 3115 8941
rect 0 8936 3115 8938
rect 0 8880 3054 8936
rect 3110 8880 3115 8936
rect 0 8878 3115 8880
rect 0 8848 800 8878
rect 3049 8875 3115 8878
rect 3509 8938 3575 8941
rect 15561 8938 15627 8941
rect 3509 8936 15627 8938
rect 3509 8880 3514 8936
rect 3570 8880 15566 8936
rect 15622 8880 15627 8936
rect 3509 8878 15627 8880
rect 3509 8875 3575 8878
rect 15561 8875 15627 8878
rect 4521 8800 4587 8805
rect 4521 8744 4526 8800
rect 4582 8744 4587 8800
rect 4521 8739 4587 8744
rect 5349 8802 5415 8805
rect 8937 8802 9003 8805
rect 5349 8800 9003 8802
rect 5349 8744 5354 8800
rect 5410 8744 8942 8800
rect 8998 8744 9003 8800
rect 5349 8742 9003 8744
rect 5349 8739 5415 8742
rect 8937 8739 9003 8742
rect 16389 8802 16455 8805
rect 19200 8802 20000 8832
rect 16389 8800 20000 8802
rect 16389 8744 16394 8800
rect 16450 8744 20000 8800
rect 16389 8742 20000 8744
rect 16389 8739 16455 8742
rect 3909 8736 4229 8737
rect 0 8666 800 8696
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 4524 8668 4584 8739
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 19200 8712 20000 8742
rect 15770 8671 16090 8672
rect 4470 8666 4476 8668
rect 0 8606 3848 8666
rect 4394 8606 4476 8666
rect 0 8576 800 8606
rect 3788 8530 3848 8606
rect 4470 8604 4476 8606
rect 4540 8666 4584 8668
rect 8569 8666 8635 8669
rect 4540 8664 8635 8666
rect 4540 8608 8574 8664
rect 8630 8608 8635 8664
rect 4540 8606 8635 8608
rect 4540 8604 4546 8606
rect 8569 8603 8635 8606
rect 6361 8530 6427 8533
rect 8569 8530 8635 8533
rect 3788 8528 8635 8530
rect 3788 8472 6366 8528
rect 6422 8472 8574 8528
rect 8630 8472 8635 8528
rect 3788 8470 8635 8472
rect 6361 8467 6427 8470
rect 8569 8467 8635 8470
rect 11053 8530 11119 8533
rect 13169 8530 13235 8533
rect 11053 8528 13235 8530
rect 11053 8472 11058 8528
rect 11114 8472 13174 8528
rect 13230 8472 13235 8528
rect 11053 8470 13235 8472
rect 11053 8467 11119 8470
rect 13169 8467 13235 8470
rect 16573 8530 16639 8533
rect 19200 8530 20000 8560
rect 16573 8528 20000 8530
rect 16573 8472 16578 8528
rect 16634 8472 20000 8528
rect 16573 8470 20000 8472
rect 16573 8467 16639 8470
rect 19200 8440 20000 8470
rect 0 8394 800 8424
rect 5809 8394 5875 8397
rect 9029 8394 9095 8397
rect 0 8392 5875 8394
rect 0 8336 5814 8392
rect 5870 8336 5875 8392
rect 0 8334 5875 8336
rect 0 8304 800 8334
rect 5809 8331 5875 8334
rect 5950 8392 9095 8394
rect 5950 8336 9034 8392
rect 9090 8336 9095 8392
rect 5950 8334 9095 8336
rect 5257 8258 5323 8261
rect 5950 8258 6010 8334
rect 9029 8331 9095 8334
rect 16113 8394 16179 8397
rect 16982 8394 16988 8396
rect 16113 8392 16988 8394
rect 16113 8336 16118 8392
rect 16174 8336 16988 8392
rect 16113 8334 16988 8336
rect 16113 8331 16179 8334
rect 16982 8332 16988 8334
rect 17052 8332 17058 8396
rect 5257 8256 6010 8258
rect 5257 8200 5262 8256
rect 5318 8200 6010 8256
rect 5257 8198 6010 8200
rect 5257 8195 5323 8198
rect 6874 8192 7194 8193
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 8127 13125 8128
rect 17769 8122 17835 8125
rect 19200 8122 20000 8152
rect 17769 8120 20000 8122
rect 17769 8064 17774 8120
rect 17830 8064 20000 8120
rect 17769 8062 20000 8064
rect 17769 8059 17835 8062
rect 19200 8032 20000 8062
rect 0 7986 800 8016
rect 1761 7986 1827 7989
rect 4245 7986 4311 7989
rect 0 7984 4311 7986
rect 0 7928 1766 7984
rect 1822 7928 4250 7984
rect 4306 7928 4311 7984
rect 0 7926 4311 7928
rect 0 7896 800 7926
rect 1761 7923 1827 7926
rect 4245 7923 4311 7926
rect 5441 7850 5507 7853
rect 3788 7848 5507 7850
rect 3788 7792 5446 7848
rect 5502 7792 5507 7848
rect 3788 7790 5507 7792
rect 0 7714 800 7744
rect 3788 7714 3848 7790
rect 5441 7787 5507 7790
rect 11973 7850 12039 7853
rect 13721 7850 13787 7853
rect 11973 7848 13787 7850
rect 11973 7792 11978 7848
rect 12034 7792 13726 7848
rect 13782 7792 13787 7848
rect 11973 7790 13787 7792
rect 11973 7787 12039 7790
rect 13721 7787 13787 7790
rect 18413 7850 18479 7853
rect 19200 7850 20000 7880
rect 18413 7848 20000 7850
rect 18413 7792 18418 7848
rect 18474 7792 20000 7848
rect 18413 7790 20000 7792
rect 18413 7787 18479 7790
rect 19200 7760 20000 7790
rect 0 7654 3848 7714
rect 0 7624 800 7654
rect 3909 7648 4229 7649
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 15561 7578 15627 7581
rect 11240 7576 15627 7578
rect 11240 7520 15566 7576
rect 15622 7520 15627 7576
rect 11240 7518 15627 7520
rect 11240 7445 11300 7518
rect 15561 7515 15627 7518
rect 9673 7444 9739 7445
rect 9622 7380 9628 7444
rect 9692 7442 9739 7444
rect 9692 7440 9784 7442
rect 9734 7384 9784 7440
rect 9692 7382 9784 7384
rect 11237 7440 11303 7445
rect 11237 7384 11242 7440
rect 11298 7384 11303 7440
rect 9692 7380 9739 7382
rect 9673 7379 9739 7380
rect 11237 7379 11303 7384
rect 15193 7442 15259 7445
rect 19200 7442 20000 7472
rect 15193 7440 20000 7442
rect 15193 7384 15198 7440
rect 15254 7384 20000 7440
rect 15193 7382 20000 7384
rect 15193 7379 15259 7382
rect 19200 7352 20000 7382
rect 0 7306 800 7336
rect 3693 7306 3759 7309
rect 0 7304 3759 7306
rect 0 7248 3698 7304
rect 3754 7248 3759 7304
rect 0 7246 3759 7248
rect 0 7216 800 7246
rect 3693 7243 3759 7246
rect 17861 7306 17927 7309
rect 17861 7304 17970 7306
rect 17861 7248 17866 7304
rect 17922 7248 17970 7304
rect 17861 7243 17970 7248
rect 17910 7170 17970 7243
rect 19200 7170 20000 7200
rect 17910 7110 20000 7170
rect 6874 7104 7194 7105
rect 0 7034 800 7064
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 19200 7080 20000 7110
rect 12805 7039 13125 7040
rect 4889 7034 4955 7037
rect 0 7032 4955 7034
rect 0 6976 4894 7032
rect 4950 6976 4955 7032
rect 0 6974 4955 6976
rect 0 6944 800 6974
rect 4889 6971 4955 6974
rect 11237 7034 11303 7037
rect 12157 7034 12223 7037
rect 11237 7032 12223 7034
rect 11237 6976 11242 7032
rect 11298 6976 12162 7032
rect 12218 6976 12223 7032
rect 11237 6974 12223 6976
rect 11237 6971 11303 6974
rect 12157 6971 12223 6974
rect 3785 6898 3851 6901
rect 2454 6896 3851 6898
rect 2454 6840 3790 6896
rect 3846 6840 3851 6896
rect 2454 6838 3851 6840
rect 0 6762 800 6792
rect 1945 6762 2011 6765
rect 2454 6762 2514 6838
rect 3785 6835 3851 6838
rect 4061 6898 4127 6901
rect 4470 6898 4476 6900
rect 4061 6896 4476 6898
rect 4061 6840 4066 6896
rect 4122 6840 4476 6896
rect 4061 6838 4476 6840
rect 4061 6835 4127 6838
rect 4470 6836 4476 6838
rect 4540 6836 4546 6900
rect 6729 6898 6795 6901
rect 7557 6898 7623 6901
rect 6729 6896 7623 6898
rect 6729 6840 6734 6896
rect 6790 6840 7562 6896
rect 7618 6840 7623 6896
rect 6729 6838 7623 6840
rect 6729 6835 6795 6838
rect 7557 6835 7623 6838
rect 12014 6836 12020 6900
rect 12084 6898 12090 6900
rect 17125 6898 17191 6901
rect 12084 6896 17191 6898
rect 12084 6840 17130 6896
rect 17186 6840 17191 6896
rect 12084 6838 17191 6840
rect 12084 6836 12090 6838
rect 17125 6835 17191 6838
rect 18321 6898 18387 6901
rect 19200 6898 20000 6928
rect 18321 6896 20000 6898
rect 18321 6840 18326 6896
rect 18382 6840 20000 6896
rect 18321 6838 20000 6840
rect 18321 6835 18387 6838
rect 19200 6808 20000 6838
rect 0 6760 2514 6762
rect 0 6704 1950 6760
rect 2006 6704 2514 6760
rect 0 6702 2514 6704
rect 2681 6762 2747 6765
rect 2865 6762 2931 6765
rect 2681 6760 2931 6762
rect 2681 6704 2686 6760
rect 2742 6704 2870 6760
rect 2926 6704 2931 6760
rect 2681 6702 2931 6704
rect 0 6672 800 6702
rect 1945 6699 2011 6702
rect 2681 6699 2747 6702
rect 2865 6699 2931 6702
rect 8937 6762 9003 6765
rect 12985 6762 13051 6765
rect 17217 6762 17283 6765
rect 8937 6760 13051 6762
rect 8937 6704 8942 6760
rect 8998 6704 12990 6760
rect 13046 6704 13051 6760
rect 8937 6702 13051 6704
rect 8937 6699 9003 6702
rect 12985 6699 13051 6702
rect 15564 6760 17283 6762
rect 15564 6704 17222 6760
rect 17278 6704 17283 6760
rect 15564 6702 17283 6704
rect 11237 6626 11303 6629
rect 15326 6626 15332 6628
rect 11237 6624 15332 6626
rect 11237 6568 11242 6624
rect 11298 6568 15332 6624
rect 11237 6566 15332 6568
rect 11237 6563 11303 6566
rect 15326 6564 15332 6566
rect 15396 6626 15402 6628
rect 15564 6626 15624 6702
rect 17217 6699 17283 6702
rect 15396 6566 15624 6626
rect 15396 6564 15402 6566
rect 3909 6560 4229 6561
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 6495 16090 6496
rect 2589 6490 2655 6493
rect 18229 6490 18295 6493
rect 19200 6490 20000 6520
rect 2589 6488 3848 6490
rect 2589 6432 2594 6488
rect 2650 6432 3848 6488
rect 2589 6430 3848 6432
rect 2589 6427 2655 6430
rect 0 6354 800 6384
rect 3417 6354 3483 6357
rect 0 6352 3483 6354
rect 0 6296 3422 6352
rect 3478 6296 3483 6352
rect 0 6294 3483 6296
rect 3788 6354 3848 6430
rect 18229 6488 20000 6490
rect 18229 6432 18234 6488
rect 18290 6432 20000 6488
rect 18229 6430 20000 6432
rect 18229 6427 18295 6430
rect 19200 6400 20000 6430
rect 9121 6354 9187 6357
rect 10409 6356 10475 6357
rect 10358 6354 10364 6356
rect 3788 6352 9187 6354
rect 3788 6296 9126 6352
rect 9182 6296 9187 6352
rect 3788 6294 9187 6296
rect 10318 6294 10364 6354
rect 10428 6352 10475 6356
rect 10470 6296 10475 6352
rect 0 6264 800 6294
rect 3417 6291 3483 6294
rect 9121 6291 9187 6294
rect 10358 6292 10364 6294
rect 10428 6292 10475 6296
rect 10409 6291 10475 6292
rect 10593 6354 10659 6357
rect 13077 6354 13143 6357
rect 10593 6352 13143 6354
rect 10593 6296 10598 6352
rect 10654 6296 13082 6352
rect 13138 6296 13143 6352
rect 10593 6294 13143 6296
rect 10593 6291 10659 6294
rect 13077 6291 13143 6294
rect 3325 6218 3391 6221
rect 11605 6220 11671 6221
rect 3325 6216 8540 6218
rect 3325 6160 3330 6216
rect 3386 6160 8540 6216
rect 3325 6158 8540 6160
rect 3325 6155 3391 6158
rect 0 6082 800 6112
rect 8480 6085 8540 6158
rect 11605 6216 11652 6220
rect 11716 6218 11722 6220
rect 14273 6218 14339 6221
rect 11605 6160 11610 6216
rect 11605 6156 11652 6160
rect 11716 6158 11762 6218
rect 11838 6216 14339 6218
rect 11838 6160 14278 6216
rect 14334 6160 14339 6216
rect 11838 6158 14339 6160
rect 11716 6156 11722 6158
rect 11605 6155 11671 6156
rect 3141 6082 3207 6085
rect 0 6080 3207 6082
rect 0 6024 3146 6080
rect 3202 6024 3207 6080
rect 0 6022 3207 6024
rect 0 5992 800 6022
rect 3141 6019 3207 6022
rect 8477 6080 8543 6085
rect 8477 6024 8482 6080
rect 8538 6024 8543 6080
rect 8477 6019 8543 6024
rect 6874 6016 7194 6017
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 11838 5813 11898 6158
rect 14273 6155 14339 6158
rect 17769 6218 17835 6221
rect 19200 6218 20000 6248
rect 17769 6216 20000 6218
rect 17769 6160 17774 6216
rect 17830 6160 20000 6216
rect 17769 6158 20000 6160
rect 17769 6155 17835 6158
rect 19200 6128 20000 6158
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 5951 13125 5952
rect 4429 5810 4495 5813
rect 4797 5810 4863 5813
rect 4429 5808 4863 5810
rect 4429 5752 4434 5808
rect 4490 5752 4802 5808
rect 4858 5752 4863 5808
rect 4429 5750 4863 5752
rect 4429 5747 4495 5750
rect 4797 5747 4863 5750
rect 6453 5810 6519 5813
rect 11838 5810 11947 5813
rect 6453 5808 12028 5810
rect 6453 5752 6458 5808
rect 6514 5752 11886 5808
rect 11942 5752 12028 5808
rect 6453 5750 12028 5752
rect 6453 5747 6519 5750
rect 11881 5747 11947 5750
rect 12382 5748 12388 5812
rect 12452 5810 12458 5812
rect 14733 5810 14799 5813
rect 12452 5808 14799 5810
rect 12452 5752 14738 5808
rect 14794 5752 14799 5808
rect 12452 5750 14799 5752
rect 12452 5748 12458 5750
rect 14733 5747 14799 5750
rect 17861 5810 17927 5813
rect 19200 5810 20000 5840
rect 17861 5808 20000 5810
rect 17861 5752 17866 5808
rect 17922 5752 20000 5808
rect 17861 5750 20000 5752
rect 17861 5747 17927 5750
rect 19200 5720 20000 5750
rect 0 5674 800 5704
rect 2773 5674 2839 5677
rect 0 5672 2839 5674
rect 0 5616 2778 5672
rect 2834 5616 2839 5672
rect 0 5614 2839 5616
rect 0 5584 800 5614
rect 2773 5611 2839 5614
rect 6637 5674 6703 5677
rect 15377 5674 15443 5677
rect 6637 5672 15443 5674
rect 6637 5616 6642 5672
rect 6698 5616 15382 5672
rect 15438 5616 15443 5672
rect 6637 5614 15443 5616
rect 6637 5611 6703 5614
rect 15377 5611 15443 5614
rect 11053 5538 11119 5541
rect 14825 5538 14891 5541
rect 11053 5536 14891 5538
rect 11053 5480 11058 5536
rect 11114 5480 14830 5536
rect 14886 5480 14891 5536
rect 11053 5478 14891 5480
rect 11053 5475 11119 5478
rect 14825 5475 14891 5478
rect 16573 5538 16639 5541
rect 19200 5538 20000 5568
rect 16573 5536 20000 5538
rect 16573 5480 16578 5536
rect 16634 5480 20000 5536
rect 16573 5478 20000 5480
rect 16573 5475 16639 5478
rect 3909 5472 4229 5473
rect 0 5402 800 5432
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 19200 5448 20000 5478
rect 15770 5407 16090 5408
rect 1577 5402 1643 5405
rect 0 5400 1643 5402
rect 0 5344 1582 5400
rect 1638 5344 1643 5400
rect 0 5342 1643 5344
rect 0 5312 800 5342
rect 1577 5339 1643 5342
rect 7281 5402 7347 5405
rect 7557 5402 7623 5405
rect 7281 5400 7623 5402
rect 7281 5344 7286 5400
rect 7342 5344 7562 5400
rect 7618 5344 7623 5400
rect 7281 5342 7623 5344
rect 7281 5339 7347 5342
rect 7557 5339 7623 5342
rect 10409 5402 10475 5405
rect 12341 5402 12407 5405
rect 12893 5402 12959 5405
rect 10409 5400 12959 5402
rect 10409 5344 10414 5400
rect 10470 5344 12346 5400
rect 12402 5344 12898 5400
rect 12954 5344 12959 5400
rect 10409 5342 12959 5344
rect 10409 5339 10475 5342
rect 12341 5339 12407 5342
rect 12893 5339 12959 5342
rect 0 5130 800 5160
rect 4245 5130 4311 5133
rect 0 5128 4311 5130
rect 0 5072 4250 5128
rect 4306 5072 4311 5128
rect 0 5070 4311 5072
rect 0 5040 800 5070
rect 4245 5067 4311 5070
rect 4613 5130 4679 5133
rect 5257 5130 5323 5133
rect 4613 5128 5323 5130
rect 4613 5072 4618 5128
rect 4674 5072 5262 5128
rect 5318 5072 5323 5128
rect 4613 5070 5323 5072
rect 4613 5067 4679 5070
rect 5257 5067 5323 5070
rect 18229 5130 18295 5133
rect 19200 5130 20000 5160
rect 18229 5128 20000 5130
rect 18229 5072 18234 5128
rect 18290 5072 20000 5128
rect 18229 5070 20000 5072
rect 18229 5067 18295 5070
rect 19200 5040 20000 5070
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 1485 4858 1551 4861
rect 4429 4858 4495 4861
rect 1485 4856 4495 4858
rect 1485 4800 1490 4856
rect 1546 4800 4434 4856
rect 4490 4800 4495 4856
rect 1485 4798 4495 4800
rect 1485 4795 1551 4798
rect 4429 4795 4495 4798
rect 17861 4858 17927 4861
rect 19200 4858 20000 4888
rect 17861 4856 20000 4858
rect 17861 4800 17866 4856
rect 17922 4800 20000 4856
rect 17861 4798 20000 4800
rect 17861 4795 17927 4798
rect 19200 4768 20000 4798
rect 0 4722 800 4752
rect 3969 4722 4035 4725
rect 0 4720 4035 4722
rect 0 4664 3974 4720
rect 4030 4664 4035 4720
rect 0 4662 4035 4664
rect 0 4632 800 4662
rect 3969 4659 4035 4662
rect 12157 4722 12223 4725
rect 14641 4722 14707 4725
rect 12157 4720 14707 4722
rect 12157 4664 12162 4720
rect 12218 4664 14646 4720
rect 14702 4664 14707 4720
rect 12157 4662 14707 4664
rect 12157 4659 12223 4662
rect 14641 4659 14707 4662
rect 3049 4586 3115 4589
rect 7925 4586 7991 4589
rect 8845 4586 8911 4589
rect 3049 4584 8911 4586
rect 3049 4528 3054 4584
rect 3110 4528 7930 4584
rect 7986 4528 8850 4584
rect 8906 4528 8911 4584
rect 3049 4526 8911 4528
rect 3049 4523 3115 4526
rect 7925 4523 7991 4526
rect 8845 4523 8911 4526
rect 0 4450 800 4480
rect 1117 4450 1183 4453
rect 0 4448 1183 4450
rect 0 4392 1122 4448
rect 1178 4392 1183 4448
rect 0 4390 1183 4392
rect 0 4360 800 4390
rect 1117 4387 1183 4390
rect 18229 4450 18295 4453
rect 19200 4450 20000 4480
rect 18229 4448 20000 4450
rect 18229 4392 18234 4448
rect 18290 4392 20000 4448
rect 18229 4390 20000 4392
rect 18229 4387 18295 4390
rect 3909 4384 4229 4385
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19200 4360 20000 4390
rect 15770 4319 16090 4320
rect 11329 4314 11395 4317
rect 11789 4314 11855 4317
rect 11329 4312 11855 4314
rect 11329 4256 11334 4312
rect 11390 4256 11794 4312
rect 11850 4256 11855 4312
rect 11329 4254 11855 4256
rect 11329 4251 11395 4254
rect 11789 4251 11855 4254
rect 1853 4178 1919 4181
rect 9121 4178 9187 4181
rect 1853 4176 9187 4178
rect 1853 4120 1858 4176
rect 1914 4120 9126 4176
rect 9182 4120 9187 4176
rect 1853 4118 9187 4120
rect 1853 4115 1919 4118
rect 9121 4115 9187 4118
rect 10317 4178 10383 4181
rect 12249 4178 12315 4181
rect 10317 4176 12315 4178
rect 10317 4120 10322 4176
rect 10378 4120 12254 4176
rect 12310 4120 12315 4176
rect 10317 4118 12315 4120
rect 10317 4115 10383 4118
rect 12249 4115 12315 4118
rect 18229 4178 18295 4181
rect 19200 4178 20000 4208
rect 18229 4176 20000 4178
rect 18229 4120 18234 4176
rect 18290 4120 20000 4176
rect 18229 4118 20000 4120
rect 18229 4115 18295 4118
rect 19200 4088 20000 4118
rect 0 4042 800 4072
rect 1485 4042 1551 4045
rect 3233 4042 3299 4045
rect 0 3982 1410 4042
rect 0 3952 800 3982
rect 1350 3906 1410 3982
rect 1485 4040 3299 4042
rect 1485 3984 1490 4040
rect 1546 3984 3238 4040
rect 3294 3984 3299 4040
rect 1485 3982 3299 3984
rect 1485 3979 1551 3982
rect 3233 3979 3299 3982
rect 5533 4042 5599 4045
rect 13721 4042 13787 4045
rect 5533 4040 13787 4042
rect 5533 3984 5538 4040
rect 5594 3984 13726 4040
rect 13782 3984 13787 4040
rect 5533 3982 13787 3984
rect 5533 3979 5599 3982
rect 13721 3979 13787 3982
rect 4521 3906 4587 3909
rect 1350 3904 4587 3906
rect 1350 3848 4526 3904
rect 4582 3848 4587 3904
rect 1350 3846 4587 3848
rect 4521 3843 4587 3846
rect 4705 3906 4771 3909
rect 5993 3906 6059 3909
rect 4705 3904 6059 3906
rect 4705 3848 4710 3904
rect 4766 3848 5998 3904
rect 6054 3848 6059 3904
rect 4705 3846 6059 3848
rect 4705 3843 4771 3846
rect 5993 3843 6059 3846
rect 12249 3906 12315 3909
rect 12382 3906 12388 3908
rect 12249 3904 12388 3906
rect 12249 3848 12254 3904
rect 12310 3848 12388 3904
rect 12249 3846 12388 3848
rect 12249 3843 12315 3846
rect 12382 3844 12388 3846
rect 12452 3844 12458 3908
rect 6874 3840 7194 3841
rect 0 3770 800 3800
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 1485 3770 1551 3773
rect 0 3768 1551 3770
rect 0 3712 1490 3768
rect 1546 3712 1551 3768
rect 0 3710 1551 3712
rect 0 3680 800 3710
rect 1485 3707 1551 3710
rect 5073 3770 5139 3773
rect 6453 3770 6519 3773
rect 5073 3768 6519 3770
rect 5073 3712 5078 3768
rect 5134 3712 6458 3768
rect 6514 3712 6519 3768
rect 5073 3710 6519 3712
rect 5073 3707 5139 3710
rect 6453 3707 6519 3710
rect 18229 3770 18295 3773
rect 19200 3770 20000 3800
rect 18229 3768 20000 3770
rect 18229 3712 18234 3768
rect 18290 3712 20000 3768
rect 18229 3710 20000 3712
rect 18229 3707 18295 3710
rect 19200 3680 20000 3710
rect 2221 3634 2287 3637
rect 4981 3634 5047 3637
rect 2221 3632 5047 3634
rect 2221 3576 2226 3632
rect 2282 3576 4986 3632
rect 5042 3576 5047 3632
rect 2221 3574 5047 3576
rect 2221 3571 2287 3574
rect 4981 3571 5047 3574
rect 6085 3634 6151 3637
rect 11697 3634 11763 3637
rect 6085 3632 11763 3634
rect 6085 3576 6090 3632
rect 6146 3576 11702 3632
rect 11758 3576 11763 3632
rect 6085 3574 11763 3576
rect 6085 3571 6151 3574
rect 11697 3571 11763 3574
rect 0 3498 800 3528
rect 2865 3498 2931 3501
rect 13629 3498 13695 3501
rect 0 3496 2931 3498
rect 0 3440 2870 3496
rect 2926 3440 2931 3496
rect 0 3438 2931 3440
rect 0 3408 800 3438
rect 2865 3435 2931 3438
rect 3742 3496 13695 3498
rect 3742 3440 13634 3496
rect 13690 3440 13695 3496
rect 3742 3438 13695 3440
rect 3509 3226 3575 3229
rect 798 3224 3575 3226
rect 798 3168 3514 3224
rect 3570 3168 3575 3224
rect 798 3166 3575 3168
rect 798 3120 858 3166
rect 3509 3163 3575 3166
rect 0 3030 858 3120
rect 3509 3090 3575 3093
rect 3742 3090 3802 3438
rect 13629 3435 13695 3438
rect 19200 3408 20000 3528
rect 5717 3362 5783 3365
rect 7925 3362 7991 3365
rect 11697 3364 11763 3365
rect 5717 3360 7991 3362
rect 5717 3304 5722 3360
rect 5778 3304 7930 3360
rect 7986 3304 7991 3360
rect 5717 3302 7991 3304
rect 5717 3299 5783 3302
rect 7925 3299 7991 3302
rect 11646 3300 11652 3364
rect 11716 3362 11763 3364
rect 11716 3360 11808 3362
rect 11758 3304 11808 3360
rect 11716 3302 11808 3304
rect 11716 3300 11763 3302
rect 11697 3299 11763 3300
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 4429 3226 4495 3229
rect 9489 3226 9555 3229
rect 4429 3224 9555 3226
rect 4429 3168 4434 3224
rect 4490 3168 9494 3224
rect 9550 3168 9555 3224
rect 4429 3166 9555 3168
rect 4429 3163 4495 3166
rect 9489 3163 9555 3166
rect 11145 3226 11211 3229
rect 12014 3226 12020 3228
rect 11145 3224 12020 3226
rect 11145 3168 11150 3224
rect 11206 3168 12020 3224
rect 11145 3166 12020 3168
rect 11145 3163 11211 3166
rect 12014 3164 12020 3166
rect 12084 3164 12090 3228
rect 19200 3136 20000 3256
rect 3509 3088 3802 3090
rect 3509 3032 3514 3088
rect 3570 3032 3802 3088
rect 3509 3030 3802 3032
rect 4061 3090 4127 3093
rect 14733 3090 14799 3093
rect 4061 3088 14799 3090
rect 4061 3032 4066 3088
rect 4122 3032 14738 3088
rect 14794 3032 14799 3088
rect 4061 3030 14799 3032
rect 0 3000 800 3030
rect 3509 3027 3575 3030
rect 4061 3027 4127 3030
rect 14733 3027 14799 3030
rect 16113 3090 16179 3093
rect 16246 3090 16252 3092
rect 16113 3088 16252 3090
rect 16113 3032 16118 3088
rect 16174 3032 16252 3088
rect 16113 3030 16252 3032
rect 16113 3027 16179 3030
rect 16246 3028 16252 3030
rect 16316 3028 16322 3092
rect 1853 2954 1919 2957
rect 13353 2954 13419 2957
rect 1853 2952 13419 2954
rect 1853 2896 1858 2952
rect 1914 2896 13358 2952
rect 13414 2896 13419 2952
rect 1853 2894 13419 2896
rect 1853 2891 1919 2894
rect 13353 2891 13419 2894
rect 0 2818 800 2848
rect 3233 2818 3299 2821
rect 0 2816 3299 2818
rect 0 2760 3238 2816
rect 3294 2760 3299 2816
rect 0 2758 3299 2760
rect 0 2728 800 2758
rect 3233 2755 3299 2758
rect 6874 2752 7194 2753
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 19200 2728 20000 2848
rect 12805 2687 13125 2688
rect 2681 2682 2747 2685
rect 6453 2682 6519 2685
rect 2681 2680 6519 2682
rect 2681 2624 2686 2680
rect 2742 2624 6458 2680
rect 6514 2624 6519 2680
rect 2681 2622 6519 2624
rect 2681 2619 2747 2622
rect 6453 2619 6519 2622
rect 15510 2620 15516 2684
rect 15580 2682 15586 2684
rect 16113 2682 16179 2685
rect 15580 2680 16179 2682
rect 15580 2624 16118 2680
rect 16174 2624 16179 2680
rect 15580 2622 16179 2624
rect 15580 2620 15586 2622
rect 16113 2619 16179 2622
rect 19200 2456 20000 2576
rect 0 2410 800 2440
rect 3877 2410 3943 2413
rect 0 2408 3943 2410
rect 0 2352 3882 2408
rect 3938 2352 3943 2408
rect 0 2350 3943 2352
rect 0 2320 800 2350
rect 3877 2347 3943 2350
rect 3909 2208 4229 2209
rect 0 2138 800 2168
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2143 16090 2144
rect 3693 2138 3759 2141
rect 0 2136 3759 2138
rect 0 2080 3698 2136
rect 3754 2080 3759 2136
rect 0 2078 3759 2080
rect 0 2048 800 2078
rect 3693 2075 3759 2078
rect 19200 2048 20000 2168
rect 0 1866 800 1896
rect 3233 1866 3299 1869
rect 0 1864 3299 1866
rect 0 1808 3238 1864
rect 3294 1808 3299 1864
rect 0 1806 3299 1808
rect 0 1776 800 1806
rect 3233 1803 3299 1806
rect 19200 1776 20000 1896
rect 0 1458 800 1488
rect 4061 1458 4127 1461
rect 0 1456 4127 1458
rect 0 1400 4066 1456
rect 4122 1400 4127 1456
rect 0 1398 4127 1400
rect 0 1368 800 1398
rect 4061 1395 4127 1398
rect 17033 1458 17099 1461
rect 19200 1458 20000 1488
rect 17033 1456 20000 1458
rect 17033 1400 17038 1456
rect 17094 1400 20000 1456
rect 17033 1398 20000 1400
rect 17033 1395 17099 1398
rect 19200 1368 20000 1398
rect 0 1186 800 1216
rect 3141 1186 3207 1189
rect 0 1184 3207 1186
rect 0 1128 3146 1184
rect 3202 1128 3207 1184
rect 0 1126 3207 1128
rect 0 1096 800 1126
rect 3141 1123 3207 1126
rect 15193 1186 15259 1189
rect 19200 1186 20000 1216
rect 15193 1184 20000 1186
rect 15193 1128 15198 1184
rect 15254 1128 20000 1184
rect 15193 1126 20000 1128
rect 15193 1123 15259 1126
rect 19200 1096 20000 1126
rect 0 778 800 808
rect 2865 778 2931 781
rect 0 776 2931 778
rect 0 720 2870 776
rect 2926 720 2931 776
rect 0 718 2931 720
rect 0 688 800 718
rect 2865 715 2931 718
rect 17493 778 17559 781
rect 19200 778 20000 808
rect 17493 776 20000 778
rect 17493 720 17498 776
rect 17554 720 20000 776
rect 17493 718 20000 720
rect 17493 715 17559 718
rect 19200 688 20000 718
rect 0 506 800 536
rect 3417 506 3483 509
rect 0 504 3483 506
rect 0 448 3422 504
rect 3478 448 3483 504
rect 0 446 3483 448
rect 0 416 800 446
rect 3417 443 3483 446
rect 18597 506 18663 509
rect 19200 506 20000 536
rect 18597 504 20000 506
rect 18597 448 18602 504
rect 18658 448 20000 504
rect 18597 446 20000 448
rect 18597 443 18663 446
rect 19200 416 20000 446
rect 0 234 800 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 800 174
rect 2773 171 2839 174
rect 15285 234 15351 237
rect 19200 234 20000 264
rect 15285 232 20000 234
rect 15285 176 15290 232
rect 15346 176 20000 232
rect 15285 174 20000 176
rect 15285 171 15351 174
rect 19200 144 20000 174
<< via3 >>
rect 15516 16764 15580 16828
rect 17172 15404 17236 15468
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 15332 13772 15396 13836
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 16252 13288 16316 13292
rect 16252 13232 16266 13288
rect 16266 13232 16316 13288
rect 16252 13228 16316 13232
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 16988 12140 17052 12204
rect 8156 12064 8220 12068
rect 8156 12008 8206 12064
rect 8206 12008 8220 12064
rect 8156 12004 8220 12008
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 9628 11188 9692 11252
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 15516 10644 15580 10708
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 16620 10432 16684 10436
rect 16620 10376 16634 10432
rect 16634 10376 16684 10432
rect 16620 10372 16684 10376
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 12388 10236 12452 10300
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 8156 9752 8220 9756
rect 8156 9696 8206 9752
rect 8206 9696 8220 9752
rect 8156 9692 8220 9696
rect 16620 9752 16684 9756
rect 16620 9696 16634 9752
rect 16634 9696 16684 9752
rect 16620 9692 16684 9696
rect 17172 9692 17236 9756
rect 12020 9420 12084 9484
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 10364 9012 10428 9076
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 4476 8604 4540 8668
rect 16988 8332 17052 8396
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 9628 7440 9692 7444
rect 9628 7384 9678 7440
rect 9678 7384 9692 7440
rect 9628 7380 9692 7384
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 4476 6836 4540 6900
rect 12020 6836 12084 6900
rect 15332 6564 15396 6628
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 10364 6352 10428 6356
rect 10364 6296 10414 6352
rect 10414 6296 10428 6352
rect 10364 6292 10428 6296
rect 11652 6216 11716 6220
rect 11652 6160 11666 6216
rect 11666 6160 11716 6216
rect 11652 6156 11716 6160
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 12388 5748 12452 5812
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 12388 3844 12452 3908
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 11652 3360 11716 3364
rect 11652 3304 11702 3360
rect 11702 3304 11716 3360
rect 11652 3300 11716 3304
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 12020 3164 12084 3228
rect 16252 3028 16316 3092
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 15516 2620 15580 2684
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 15515 16828 15581 16829
rect 15515 16764 15516 16828
rect 15580 16764 15581 16828
rect 15515 16763 15581 16764
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 8155 12068 8221 12069
rect 8155 12004 8156 12068
rect 8220 12004 8221 12068
rect 8155 12003 8221 12004
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 8158 9757 8218 12003
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9627 11252 9693 11253
rect 9627 11188 9628 11252
rect 9692 11188 9693 11252
rect 9627 11187 9693 11188
rect 8155 9756 8221 9757
rect 8155 9692 8156 9756
rect 8220 9692 8221 9756
rect 8155 9691 8221 9692
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 4475 8668 4541 8669
rect 4475 8604 4476 8668
rect 4540 8604 4541 8668
rect 4475 8603 4541 8604
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 4478 6901 4538 8603
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 9630 7445 9690 11187
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 15331 13836 15397 13837
rect 15331 13772 15332 13836
rect 15396 13772 15397 13836
rect 15331 13771 15397 13772
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12387 10300 12453 10301
rect 12387 10236 12388 10300
rect 12452 10236 12453 10300
rect 12387 10235 12453 10236
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 12019 9484 12085 9485
rect 12019 9420 12020 9484
rect 12084 9420 12085 9484
rect 12019 9419 12085 9420
rect 10363 9076 10429 9077
rect 10363 9012 10364 9076
rect 10428 9012 10429 9076
rect 10363 9011 10429 9012
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9627 7444 9693 7445
rect 9627 7380 9628 7444
rect 9692 7380 9693 7444
rect 9627 7379 9693 7380
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 4475 6900 4541 6901
rect 4475 6836 4476 6900
rect 4540 6836 4541 6900
rect 4475 6835 4541 6836
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 10366 6357 10426 9011
rect 12022 6901 12082 9419
rect 12019 6900 12085 6901
rect 12019 6836 12020 6900
rect 12084 6836 12085 6900
rect 12019 6835 12085 6836
rect 10363 6356 10429 6357
rect 10363 6292 10364 6356
rect 10428 6292 10429 6356
rect 10363 6291 10429 6292
rect 11651 6220 11717 6221
rect 11651 6156 11652 6220
rect 11716 6156 11717 6220
rect 11651 6155 11717 6156
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 11654 3365 11714 6155
rect 11651 3364 11717 3365
rect 11651 3300 11652 3364
rect 11716 3300 11717 3364
rect 11651 3299 11717 3300
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 12022 3229 12082 6835
rect 12390 5813 12450 10235
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 15334 6629 15394 13771
rect 15518 10709 15578 16763
rect 17171 15468 17237 15469
rect 17171 15404 17172 15468
rect 17236 15404 17237 15468
rect 17171 15403 17237 15404
rect 15770 14176 16090 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 15770 13088 16090 14112
rect 16251 13292 16317 13293
rect 16251 13228 16252 13292
rect 16316 13228 16317 13292
rect 16251 13227 16317 13228
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 12000 16090 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 10912 16090 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15515 10708 15581 10709
rect 15515 10644 15516 10708
rect 15580 10644 15581 10708
rect 15515 10643 15581 10644
rect 15331 6628 15397 6629
rect 15331 6564 15332 6628
rect 15396 6564 15397 6628
rect 15331 6563 15397 6564
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12387 5812 12453 5813
rect 12387 5748 12388 5812
rect 12452 5748 12453 5812
rect 12387 5747 12453 5748
rect 12390 3909 12450 5747
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12387 3908 12453 3909
rect 12387 3844 12388 3908
rect 12452 3844 12453 3908
rect 12387 3843 12453 3844
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12019 3228 12085 3229
rect 12019 3164 12020 3228
rect 12084 3164 12085 3228
rect 12019 3163 12085 3164
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 15518 2685 15578 10643
rect 15770 9824 16090 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 8736 16090 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 7648 16090 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 6560 16090 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 5472 16090 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 4384 16090 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15770 3296 16090 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15515 2684 15581 2685
rect 15515 2620 15516 2684
rect 15580 2620 15581 2684
rect 15515 2619 15581 2620
rect 15770 2208 16090 3232
rect 16254 3093 16314 13227
rect 16987 12204 17053 12205
rect 16987 12140 16988 12204
rect 17052 12140 17053 12204
rect 16987 12139 17053 12140
rect 16619 10436 16685 10437
rect 16619 10372 16620 10436
rect 16684 10372 16685 10436
rect 16619 10371 16685 10372
rect 16622 9757 16682 10371
rect 16619 9756 16685 9757
rect 16619 9692 16620 9756
rect 16684 9692 16685 9756
rect 16619 9691 16685 9692
rect 16990 8397 17050 12139
rect 17174 9757 17234 15403
rect 17171 9756 17237 9757
rect 17171 9692 17172 9756
rect 17236 9692 17237 9756
rect 17171 9691 17237 9692
rect 16987 8396 17053 8397
rect 16987 8332 16988 8396
rect 17052 8332 17053 8396
rect 16987 8331 17053 8332
rect 16251 3092 16317 3093
rect 16251 3028 16252 3092
rect 16316 3028 16317 3092
rect 16251 3027 16317 3028
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2128 16090 2144
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608763783
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608763783
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1608763783
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_180
timestamp 1608763783
transform 1 0 17664 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1608763783
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608763783
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1608763783
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1608763783
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1608763783
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608763783
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1608763783
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1608763783
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1608763783
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608763783
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1608763783
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1608763783
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1608763783
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1608763783
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608763783
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1608763783
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1608763783
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608763783
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_23
timestamp 1608763783
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608763783
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1608763783
transform 1 0 1564 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608763783
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1608763783
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_11
timestamp 1608763783
transform 1 0 2116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608763783
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1608763783
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1608763783
transform 1 0 16468 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608763783
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1608763783
transform 1 0 17020 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608763783
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1608763783
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1608763783
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1608763783
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1608763783
transform 1 0 15732 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1608763783
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608763783
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_107
timestamp 1608763783
transform 1 0 10948 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1608763783
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1608763783
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  clk_1_N_FTB01
timestamp 1608763783
transform 1 0 10396 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1608763783
transform 1 0 9384 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1608763783
transform 1 0 9016 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1608763783
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1608763783
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608763783
transform 1 0 6072 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608763783
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_43
timestamp 1608763783
transform 1 0 5060 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_51
timestamp 1608763783
transform 1 0 5796 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_58
timestamp 1608763783
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1608763783
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1608763783
transform 1 0 3956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  clk_2_W_FTB01
timestamp 1608763783
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_W_FTB01
timestamp 1608763783
transform 1 0 2300 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608763783
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1608763783
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1608763783
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_19
timestamp 1608763783
transform 1 0 2852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608763783
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608763783
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_188
timestamp 1608763783
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608763783
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_1_S_FTB01
timestamp 1608763783
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608763783
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1608763783
transform 1 0 17480 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1608763783
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 1608763783
transform 1 0 17480 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1608763783
transform 1 0 18216 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_E_FTB01
timestamp 1608763783
transform 1 0 16928 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1608763783
transform 1 0 16652 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_167
timestamp 1608763783
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608763783
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1608763783
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1608763783
transform 1 0 15732 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1608763783
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1608763783
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_166
timestamp 1608763783
transform 1 0 16376 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1608763783
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_128
timestamp 1608763783
transform 1 0 12880 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_140
timestamp 1608763783
transform 1 0 13984 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1608763783
transform 1 0 11316 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1608763783
transform 1 0 10948 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608763783
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_109
timestamp 1608763783
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1608763783
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1608763783
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_105
timestamp 1608763783
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_116
timestamp 1608763783
transform 1 0 11776 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1608763783
transform 1 0 10304 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1608763783
transform 1 0 9292 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1608763783
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608763783
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_88
timestamp 1608763783
transform 1 0 9200 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_98
timestamp 1608763783
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1608763783
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1608763783
transform 1 0 7820 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1608763783
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_82
timestamp 1608763783
transform 1 0 8648 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1608763783
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1608763783
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1608763783
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608763783
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_42
timestamp 1608763783
transform 1 0 4968 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_54
timestamp 1608763783
transform 1 0 6072 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1608763783
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1608763783
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1608763783
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1608763783
transform 1 0 3036 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608763783
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_30
timestamp 1608763783
transform 1 0 3864 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1608763783
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1608763783
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1608763783
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1608763783
transform 1 0 2944 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1608763783
transform 1 0 2576 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_11
timestamp 1608763783
transform 1 0 2116 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_14
timestamp 1608763783
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_3_E_FTB01
timestamp 1608763783
transform 1 0 1840 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_W_FTB01
timestamp 1608763783
transform 1 0 1564 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608763783
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608763783
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1608763783
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1608763783
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1608763783
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608763783
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1608763783
transform 1 0 18492 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1608763783
transform 1 0 17296 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_174
timestamp 1608763783
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_185
timestamp 1608763783
transform 1 0 18124 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1608763783
transform 1 0 16284 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_E_FTB01
timestamp 1608763783
transform 1 0 15548 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608763783
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1608763783
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1608763783
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1608763783
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608763783
transform 1 0 13892 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_136
timestamp 1608763783
transform 1 0 13616 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1608763783
transform 1 0 11684 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_113
timestamp 1608763783
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_124
timestamp 1608763783
transform 1 0 12512 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1608763783
transform 1 0 10672 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1608763783
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608763783
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1608763783
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1608763783
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1608763783
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1608763783
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1608763783
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1608763783
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 5888 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_44
timestamp 1608763783
transform 1 0 5152 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608763783
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_28
timestamp 1608763783
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608763783
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1608763783
transform 1 0 1840 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1608763783
transform 1 0 2852 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608763783
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1608763783
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1608763783
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_17
timestamp 1608763783
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608763783
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1608763783
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608763783
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608763783
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608763783
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_176
timestamp 1608763783
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1608763783
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 15824 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_S_FTB01
timestamp 1608763783
transform 1 0 15088 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1608763783
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1608763783
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1608763783
transform 1 0 13340 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1608763783
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_142
timestamp 1608763783
transform 1 0 14168 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608763783
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1608763783
transform 1 0 11500 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608763783
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1608763783
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1608763783
transform 1 0 8832 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1608763783
transform 1 0 10672 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp 1608763783
transform 1 0 9660 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_101
timestamp 1608763783
transform 1 0 10396 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1608763783
transform 1 0 7820 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1608763783
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1608763783
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1608763783
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1608763783
transform 1 0 5704 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608763783
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_47
timestamp 1608763783
transform 1 0 5428 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608763783
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1608763783
transform 1 0 3128 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1608763783
transform 1 0 4600 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_31
timestamp 1608763783
transform 1 0 3956 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_37
timestamp 1608763783
transform 1 0 4508 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1608763783
transform 1 0 2116 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608763783
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1608763783
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_20
timestamp 1608763783
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608763783
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1608763783
transform 1 0 17204 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1608763783
transform 1 0 16744 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_174
timestamp 1608763783
transform 1 0 17112 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_184
timestamp 1608763783
transform 1 0 18032 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608763783
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1608763783
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1608763783
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 13248 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_130
timestamp 1608763783
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1608763783
transform 1 0 11316 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1608763783
transform 1 0 12236 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1608763783
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_114
timestamp 1608763783
transform 1 0 11592 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_120
timestamp 1608763783
transform 1 0 12144 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608763783
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608763783
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608763783
transform 1 0 7452 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 7912 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_66
timestamp 1608763783
transform 1 0 7176 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_72
timestamp 1608763783
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 5704 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1608763783
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608763783
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608763783
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608763783
transform 1 0 1656 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 2116 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608763783
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1608763783
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_9
timestamp 1608763783
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608763783
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp 1608763783
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608763783
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1608763783
transform 1 0 16928 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608763783
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_170
timestamp 1608763783
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608763783
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608763783
transform 1 0 16376 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 14720 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_146
timestamp 1608763783
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_164
timestamp 1608763783
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608763783
transform 1 0 14168 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_139
timestamp 1608763783
transform 1 0 13892 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1608763783
transform 1 0 11132 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608763783
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1608763783
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1608763783
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1608763783
transform 1 0 10120 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1608763783
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 8464 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 7820 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1608763783
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_76
timestamp 1608763783
transform 1 0 8096 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1608763783
transform 1 0 5428 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1608763783
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608763783
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_45
timestamp 1608763783
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_56
timestamp 1608763783
transform 1 0 6256 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1608763783
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1608763783
transform 1 0 4416 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1608763783
transform 1 0 3404 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_24
timestamp 1608763783
transform 1 0 3312 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 1608763783
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608763783
transform 1 0 1564 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1608763783
transform 1 0 2116 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608763783
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1608763783
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1608763783
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_20
timestamp 1608763783
transform 1 0 2944 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608763783
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608763783
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1608763783
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1608763783
transform 1 0 18492 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608763783
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1608763783
transform 1 0 17296 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_N_FTB01
timestamp 1608763783
transform 1 0 17204 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608763783
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_173
timestamp 1608763783
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1608763783
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_174
timestamp 1608763783
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_185
timestamp 1608763783
transform 1 0 18124 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 15548 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1608763783
transform 1 0 16284 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1608763783
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608763783
transform 1 0 14996 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1608763783
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608763783
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_149
timestamp 1608763783
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1608763783
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 1608763783
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1608763783
transform 1 0 12972 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1608763783
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1608763783
transform 1 0 13892 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_127
timestamp 1608763783
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_138
timestamp 1608763783
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_136
timestamp 1608763783
transform 1 0 13616 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 12144 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608763783
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608763783
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1608763783
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_118
timestamp 1608763783
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1608763783
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1608763783
transform 1 0 11132 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 11040 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 10764 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_107
timestamp 1608763783
transform 1 0 10948 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_108
timestamp 1608763783
transform 1 0 11040 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 9108 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1608763783
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608763783
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_85
timestamp 1608763783
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_103
timestamp 1608763783
transform 1 0 10580 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1608763783
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_102
timestamp 1608763783
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 7452 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1608763783
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 6992 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_67
timestamp 1608763783
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_73
timestamp 1608763783
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 5060 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 6348 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608763783
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 5428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608763783
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1608763783
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1608763783
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_50
timestamp 1608763783
transform 1 0 5704 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp 1608763783
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_41
timestamp 1608763783
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1608763783
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1608763783
transform 1 0 4048 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608763783
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1608763783
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608763783
transform 1 0 3036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 3588 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_25
timestamp 1608763783
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_30
timestamp 1608763783
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_25
timestamp 1608763783
transform 1 0 3404 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608763783
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 1380 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 1932 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608763783
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608763783
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1608763783
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1608763783
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608763783
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 1608763783
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608763783
transform 1 0 18032 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1608763783
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 16376 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1608763783
transform 1 0 15364 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608763783
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1608763783
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_154
timestamp 1608763783
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_164
timestamp 1608763783
transform 1 0 16192 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 13432 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_132
timestamp 1608763783
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1608763783
transform 1 0 12420 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1608763783
transform 1 0 11408 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1608763783
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_121
timestamp 1608763783
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1608763783
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1608763783
transform 1 0 10672 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608763783
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1608763783
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1608763783
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1608763783
transform 1 0 7912 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1608763783
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_83
timestamp 1608763783
transform 1 0 8740 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608763783
transform 1 0 5704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 6256 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1608763783
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_53
timestamp 1608763783
transform 1 0 5980 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608763783
transform 1 0 3036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608763783
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_25
timestamp 1608763783
transform 1 0 3404 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 1380 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608763783
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_19
timestamp 1608763783
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608763783
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1608763783
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608763783
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1608763783
transform 1 0 16652 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608763783
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_167
timestamp 1608763783
transform 1 0 16468 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1608763783
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1608763783
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608763783
transform 1 0 14536 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 14996 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_149
timestamp 1608763783
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1608763783
transform 1 0 13524 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_132
timestamp 1608763783
transform 1 0 13248 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_144
timestamp 1608763783
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1608763783
transform 1 0 11500 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1608763783
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608763783
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 10028 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1608763783
transform 1 0 9200 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_86
timestamp 1608763783
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1608763783
transform 1 0 7084 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 7544 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_68
timestamp 1608763783
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608763783
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1608763783
transform 1 0 4968 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608763783
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_51
timestamp 1608763783
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1608763783
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1608763783
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1608763783
transform 1 0 3956 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_29
timestamp 1608763783
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_40
timestamp 1608763783
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1608763783
transform 1 0 1656 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 2300 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608763783
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1608763783
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_10
timestamp 1608763783
transform 1 0 2024 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608763783
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608763783
transform 1 0 17940 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1608763783
transform 1 0 16928 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_170
timestamp 1608763783
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1608763783
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_187
timestamp 1608763783
transform 1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608763783
transform 1 0 14628 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608763783
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1608763783
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 12972 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1608763783
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1608763783
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 11316 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1608763783
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1608763783
transform 1 0 10304 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 9660 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608763783
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1608763783
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_99
timestamp 1608763783
transform 1 0 10212 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1608763783
transform 1 0 8372 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_77
timestamp 1608763783
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 5060 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 6716 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1608763783
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1608763783
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608763783
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1608763783
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1608763783
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1608763783
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1608763783
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1608763783
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608763783
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1608763783
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1608763783
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608763783
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1608763783
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608763783
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 17020 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608763783
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_171
timestamp 1608763783
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1608763783
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608763783
transform 1 0 15548 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1608763783
transform 1 0 16008 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_155
timestamp 1608763783
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_160
timestamp 1608763783
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 13892 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1608763783
transform 1 0 12880 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_137
timestamp 1608763783
transform 1 0 13708 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1608763783
transform 1 0 10764 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1608763783
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608763783
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 12604 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_108
timestamp 1608763783
transform 1 0 11040 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1608763783
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1608763783
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 8924 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 7820 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1608763783
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_79
timestamp 1608763783
transform 1 0 8372 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608763783
transform 1 0 6164 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1608763783
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608763783
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1608763783
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608763783
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1608763783
transform 1 0 3864 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 4508 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_28
timestamp 1608763783
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_34
timestamp 1608763783
transform 1 0 4232 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1608763783
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1608763783
transform 1 0 2852 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1608763783
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608763783
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_6
timestamp 1608763783
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_17
timestamp 1608763783
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608763783
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1608763783
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608763783
transform 1 0 18124 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1608763783
transform 1 0 17112 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_172
timestamp 1608763783
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_183
timestamp 1608763783
transform 1 0 17940 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 15456 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608763783
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1608763783
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1608763783
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1608763783
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1608763783
transform 1 0 13892 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 13156 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1608763783
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1608763783
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 11500 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_111
timestamp 1608763783
transform 1 0 11316 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1608763783
transform 1 0 10488 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608763783
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608763783
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_99
timestamp 1608763783
transform 1 0 10212 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1608763783
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1608763783
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1608763783
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1608763783
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1608763783
transform 1 0 6532 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_57
timestamp 1608763783
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608763783
transform 1 0 3036 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608763783
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 4876 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608763783
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 4600 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 3588 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_25
timestamp 1608763783
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1608763783
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_36
timestamp 1608763783
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 1380 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608763783
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1608763783
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608763783
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608763783
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1608763783
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608763783
transform 1 0 17940 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608763783
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1608763783
transform 1 0 16928 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608763783
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1608763783
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_181
timestamp 1608763783
transform 1 0 17756 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_187
timestamp 1608763783
transform 1 0 18308 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1608763783
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 16284 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608763783
transform 1 0 16376 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_164
timestamp 1608763783
transform 1 0 16192 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_160
timestamp 1608763783
transform 1 0 15824 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_164
timestamp 1608763783
transform 1 0 16192 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1608763783
transform 1 0 14996 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1608763783
transform 1 0 15364 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608763783
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608763783
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_154
timestamp 1608763783
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 1608763783
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 12788 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1608763783
transform 1 0 12972 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1608763783
transform 1 0 13984 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 14444 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_143
timestamp 1608763783
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_126
timestamp 1608763783
transform 1 0 12696 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_138
timestamp 1608763783
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1608763783
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 11132 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608763783
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_125
timestamp 1608763783
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_114
timestamp 1608763783
transform 1 0 11592 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_118
timestamp 1608763783
transform 1 0 11960 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608763783
transform 1 0 10028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608763783
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 10120 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1608763783
transform 1 0 10304 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608763783
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 8648 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1608763783
transform 1 0 6900 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1608763783
transform 1 0 7912 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1608763783
transform 1 0 8740 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_72
timestamp 1608763783
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1608763783
transform 1 0 8280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1608763783
transform 1 0 6072 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1608763783
transform 1 0 5060 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 6072 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608763783
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_52
timestamp 1608763783
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_60
timestamp 1608763783
transform 1 0 6624 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_52
timestamp 1608763783
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1608763783
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 4416 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1608763783
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608763783
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_28
timestamp 1608763783
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1608763783
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_34
timestamp 1608763783
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 2760 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1608763783
transform 1 0 2852 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_17
timestamp 1608763783
transform 1 0 2668 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_16
timestamp 1608763783
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1608763783
transform 1 0 1840 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1608763783
transform 1 0 1748 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608763783
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608763783
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1608763783
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1608763783
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1608763783
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608763783
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1608763783
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608763783
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1608763783
transform 1 0 16744 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608763783
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_168
timestamp 1608763783
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_179
timestamp 1608763783
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1608763783
transform 1 0 14536 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 15088 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp 1608763783
transform 1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1608763783
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_132
timestamp 1608763783
transform 1 0 13248 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1608763783
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1608763783
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1608763783
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1608763783
transform 1 0 11316 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608763783
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_109
timestamp 1608763783
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1608763783
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 9016 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_102
timestamp 1608763783
transform 1 0 10488 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1608763783
transform 1 0 7820 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1608763783
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_82
timestamp 1608763783
transform 1 0 8648 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1608763783
transform 1 0 6256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1608763783
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608763783
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1608763783
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608763783
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608763783
transform 1 0 3956 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 4600 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_29
timestamp 1608763783
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_35
timestamp 1608763783
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608763783
transform 1 0 1656 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 2300 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608763783
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1608763783
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_10
timestamp 1608763783
transform 1 0 2024 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608763783
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp 1608763783
transform 1 0 18492 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1608763783
transform 1 0 17112 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_171
timestamp 1608763783
transform 1 0 16836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_183
timestamp 1608763783
transform 1 0 17940 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1608763783
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 16284 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608763783
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1608763783
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1608763783
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 13524 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_131
timestamp 1608763783
transform 1 0 13156 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1608763783
transform 1 0 12328 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 11592 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1608763783
transform 1 0 11224 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_120
timestamp 1608763783
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 9752 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608763783
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1608763783
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1608763783
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 7084 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 8740 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1608763783
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_81
timestamp 1608763783
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1608763783
transform 1 0 5060 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1608763783
transform 1 0 6072 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_52
timestamp 1608763783
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1608763783
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608763783
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_25
timestamp 1608763783
transform 1 0 3404 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1608763783
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608763783
transform 1 0 2024 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608763783
transform 1 0 1472 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1608763783
transform 1 0 2576 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608763783
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1608763783
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_8
timestamp 1608763783
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_14
timestamp 1608763783
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608763783
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1608763783
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608763783
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1608763783
transform 1 0 16928 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608763783
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1608763783
transform 1 0 16652 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1608763783
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 15180 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 14628 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_150
timestamp 1608763783
transform 1 0 14904 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1608763783
transform 1 0 13616 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_133
timestamp 1608763783
transform 1 0 13340 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp 1608763783
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1608763783
transform 1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1608763783
transform 1 0 11316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608763783
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1608763783
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608763783
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1608763783
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1608763783
transform 1 0 10304 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1608763783
transform 1 0 9936 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 8464 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1608763783
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608763783
transform 1 0 6164 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1608763783
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608763783
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_42
timestamp 1608763783
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_53
timestamp 1608763783
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608763783
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763783
transform 1 0 3496 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_24
timestamp 1608763783
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1608763783
transform 1 0 2484 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1608763783
transform 1 0 1472 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608763783
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608763783
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1608763783
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608763783
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1608763783
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608763783
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1608763783
transform 1 0 17020 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_171
timestamp 1608763783
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1608763783
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1608763783
transform 1 0 16008 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608763783
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1608763783
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_160
timestamp 1608763783
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763783
transform 1 0 12880 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_126
timestamp 1608763783
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1608763783
transform 1 0 14352 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 11224 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_108
timestamp 1608763783
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1608763783
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1608763783
transform 1 0 10212 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608763783
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_87
timestamp 1608763783
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1608763783
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1608763783
transform 1 0 7268 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1608763783
transform 1 0 8280 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_top_ipin_0.prog_clk
timestamp 1608763783
transform 1 0 6900 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_66
timestamp 1608763783
transform 1 0 7176 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_76
timestamp 1608763783
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 5244 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_43
timestamp 1608763783
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_61
timestamp 1608763783
transform 1 0 6716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1608763783
transform 1 0 4232 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 3220 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1608763783
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1608763783
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1608763783
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763783
transform 1 0 1380 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608763783
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1608763783
transform 1 0 2852 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608763783
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608763783
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1608763783
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1608763783
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1608763783
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_178
timestamp 1608763783
transform 1 0 17480 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1608763783
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_184
timestamp 1608763783
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1608763783
transform 1 0 16744 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1608763783
transform 1 0 16652 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_167
timestamp 1608763783
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_168
timestamp 1608763783
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 14628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1608763783
transform 1 0 15732 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1608763783
transform 1 0 15640 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1608763783
transform 1 0 14720 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1608763783
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1608763783
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1608763783
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1608763783
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_157
timestamp 1608763783
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1608763783
transform 1 0 13708 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1608763783
transform 1 0 13616 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1608763783
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1608763783
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1608763783
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_136
timestamp 1608763783
transform 1 0 13616 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1608763783
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1608763783
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1608763783
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1608763783
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115
timestamp 1608763783
transform 1 0 11684 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1608763783
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_115
timestamp 1608763783
transform 1 0 11684 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1608763783
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1608763783
transform 1 0 10856 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1608763783
transform 1 0 10856 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763783
transform 1 0 9200 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1608763783
transform 1 0 9844 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1608763783
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1608763783
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1608763783
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_104
timestamp 1608763783
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_85
timestamp 1608763783
transform 1 0 8924 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_104
timestamp 1608763783
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 7912 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1608763783
transform 1 0 7084 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1608763783
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1608763783
transform 1 0 8096 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1608763783
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1608763783
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1608763783
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_74
timestamp 1608763783
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1608763783
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_62
timestamp 1608763783
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 5980 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1608763783
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1608763783
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1608763783
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1608763783
transform 1 0 4968 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1608763783
transform 1 0 5796 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1608763783
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50
timestamp 1608763783
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_51
timestamp 1608763783
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1608763783
transform 1 0 4508 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1608763783
transform 1 0 3864 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1608763783
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1608763783
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1608763783
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36
timestamp 1608763783
transform 1 0 4416 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_28
timestamp 1608763783
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_39
timestamp 1608763783
transform 1 0 4692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1608763783
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1608763783
transform 1 0 2852 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1608763783
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19
timestamp 1608763783
transform 1 0 2852 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_17
timestamp 1608763783
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608763783
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763783
transform 1 0 1932 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1608763783
transform 1 0 1840 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608763783
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608763783
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7
timestamp 1608763783
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1608763783
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1608763783
transform 1 0 1748 0 1 2720
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 13472 800 13592 4 REGIN_FEEDTHROUGH
port 1 nsew
rlabel metal3 s 0 13200 800 13320 4 REGOUT_FEEDTHROUGH
port 2 nsew
rlabel metal2 s 16670 0 16726 800 4 SC_IN_BOT
port 3 nsew
rlabel metal2 s 1950 16200 2006 17000 4 SC_IN_TOP
port 4 nsew
rlabel metal2 s 17590 0 17646 800 4 SC_OUT_BOT
port 5 nsew
rlabel metal2 s 5906 16200 5962 17000 4 SC_OUT_TOP
port 6 nsew
rlabel metal2 s 2134 0 2190 800 4 bottom_grid_pin_0_
port 7 nsew
rlabel metal2 s 11242 0 11298 800 4 bottom_grid_pin_10_
port 8 nsew
rlabel metal2 s 12162 0 12218 800 4 bottom_grid_pin_11_
port 9 nsew
rlabel metal2 s 13082 0 13138 800 4 bottom_grid_pin_12_
port 10 nsew
rlabel metal2 s 13910 0 13966 800 4 bottom_grid_pin_13_
port 11 nsew
rlabel metal2 s 14830 0 14886 800 4 bottom_grid_pin_14_
port 12 nsew
rlabel metal2 s 15750 0 15806 800 4 bottom_grid_pin_15_
port 13 nsew
rlabel metal2 s 3054 0 3110 800 4 bottom_grid_pin_1_
port 14 nsew
rlabel metal2 s 3974 0 4030 800 4 bottom_grid_pin_2_
port 15 nsew
rlabel metal2 s 4894 0 4950 800 4 bottom_grid_pin_3_
port 16 nsew
rlabel metal2 s 5814 0 5870 800 4 bottom_grid_pin_4_
port 17 nsew
rlabel metal2 s 6734 0 6790 800 4 bottom_grid_pin_5_
port 18 nsew
rlabel metal2 s 7562 0 7618 800 4 bottom_grid_pin_6_
port 19 nsew
rlabel metal2 s 8482 0 8538 800 4 bottom_grid_pin_7_
port 20 nsew
rlabel metal2 s 9402 0 9458 800 4 bottom_grid_pin_8_
port 21 nsew
rlabel metal2 s 10322 0 10378 800 4 bottom_grid_pin_9_
port 22 nsew
rlabel metal2 s 386 0 442 800 4 ccff_head
port 23 nsew
rlabel metal2 s 1214 0 1270 800 4 ccff_tail
port 24 nsew
rlabel metal3 s 0 6672 800 6792 4 chanx_left_in[0]
port 25 nsew
rlabel metal3 s 0 9936 800 10056 4 chanx_left_in[10]
port 26 nsew
rlabel metal3 s 0 10208 800 10328 4 chanx_left_in[11]
port 27 nsew
rlabel metal3 s 0 10480 800 10600 4 chanx_left_in[12]
port 28 nsew
rlabel metal3 s 0 10888 800 11008 4 chanx_left_in[13]
port 29 nsew
rlabel metal3 s 0 11160 800 11280 4 chanx_left_in[14]
port 30 nsew
rlabel metal3 s 0 11568 800 11688 4 chanx_left_in[15]
port 31 nsew
rlabel metal3 s 0 11840 800 11960 4 chanx_left_in[16]
port 32 nsew
rlabel metal3 s 0 12112 800 12232 4 chanx_left_in[17]
port 33 nsew
rlabel metal3 s 0 12520 800 12640 4 chanx_left_in[18]
port 34 nsew
rlabel metal3 s 0 12792 800 12912 4 chanx_left_in[19]
port 35 nsew
rlabel metal3 s 0 6944 800 7064 4 chanx_left_in[1]
port 36 nsew
rlabel metal3 s 0 7216 800 7336 4 chanx_left_in[2]
port 37 nsew
rlabel metal3 s 0 7624 800 7744 4 chanx_left_in[3]
port 38 nsew
rlabel metal3 s 0 7896 800 8016 4 chanx_left_in[4]
port 39 nsew
rlabel metal3 s 0 8304 800 8424 4 chanx_left_in[5]
port 40 nsew
rlabel metal3 s 0 8576 800 8696 4 chanx_left_in[6]
port 41 nsew
rlabel metal3 s 0 8848 800 8968 4 chanx_left_in[7]
port 42 nsew
rlabel metal3 s 0 9256 800 9376 4 chanx_left_in[8]
port 43 nsew
rlabel metal3 s 0 9528 800 9648 4 chanx_left_in[9]
port 44 nsew
rlabel metal3 s 0 144 800 264 4 chanx_left_out[0]
port 45 nsew
rlabel metal3 s 0 3408 800 3528 4 chanx_left_out[10]
port 46 nsew
rlabel metal3 s 0 3680 800 3800 4 chanx_left_out[11]
port 47 nsew
rlabel metal3 s 0 3952 800 4072 4 chanx_left_out[12]
port 48 nsew
rlabel metal3 s 0 4360 800 4480 4 chanx_left_out[13]
port 49 nsew
rlabel metal3 s 0 4632 800 4752 4 chanx_left_out[14]
port 50 nsew
rlabel metal3 s 0 5040 800 5160 4 chanx_left_out[15]
port 51 nsew
rlabel metal3 s 0 5312 800 5432 4 chanx_left_out[16]
port 52 nsew
rlabel metal3 s 0 5584 800 5704 4 chanx_left_out[17]
port 53 nsew
rlabel metal3 s 0 5992 800 6112 4 chanx_left_out[18]
port 54 nsew
rlabel metal3 s 0 6264 800 6384 4 chanx_left_out[19]
port 55 nsew
rlabel metal3 s 0 416 800 536 4 chanx_left_out[1]
port 56 nsew
rlabel metal3 s 0 688 800 808 4 chanx_left_out[2]
port 57 nsew
rlabel metal3 s 0 1096 800 1216 4 chanx_left_out[3]
port 58 nsew
rlabel metal3 s 0 1368 800 1488 4 chanx_left_out[4]
port 59 nsew
rlabel metal3 s 0 1776 800 1896 4 chanx_left_out[5]
port 60 nsew
rlabel metal3 s 0 2048 800 2168 4 chanx_left_out[6]
port 61 nsew
rlabel metal3 s 0 2320 800 2440 4 chanx_left_out[7]
port 62 nsew
rlabel metal3 s 0 2728 800 2848 4 chanx_left_out[8]
port 63 nsew
rlabel metal3 s 0 3000 800 3120 4 chanx_left_out[9]
port 64 nsew
rlabel metal3 s 19200 10344 20000 10464 4 chanx_right_in[0]
port 65 nsew
rlabel metal3 s 19200 13744 20000 13864 4 chanx_right_in[10]
port 66 nsew
rlabel metal3 s 19200 14016 20000 14136 4 chanx_right_in[11]
port 67 nsew
rlabel metal3 s 19200 14424 20000 14544 4 chanx_right_in[12]
port 68 nsew
rlabel metal3 s 19200 14696 20000 14816 4 chanx_right_in[13]
port 69 nsew
rlabel metal3 s 19200 15104 20000 15224 4 chanx_right_in[14]
port 70 nsew
rlabel metal3 s 19200 15376 20000 15496 4 chanx_right_in[15]
port 71 nsew
rlabel metal3 s 19200 15784 20000 15904 4 chanx_right_in[16]
port 72 nsew
rlabel metal3 s 19200 16056 20000 16176 4 chanx_right_in[17]
port 73 nsew
rlabel metal3 s 19200 16464 20000 16584 4 chanx_right_in[18]
port 74 nsew
rlabel metal3 s 19200 16736 20000 16856 4 chanx_right_in[19]
port 75 nsew
rlabel metal3 s 19200 10752 20000 10872 4 chanx_right_in[1]
port 76 nsew
rlabel metal3 s 19200 11024 20000 11144 4 chanx_right_in[2]
port 77 nsew
rlabel metal3 s 19200 11432 20000 11552 4 chanx_right_in[3]
port 78 nsew
rlabel metal3 s 19200 11704 20000 11824 4 chanx_right_in[4]
port 79 nsew
rlabel metal3 s 19200 12112 20000 12232 4 chanx_right_in[5]
port 80 nsew
rlabel metal3 s 19200 12384 20000 12504 4 chanx_right_in[6]
port 81 nsew
rlabel metal3 s 19200 12792 20000 12912 4 chanx_right_in[7]
port 82 nsew
rlabel metal3 s 19200 13064 20000 13184 4 chanx_right_in[8]
port 83 nsew
rlabel metal3 s 19200 13472 20000 13592 4 chanx_right_in[9]
port 84 nsew
rlabel metal3 s 19200 3680 20000 3800 4 chanx_right_out[0]
port 85 nsew
rlabel metal3 s 19200 7080 20000 7200 4 chanx_right_out[10]
port 86 nsew
rlabel metal3 s 19200 7352 20000 7472 4 chanx_right_out[11]
port 87 nsew
rlabel metal3 s 19200 7760 20000 7880 4 chanx_right_out[12]
port 88 nsew
rlabel metal3 s 19200 8032 20000 8152 4 chanx_right_out[13]
port 89 nsew
rlabel metal3 s 19200 8440 20000 8560 4 chanx_right_out[14]
port 90 nsew
rlabel metal3 s 19200 8712 20000 8832 4 chanx_right_out[15]
port 91 nsew
rlabel metal3 s 19200 9120 20000 9240 4 chanx_right_out[16]
port 92 nsew
rlabel metal3 s 19200 9392 20000 9512 4 chanx_right_out[17]
port 93 nsew
rlabel metal3 s 19200 9800 20000 9920 4 chanx_right_out[18]
port 94 nsew
rlabel metal3 s 19200 10072 20000 10192 4 chanx_right_out[19]
port 95 nsew
rlabel metal3 s 19200 4088 20000 4208 4 chanx_right_out[1]
port 96 nsew
rlabel metal3 s 19200 4360 20000 4480 4 chanx_right_out[2]
port 97 nsew
rlabel metal3 s 19200 4768 20000 4888 4 chanx_right_out[3]
port 98 nsew
rlabel metal3 s 19200 5040 20000 5160 4 chanx_right_out[4]
port 99 nsew
rlabel metal3 s 19200 5448 20000 5568 4 chanx_right_out[5]
port 100 nsew
rlabel metal3 s 19200 5720 20000 5840 4 chanx_right_out[6]
port 101 nsew
rlabel metal3 s 19200 6128 20000 6248 4 chanx_right_out[7]
port 102 nsew
rlabel metal3 s 19200 6400 20000 6520 4 chanx_right_out[8]
port 103 nsew
rlabel metal3 s 19200 6808 20000 6928 4 chanx_right_out[9]
port 104 nsew
rlabel metal3 s 19200 3408 20000 3528 4 clk_1_E_in
port 105 nsew
rlabel metal2 s 9862 16200 9918 17000 4 clk_1_N_out
port 106 nsew
rlabel metal2 s 18510 0 18566 800 4 clk_1_S_out
port 107 nsew
rlabel metal3 s 0 16736 800 16856 4 clk_1_W_in
port 108 nsew
rlabel metal3 s 19200 3136 20000 3256 4 clk_2_E_in
port 109 nsew
rlabel metal3 s 19200 1368 20000 1488 4 clk_2_E_out
port 110 nsew
rlabel metal3 s 0 16464 800 16584 4 clk_2_W_in
port 111 nsew
rlabel metal3 s 0 14832 800 14952 4 clk_2_W_out
port 112 nsew
rlabel metal3 s 19200 2728 20000 2848 4 clk_3_E_in
port 113 nsew
rlabel metal3 s 19200 1096 20000 1216 4 clk_3_E_out
port 114 nsew
rlabel metal3 s 0 16056 800 16176 4 clk_3_W_in
port 115 nsew
rlabel metal3 s 0 14424 800 14544 4 clk_3_W_out
port 116 nsew
rlabel metal2 s 13910 16200 13966 17000 4 prog_clk_0_N_in
port 117 nsew
rlabel metal2 s 17866 16200 17922 17000 4 prog_clk_0_W_out
port 118 nsew
rlabel metal3 s 19200 2456 20000 2576 4 prog_clk_1_E_in
port 119 nsew
rlabel metal3 s 19200 688 20000 808 4 prog_clk_1_N_out
port 120 nsew
rlabel metal2 s 19430 0 19486 800 4 prog_clk_1_S_out
port 121 nsew
rlabel metal3 s 0 15784 800 15904 4 prog_clk_1_W_in
port 122 nsew
rlabel metal3 s 19200 2048 20000 2168 4 prog_clk_2_E_in
port 123 nsew
rlabel metal3 s 19200 416 20000 536 4 prog_clk_2_E_out
port 124 nsew
rlabel metal3 s 0 15376 800 15496 4 prog_clk_2_W_in
port 125 nsew
rlabel metal3 s 0 14152 800 14272 4 prog_clk_2_W_out
port 126 nsew
rlabel metal3 s 19200 1776 20000 1896 4 prog_clk_3_E_in
port 127 nsew
rlabel metal3 s 19200 144 20000 264 4 prog_clk_3_E_out
port 128 nsew
rlabel metal3 s 0 15104 800 15224 4 prog_clk_3_W_in
port 129 nsew
rlabel metal3 s 0 13744 800 13864 4 prog_clk_3_W_out
port 130 nsew
rlabel metal4 s 3909 2128 4229 14736 4 VPWR
port 131 nsew
rlabel metal4 s 6875 2128 7195 14736 4 VGND
port 132 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 17000
string GDS_FILE /ef/openfpga/openlane/runs/cbx_1__1_/results/magic/cbx_1__1_.gds
string GDS_END 1008916
string GDS_START 78434
<< end >>
