VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__0_
  CLASS BLOCK ;
  FOREIGN cbx_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 120.000 ;
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END bottom_grid_pin_0_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.400 61.840 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 2.400 91.760 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 2.400 94.480 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 2.400 97.200 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 2.400 103.320 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.400 106.720 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 2.400 112.160 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 2.400 115.560 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 2.400 118.280 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 2.400 67.280 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 2.400 76.800 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 2.400 82.240 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 2.400 88.360 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 2.400 2.000 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 2.400 34.640 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.400 37.360 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 2.400 40.760 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 2.400 46.880 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.400 49.600 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.400 52.320 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.400 58.440 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.400 13.560 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 2.400 16.960 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 2.400 19.680 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 61.240 150.000 61.840 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 91.160 150.000 91.760 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 93.880 150.000 94.480 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 96.600 150.000 97.200 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 100.000 150.000 100.600 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 102.720 150.000 103.320 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 106.120 150.000 106.720 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 108.840 150.000 109.440 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 111.560 150.000 112.160 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 114.960 150.000 115.560 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 117.680 150.000 118.280 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 63.960 150.000 64.560 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 66.680 150.000 67.280 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 70.080 150.000 70.680 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 72.800 150.000 73.400 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 76.200 150.000 76.800 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 78.920 150.000 79.520 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 81.640 150.000 82.240 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 85.040 150.000 85.640 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 87.760 150.000 88.360 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 1.400 150.000 2.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 31.320 150.000 31.920 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 34.040 150.000 34.640 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 36.760 150.000 37.360 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 40.160 150.000 40.760 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 42.880 150.000 43.480 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 46.280 150.000 46.880 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 49.000 150.000 49.600 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 51.720 150.000 52.320 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 55.120 150.000 55.720 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 57.840 150.000 58.440 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 4.120 150.000 4.720 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 6.840 150.000 7.440 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 10.240 150.000 10.840 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 12.960 150.000 13.560 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 16.360 150.000 16.960 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 19.080 150.000 19.680 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 21.800 150.000 22.400 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 25.200 150.000 25.800 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 27.920 150.000 28.520 ;
    END
  END chanx_right_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 2.400 ;
    END
  END prog_clk
  PIN top_grid_pin_16_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.690 117.600 4.970 120.000 ;
    END
  END top_grid_pin_16_
  PIN top_grid_pin_17_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 117.600 14.170 120.000 ;
    END
  END top_grid_pin_17_
  PIN top_grid_pin_18_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 117.600 23.370 120.000 ;
    END
  END top_grid_pin_18_
  PIN top_grid_pin_19_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.750 117.600 33.030 120.000 ;
    END
  END top_grid_pin_19_
  PIN top_grid_pin_20_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.950 117.600 42.230 120.000 ;
    END
  END top_grid_pin_20_
  PIN top_grid_pin_21_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.150 117.600 51.430 120.000 ;
    END
  END top_grid_pin_21_
  PIN top_grid_pin_22_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 117.600 61.090 120.000 ;
    END
  END top_grid_pin_22_
  PIN top_grid_pin_23_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 117.600 70.290 120.000 ;
    END
  END top_grid_pin_23_
  PIN top_grid_pin_24_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.670 117.600 79.950 120.000 ;
    END
  END top_grid_pin_24_
  PIN top_grid_pin_25_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 117.600 89.150 120.000 ;
    END
  END top_grid_pin_25_
  PIN top_grid_pin_26_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 117.600 98.350 120.000 ;
    END
  END top_grid_pin_26_
  PIN top_grid_pin_27_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 117.600 108.010 120.000 ;
    END
  END top_grid_pin_27_
  PIN top_grid_pin_28_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.930 117.600 117.210 120.000 ;
    END
  END top_grid_pin_28_
  PIN top_grid_pin_29_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.130 117.600 126.410 120.000 ;
    END
  END top_grid_pin_29_
  PIN top_grid_pin_30_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.790 117.600 136.070 120.000 ;
    END
  END top_grid_pin_30_
  PIN top_grid_pin_31_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 144.990 117.600 145.270 120.000 ;
    END
  END top_grid_pin_31_
  PIN vpwr
    USE POWER ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 29.720 10.640 31.320 109.040 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 54.720 10.640 56.320 109.040 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 108.885 ;
      LAYER met1 ;
        RECT 2.830 9.900 145.290 114.200 ;
      LAYER met2 ;
        RECT 2.850 117.320 4.410 118.165 ;
        RECT 5.250 117.320 13.610 118.165 ;
        RECT 14.450 117.320 22.810 118.165 ;
        RECT 23.650 117.320 32.470 118.165 ;
        RECT 33.310 117.320 41.670 118.165 ;
        RECT 42.510 117.320 50.870 118.165 ;
        RECT 51.710 117.320 60.530 118.165 ;
        RECT 61.370 117.320 69.730 118.165 ;
        RECT 70.570 117.320 79.390 118.165 ;
        RECT 80.230 117.320 88.590 118.165 ;
        RECT 89.430 117.320 97.790 118.165 ;
        RECT 98.630 117.320 107.450 118.165 ;
        RECT 108.290 117.320 116.650 118.165 ;
        RECT 117.490 117.320 125.850 118.165 ;
        RECT 126.690 117.320 135.510 118.165 ;
        RECT 136.350 117.320 144.710 118.165 ;
        RECT 2.850 2.680 145.260 117.320 ;
        RECT 2.850 1.515 18.210 2.680 ;
        RECT 19.050 1.515 55.470 2.680 ;
        RECT 56.310 1.515 93.190 2.680 ;
        RECT 94.030 1.515 130.450 2.680 ;
        RECT 131.290 1.515 145.260 2.680 ;
      LAYER met3 ;
        RECT 2.800 117.280 147.200 118.145 ;
        RECT 2.400 115.960 147.600 117.280 ;
        RECT 2.800 114.560 147.200 115.960 ;
        RECT 2.400 112.560 147.600 114.560 ;
        RECT 2.800 111.160 147.200 112.560 ;
        RECT 2.400 109.840 147.600 111.160 ;
        RECT 2.800 108.440 147.200 109.840 ;
        RECT 2.400 107.120 147.600 108.440 ;
        RECT 2.800 105.720 147.200 107.120 ;
        RECT 2.400 103.720 147.600 105.720 ;
        RECT 2.800 102.320 147.200 103.720 ;
        RECT 2.400 101.000 147.600 102.320 ;
        RECT 2.800 99.600 147.200 101.000 ;
        RECT 2.400 97.600 147.600 99.600 ;
        RECT 2.800 96.200 147.200 97.600 ;
        RECT 2.400 94.880 147.600 96.200 ;
        RECT 2.800 93.480 147.200 94.880 ;
        RECT 2.400 92.160 147.600 93.480 ;
        RECT 2.800 90.760 147.200 92.160 ;
        RECT 2.400 88.760 147.600 90.760 ;
        RECT 2.800 87.360 147.200 88.760 ;
        RECT 2.400 86.040 147.600 87.360 ;
        RECT 2.800 84.640 147.200 86.040 ;
        RECT 2.400 82.640 147.600 84.640 ;
        RECT 2.800 81.240 147.200 82.640 ;
        RECT 2.400 79.920 147.600 81.240 ;
        RECT 2.800 78.520 147.200 79.920 ;
        RECT 2.400 77.200 147.600 78.520 ;
        RECT 2.800 75.800 147.200 77.200 ;
        RECT 2.400 73.800 147.600 75.800 ;
        RECT 2.800 72.400 147.200 73.800 ;
        RECT 2.400 71.080 147.600 72.400 ;
        RECT 2.800 69.680 147.200 71.080 ;
        RECT 2.400 67.680 147.600 69.680 ;
        RECT 2.800 66.280 147.200 67.680 ;
        RECT 2.400 64.960 147.600 66.280 ;
        RECT 2.800 63.560 147.200 64.960 ;
        RECT 2.400 62.240 147.600 63.560 ;
        RECT 2.800 60.840 147.200 62.240 ;
        RECT 2.400 58.840 147.600 60.840 ;
        RECT 2.800 57.440 147.200 58.840 ;
        RECT 2.400 56.120 147.600 57.440 ;
        RECT 2.800 54.720 147.200 56.120 ;
        RECT 2.400 52.720 147.600 54.720 ;
        RECT 2.800 51.320 147.200 52.720 ;
        RECT 2.400 50.000 147.600 51.320 ;
        RECT 2.800 48.600 147.200 50.000 ;
        RECT 2.400 47.280 147.600 48.600 ;
        RECT 2.800 45.880 147.200 47.280 ;
        RECT 2.400 43.880 147.600 45.880 ;
        RECT 2.800 42.480 147.200 43.880 ;
        RECT 2.400 41.160 147.600 42.480 ;
        RECT 2.800 39.760 147.200 41.160 ;
        RECT 2.400 37.760 147.600 39.760 ;
        RECT 2.800 36.360 147.200 37.760 ;
        RECT 2.400 35.040 147.600 36.360 ;
        RECT 2.800 33.640 147.200 35.040 ;
        RECT 2.400 32.320 147.600 33.640 ;
        RECT 2.800 30.920 147.200 32.320 ;
        RECT 2.400 28.920 147.600 30.920 ;
        RECT 2.800 27.520 147.200 28.920 ;
        RECT 2.400 26.200 147.600 27.520 ;
        RECT 2.800 24.800 147.200 26.200 ;
        RECT 2.400 22.800 147.600 24.800 ;
        RECT 2.800 21.400 147.200 22.800 ;
        RECT 2.400 20.080 147.600 21.400 ;
        RECT 2.800 18.680 147.200 20.080 ;
        RECT 2.400 17.360 147.600 18.680 ;
        RECT 2.800 15.960 147.200 17.360 ;
        RECT 2.400 13.960 147.600 15.960 ;
        RECT 2.800 12.560 147.200 13.960 ;
        RECT 2.400 11.240 147.600 12.560 ;
        RECT 2.800 9.840 147.200 11.240 ;
        RECT 2.400 7.840 147.600 9.840 ;
        RECT 2.800 6.440 147.200 7.840 ;
        RECT 2.400 5.120 147.600 6.440 ;
        RECT 2.800 3.720 147.200 5.120 ;
        RECT 2.400 2.400 147.600 3.720 ;
        RECT 2.800 1.535 147.200 2.400 ;
      LAYER met4 ;
        RECT 32.070 10.640 54.320 109.040 ;
        RECT 56.720 10.640 131.320 109.040 ;
      LAYER met5 ;
        RECT 31.860 58.700 64.740 60.300 ;
  END
END cbx_1__0_
END LIBRARY

