magic
tech sky130A
magscale 1 2
timestamp 1606425701
<< locali >>
rect 3893 13243 3927 13413
rect 12173 9435 12207 9605
rect 8309 9027 8343 9129
rect 18981 5695 19015 6613
<< viali >>
rect 1869 14569 1903 14603
rect 2697 14569 2731 14603
rect 1685 14433 1719 14467
rect 2513 14433 2547 14467
rect 15485 14433 15519 14467
rect 15669 14229 15703 14263
rect 2053 14025 2087 14059
rect 3249 14025 3283 14059
rect 6193 14025 6227 14059
rect 14657 14025 14691 14059
rect 15853 14025 15887 14059
rect 7021 13957 7055 13991
rect 1869 13821 1903 13855
rect 3065 13821 3099 13855
rect 6009 13821 6043 13855
rect 6837 13821 6871 13855
rect 13645 13821 13679 13855
rect 14473 13821 14507 13855
rect 15669 13821 15703 13855
rect 13829 13685 13863 13719
rect 1777 13481 1811 13515
rect 2789 13413 2823 13447
rect 3893 13413 3927 13447
rect 1593 13345 1627 13379
rect 2697 13345 2731 13379
rect 2973 13277 3007 13311
rect 4077 13345 4111 13379
rect 15460 13345 15494 13379
rect 17877 13345 17911 13379
rect 3893 13209 3927 13243
rect 2329 13141 2363 13175
rect 15531 13141 15565 13175
rect 18061 13141 18095 13175
rect 1593 12937 1627 12971
rect 16681 12869 16715 12903
rect 2145 12801 2179 12835
rect 6193 12801 6227 12835
rect 1961 12733 1995 12767
rect 2789 12733 2823 12767
rect 5457 12733 5491 12767
rect 5917 12733 5951 12767
rect 7941 12733 7975 12767
rect 12852 12733 12886 12767
rect 14232 12733 14266 12767
rect 14968 12733 15002 12767
rect 15577 12733 15611 12767
rect 16497 12733 16531 12767
rect 17233 12733 17267 12767
rect 3034 12665 3068 12699
rect 8585 12665 8619 12699
rect 2053 12597 2087 12631
rect 4169 12597 4203 12631
rect 4629 12597 4663 12631
rect 5549 12597 5583 12631
rect 6009 12597 6043 12631
rect 6837 12597 6871 12631
rect 12955 12597 12989 12631
rect 14335 12597 14369 12631
rect 15071 12597 15105 12631
rect 15761 12597 15795 12631
rect 17417 12597 17451 12631
rect 2329 12393 2363 12427
rect 2697 12393 2731 12427
rect 6714 12325 6748 12359
rect 1593 12257 1627 12291
rect 4896 12257 4930 12291
rect 8677 12257 8711 12291
rect 8769 12257 8803 12291
rect 12484 12257 12518 12291
rect 13404 12257 13438 12291
rect 14473 12257 14507 12291
rect 15669 12257 15703 12291
rect 16405 12257 16439 12291
rect 17141 12257 17175 12291
rect 17877 12257 17911 12291
rect 2789 12189 2823 12223
rect 2973 12189 3007 12223
rect 4629 12189 4663 12223
rect 6469 12189 6503 12223
rect 8953 12189 8987 12223
rect 16589 12121 16623 12155
rect 1777 12053 1811 12087
rect 6009 12053 6043 12087
rect 7849 12053 7883 12087
rect 8309 12053 8343 12087
rect 12587 12053 12621 12087
rect 13507 12053 13541 12087
rect 14657 12053 14691 12087
rect 15853 12053 15887 12087
rect 17325 12053 17359 12087
rect 18061 12053 18095 12087
rect 4997 11849 5031 11883
rect 15209 11849 15243 11883
rect 8677 11781 8711 11815
rect 2881 11713 2915 11747
rect 3617 11713 3651 11747
rect 5917 11713 5951 11747
rect 6101 11713 6135 11747
rect 9229 11713 9263 11747
rect 13093 11713 13127 11747
rect 14197 11713 14231 11747
rect 1593 11645 1627 11679
rect 2697 11645 2731 11679
rect 6837 11645 6871 11679
rect 15025 11645 15059 11679
rect 15761 11645 15795 11679
rect 16497 11645 16531 11679
rect 17233 11645 17267 11679
rect 3862 11577 3896 11611
rect 7082 11577 7116 11611
rect 12817 11577 12851 11611
rect 14013 11577 14047 11611
rect 1777 11509 1811 11543
rect 2329 11509 2363 11543
rect 2789 11509 2823 11543
rect 5457 11509 5491 11543
rect 5825 11509 5859 11543
rect 8217 11509 8251 11543
rect 9045 11509 9079 11543
rect 9137 11509 9171 11543
rect 12449 11509 12483 11543
rect 12909 11509 12943 11543
rect 13645 11509 13679 11543
rect 14105 11509 14139 11543
rect 15945 11509 15979 11543
rect 16681 11509 16715 11543
rect 17417 11509 17451 11543
rect 1869 11305 1903 11339
rect 2697 11305 2731 11339
rect 3157 11305 3191 11339
rect 4077 11305 4111 11339
rect 4445 11305 4479 11339
rect 15669 11305 15703 11339
rect 16497 11305 16531 11339
rect 3065 11237 3099 11271
rect 7748 11237 7782 11271
rect 5733 11169 5767 11203
rect 6745 11169 6779 11203
rect 10784 11169 10818 11203
rect 12541 11169 12575 11203
rect 12808 11169 12842 11203
rect 14473 11169 14507 11203
rect 16865 11169 16899 11203
rect 17877 11169 17911 11203
rect 1961 11101 1995 11135
rect 2145 11101 2179 11135
rect 3341 11101 3375 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 5825 11101 5859 11135
rect 6009 11101 6043 11135
rect 7481 11101 7515 11135
rect 9689 11101 9723 11135
rect 10517 11101 10551 11135
rect 15761 11101 15795 11135
rect 15853 11101 15887 11135
rect 16957 11101 16991 11135
rect 17049 11101 17083 11135
rect 1501 11033 1535 11067
rect 6929 11033 6963 11067
rect 18061 11033 18095 11067
rect 5365 10965 5399 10999
rect 8861 10965 8895 10999
rect 11897 10965 11931 10999
rect 13921 10965 13955 10999
rect 14657 10965 14691 10999
rect 15301 10965 15335 10999
rect 13001 10761 13035 10795
rect 3801 10693 3835 10727
rect 4353 10693 4387 10727
rect 6837 10693 6871 10727
rect 5273 10625 5307 10659
rect 7481 10625 7515 10659
rect 11161 10625 11195 10659
rect 11345 10625 11379 10659
rect 13553 10625 13587 10659
rect 1685 10557 1719 10591
rect 2421 10557 2455 10591
rect 4537 10557 4571 10591
rect 4997 10557 5031 10591
rect 5825 10557 5859 10591
rect 7205 10557 7239 10591
rect 8033 10557 8067 10591
rect 8861 10557 8895 10591
rect 11069 10557 11103 10591
rect 12817 10557 12851 10591
rect 15393 10557 15427 10591
rect 17233 10557 17267 10591
rect 2688 10489 2722 10523
rect 6101 10489 6135 10523
rect 9128 10489 9162 10523
rect 13820 10489 13854 10523
rect 15660 10489 15694 10523
rect 1869 10421 1903 10455
rect 4629 10421 4663 10455
rect 5089 10421 5123 10455
rect 7297 10421 7331 10455
rect 8217 10421 8251 10455
rect 10241 10421 10275 10455
rect 10701 10421 10735 10455
rect 14933 10421 14967 10455
rect 16773 10421 16807 10455
rect 17417 10421 17451 10455
rect 1593 10217 1627 10251
rect 1961 10217 1995 10251
rect 2789 10217 2823 10251
rect 3157 10217 3191 10251
rect 4997 10217 5031 10251
rect 5365 10217 5399 10251
rect 6193 10217 6227 10251
rect 6561 10217 6595 10251
rect 9781 10217 9815 10251
rect 10149 10217 10183 10251
rect 10977 10217 11011 10251
rect 12541 10217 12575 10251
rect 13369 10217 13403 10251
rect 13737 10217 13771 10251
rect 15853 10217 15887 10251
rect 17233 10217 17267 10251
rect 17693 10217 17727 10251
rect 4353 10149 4387 10183
rect 6653 10149 6687 10183
rect 7840 10149 7874 10183
rect 11437 10149 11471 10183
rect 2053 10081 2087 10115
rect 4077 10081 4111 10115
rect 7573 10081 7607 10115
rect 11345 10081 11379 10115
rect 13829 10081 13863 10115
rect 14632 10081 14666 10115
rect 16221 10081 16255 10115
rect 17601 10081 17635 10115
rect 2237 10013 2271 10047
rect 3249 10013 3283 10047
rect 3341 10013 3375 10047
rect 5457 10013 5491 10047
rect 5641 10013 5675 10047
rect 6837 10013 6871 10047
rect 10241 10013 10275 10047
rect 10333 10013 10367 10047
rect 11621 10013 11655 10047
rect 12633 10013 12667 10047
rect 12725 10013 12759 10047
rect 13921 10013 13955 10047
rect 16313 10013 16347 10047
rect 16497 10013 16531 10047
rect 17785 10013 17819 10047
rect 12173 9945 12207 9979
rect 8953 9877 8987 9911
rect 14703 9877 14737 9911
rect 3709 9673 3743 9707
rect 5457 9673 5491 9707
rect 12449 9673 12483 9707
rect 15669 9673 15703 9707
rect 3249 9605 3283 9639
rect 8861 9605 8895 9639
rect 9781 9605 9815 9639
rect 10701 9605 10735 9639
rect 12173 9605 12207 9639
rect 16773 9605 16807 9639
rect 4261 9537 4295 9571
rect 6101 9537 6135 9571
rect 9413 9537 9447 9571
rect 10425 9537 10459 9571
rect 11253 9537 11287 9571
rect 1869 9469 1903 9503
rect 5365 9469 5399 9503
rect 7021 9469 7055 9503
rect 7288 9469 7322 9503
rect 12081 9469 12115 9503
rect 13001 9537 13035 9571
rect 14289 9537 14323 9571
rect 16129 9537 16163 9571
rect 17325 9537 17359 9571
rect 14556 9469 14590 9503
rect 2136 9401 2170 9435
rect 4169 9401 4203 9435
rect 5825 9401 5859 9435
rect 9229 9401 9263 9435
rect 12173 9401 12207 9435
rect 12909 9401 12943 9435
rect 17141 9401 17175 9435
rect 17233 9401 17267 9435
rect 4077 9333 4111 9367
rect 5181 9333 5215 9367
rect 5917 9333 5951 9367
rect 8401 9333 8435 9367
rect 9321 9333 9355 9367
rect 10149 9333 10183 9367
rect 10241 9333 10275 9367
rect 11069 9333 11103 9367
rect 11161 9333 11195 9367
rect 11897 9333 11931 9367
rect 12817 9333 12851 9367
rect 13645 9333 13679 9367
rect 2973 9129 3007 9163
rect 5457 9129 5491 9163
rect 5917 9129 5951 9163
rect 6377 9129 6411 9163
rect 7113 9129 7147 9163
rect 8309 9129 8343 9163
rect 8401 9129 8435 9163
rect 10517 9129 10551 9163
rect 12357 9129 12391 9163
rect 12909 9129 12943 9163
rect 14105 9129 14139 9163
rect 16681 9129 16715 9163
rect 17141 9129 17175 9163
rect 17509 9129 17543 9163
rect 1860 9061 1894 9095
rect 7573 9061 7607 9095
rect 15568 9061 15602 9095
rect 1593 8993 1627 9027
rect 4344 8993 4378 9027
rect 6285 8993 6319 9027
rect 7481 8993 7515 9027
rect 8309 8993 8343 9027
rect 8769 8993 8803 9027
rect 10057 8993 10091 9027
rect 10977 8993 11011 9027
rect 11244 8993 11278 9027
rect 13277 8993 13311 9027
rect 14289 8993 14323 9027
rect 14473 8993 14507 9027
rect 15301 8993 15335 9027
rect 4077 8925 4111 8959
rect 6561 8925 6595 8959
rect 7665 8925 7699 8959
rect 8861 8925 8895 8959
rect 8953 8925 8987 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 13369 8925 13403 8959
rect 13553 8925 13587 8959
rect 17601 8925 17635 8959
rect 17785 8925 17819 8959
rect 9689 8789 9723 8823
rect 14657 8789 14691 8823
rect 4261 8585 4295 8619
rect 9873 8585 9907 8619
rect 12909 8585 12943 8619
rect 15945 8585 15979 8619
rect 16405 8585 16439 8619
rect 1869 8517 1903 8551
rect 7021 8517 7055 8551
rect 7389 8517 7423 8551
rect 11805 8517 11839 8551
rect 2513 8449 2547 8483
rect 3709 8449 3743 8483
rect 4905 8449 4939 8483
rect 6101 8449 6135 8483
rect 7849 8449 7883 8483
rect 8033 8449 8067 8483
rect 10425 8449 10459 8483
rect 13553 8449 13587 8483
rect 14565 8449 14599 8483
rect 16957 8449 16991 8483
rect 3433 8381 3467 8415
rect 3525 8381 3559 8415
rect 4629 8381 4663 8415
rect 6837 8381 6871 8415
rect 8585 8381 8619 8415
rect 10692 8381 10726 8415
rect 2329 8313 2363 8347
rect 5917 8313 5951 8347
rect 6009 8313 6043 8347
rect 7757 8313 7791 8347
rect 13277 8313 13311 8347
rect 14832 8313 14866 8347
rect 16865 8313 16899 8347
rect 2237 8245 2271 8279
rect 3065 8245 3099 8279
rect 4721 8245 4755 8279
rect 5549 8245 5583 8279
rect 13369 8245 13403 8279
rect 16773 8245 16807 8279
rect 1501 8041 1535 8075
rect 1961 8041 1995 8075
rect 4537 8041 4571 8075
rect 4997 8041 5031 8075
rect 7113 8041 7147 8075
rect 8033 8041 8067 8075
rect 8953 8041 8987 8075
rect 12173 8041 12207 8075
rect 15761 8041 15795 8075
rect 16957 8041 16991 8075
rect 1869 7973 1903 8007
rect 13369 7973 13403 8007
rect 17325 7973 17359 8007
rect 3065 7905 3099 7939
rect 4905 7905 4939 7939
rect 6000 7905 6034 7939
rect 7941 7905 7975 7939
rect 8769 7905 8803 7939
rect 9945 7905 9979 7939
rect 12081 7905 12115 7939
rect 13277 7905 13311 7939
rect 14473 7905 14507 7939
rect 16129 7905 16163 7939
rect 17417 7905 17451 7939
rect 2145 7837 2179 7871
rect 3157 7837 3191 7871
rect 3341 7837 3375 7871
rect 5181 7837 5215 7871
rect 5733 7837 5767 7871
rect 8217 7837 8251 7871
rect 9689 7837 9723 7871
rect 12311 7837 12345 7871
rect 13461 7837 13495 7871
rect 16221 7837 16255 7871
rect 16313 7837 16347 7871
rect 17509 7837 17543 7871
rect 12909 7769 12943 7803
rect 2697 7701 2731 7735
rect 7573 7701 7607 7735
rect 11069 7701 11103 7735
rect 11713 7701 11747 7735
rect 14657 7701 14691 7735
rect 2237 7497 2271 7531
rect 4353 7497 4387 7531
rect 5549 7497 5583 7531
rect 7205 7497 7239 7531
rect 9781 7497 9815 7531
rect 11713 7497 11747 7531
rect 15117 7497 15151 7531
rect 2789 7361 2823 7395
rect 4813 7361 4847 7395
rect 4997 7361 5031 7395
rect 6009 7361 6043 7395
rect 6193 7361 6227 7395
rect 7849 7361 7883 7395
rect 13093 7361 13127 7395
rect 1501 7293 1535 7327
rect 2605 7293 2639 7327
rect 2697 7293 2731 7327
rect 3433 7293 3467 7327
rect 5917 7293 5951 7327
rect 7573 7293 7607 7327
rect 8401 7293 8435 7327
rect 10333 7293 10367 7327
rect 10600 7293 10634 7327
rect 12817 7293 12851 7327
rect 13737 7293 13771 7327
rect 15577 7293 15611 7327
rect 7665 7225 7699 7259
rect 8646 7225 8680 7259
rect 12909 7225 12943 7259
rect 14004 7225 14038 7259
rect 15844 7225 15878 7259
rect 1685 7157 1719 7191
rect 3617 7157 3651 7191
rect 4721 7157 4755 7191
rect 12449 7157 12483 7191
rect 16957 7157 16991 7191
rect 2789 6953 2823 6987
rect 5457 6953 5491 6987
rect 6377 6953 6411 6987
rect 7113 6953 7147 6987
rect 7481 6953 7515 6987
rect 11989 6953 12023 6987
rect 12817 6953 12851 6987
rect 13185 6953 13219 6987
rect 14381 6953 14415 6987
rect 15669 6953 15703 6987
rect 17049 6953 17083 6987
rect 3157 6885 3191 6919
rect 8769 6885 8803 6919
rect 10793 6885 10827 6919
rect 17141 6885 17175 6919
rect 1685 6817 1719 6851
rect 4333 6817 4367 6851
rect 6285 6817 6319 6851
rect 7573 6817 7607 6851
rect 9689 6817 9723 6851
rect 10885 6817 10919 6851
rect 12081 6817 12115 6851
rect 17877 6817 17911 6851
rect 3249 6749 3283 6783
rect 3433 6749 3467 6783
rect 4077 6749 4111 6783
rect 6561 6749 6595 6783
rect 7665 6749 7699 6783
rect 8861 6749 8895 6783
rect 8953 6749 8987 6783
rect 10977 6749 11011 6783
rect 12265 6749 12299 6783
rect 13277 6749 13311 6783
rect 13369 6749 13403 6783
rect 14473 6749 14507 6783
rect 14657 6749 14691 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 17233 6749 17267 6783
rect 10425 6681 10459 6715
rect 16681 6681 16715 6715
rect 1869 6613 1903 6647
rect 5917 6613 5951 6647
rect 8401 6613 8435 6647
rect 9873 6613 9907 6647
rect 11621 6613 11655 6647
rect 14013 6613 14047 6647
rect 15301 6613 15335 6647
rect 18061 6613 18095 6647
rect 18981 6613 19015 6647
rect 3801 6409 3835 6443
rect 6837 6409 6871 6443
rect 8033 6409 8067 6443
rect 11161 6409 11195 6443
rect 15945 6409 15979 6443
rect 15485 6341 15519 6375
rect 2421 6273 2455 6307
rect 7481 6273 7515 6307
rect 8493 6273 8527 6307
rect 8585 6273 8619 6307
rect 9229 6273 9263 6307
rect 11621 6273 11655 6307
rect 11805 6273 11839 6307
rect 12541 6273 12575 6307
rect 13553 6273 13587 6307
rect 16497 6273 16531 6307
rect 1685 6205 1719 6239
rect 4629 6205 4663 6239
rect 4896 6205 4930 6239
rect 6653 6205 6687 6239
rect 7205 6205 7239 6239
rect 9496 6205 9530 6239
rect 11529 6205 11563 6239
rect 14105 6205 14139 6239
rect 17233 6205 17267 6239
rect 2666 6137 2700 6171
rect 12633 6137 12667 6171
rect 14372 6137 14406 6171
rect 16313 6137 16347 6171
rect 1869 6069 1903 6103
rect 6009 6069 6043 6103
rect 6469 6069 6503 6103
rect 7297 6069 7331 6103
rect 8401 6069 8435 6103
rect 10609 6069 10643 6103
rect 16405 6069 16439 6103
rect 17417 6069 17451 6103
rect 3249 5865 3283 5899
rect 4077 5865 4111 5899
rect 12909 5865 12943 5899
rect 16497 5865 16531 5899
rect 17325 5865 17359 5899
rect 17693 5865 17727 5899
rect 3157 5797 3191 5831
rect 6552 5797 6586 5831
rect 9137 5797 9171 5831
rect 13614 5797 13648 5831
rect 17785 5797 17819 5831
rect 1685 5729 1719 5763
rect 4445 5729 4479 5763
rect 5549 5729 5583 5763
rect 8769 5729 8803 5763
rect 9945 5729 9979 5763
rect 11796 5729 11830 5763
rect 13369 5729 13403 5763
rect 15393 5729 15427 5763
rect 1869 5661 1903 5695
rect 3433 5661 3467 5695
rect 4537 5661 4571 5695
rect 4629 5661 4663 5695
rect 6285 5661 6319 5695
rect 8401 5661 8435 5695
rect 9689 5661 9723 5695
rect 11529 5661 11563 5695
rect 16589 5661 16623 5695
rect 16681 5661 16715 5695
rect 17877 5661 17911 5695
rect 18981 5661 19015 5695
rect 2789 5593 2823 5627
rect 5733 5525 5767 5559
rect 7665 5525 7699 5559
rect 11069 5525 11103 5559
rect 14749 5525 14783 5559
rect 15577 5525 15611 5559
rect 16129 5525 16163 5559
rect 1869 5321 1903 5355
rect 3709 5321 3743 5355
rect 9505 5321 9539 5355
rect 9965 5321 9999 5355
rect 15485 5321 15519 5355
rect 16681 5321 16715 5355
rect 6285 5253 6319 5287
rect 7297 5253 7331 5287
rect 12725 5253 12759 5287
rect 4353 5185 4387 5219
rect 13369 5185 13403 5219
rect 14197 5185 14231 5219
rect 16037 5185 16071 5219
rect 17233 5185 17267 5219
rect 1685 5117 1719 5151
rect 2605 5117 2639 5151
rect 4077 5117 4111 5151
rect 4905 5117 4939 5151
rect 6837 5117 6871 5151
rect 7205 5117 7239 5151
rect 8125 5117 8159 5151
rect 10149 5117 10183 5151
rect 10241 5117 10275 5151
rect 12541 5117 12575 5151
rect 15853 5117 15887 5151
rect 17141 5117 17175 5151
rect 2881 5049 2915 5083
rect 5150 5049 5184 5083
rect 8392 5049 8426 5083
rect 10486 5049 10520 5083
rect 13461 5049 13495 5083
rect 14841 5049 14875 5083
rect 17049 5049 17083 5083
rect 4169 4981 4203 5015
rect 11621 4981 11655 5015
rect 15945 4981 15979 5015
rect 1869 4777 1903 4811
rect 2605 4777 2639 4811
rect 4905 4777 4939 4811
rect 5641 4777 5675 4811
rect 9045 4777 9079 4811
rect 16865 4777 16899 4811
rect 17233 4777 17267 4811
rect 6009 4709 6043 4743
rect 11161 4709 11195 4743
rect 11989 4709 12023 4743
rect 12081 4709 12115 4743
rect 13737 4709 13771 4743
rect 13829 4709 13863 4743
rect 15485 4709 15519 4743
rect 16405 4709 16439 4743
rect 1685 4641 1719 4675
rect 2421 4641 2455 4675
rect 3157 4641 3191 4675
rect 4813 4641 4847 4675
rect 6929 4641 6963 4675
rect 7932 4641 7966 4675
rect 9689 4641 9723 4675
rect 10793 4641 10827 4675
rect 5089 4573 5123 4607
rect 6101 4573 6135 4607
rect 6193 4573 6227 4607
rect 7665 4573 7699 4607
rect 13001 4573 13035 4607
rect 14381 4573 14415 4607
rect 15393 4573 15427 4607
rect 17325 4573 17359 4607
rect 17417 4573 17451 4607
rect 10425 4505 10459 4539
rect 3341 4437 3375 4471
rect 4445 4437 4479 4471
rect 7113 4437 7147 4471
rect 9873 4437 9907 4471
rect 1869 4233 1903 4267
rect 9137 4165 9171 4199
rect 9689 4165 9723 4199
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 5733 4097 5767 4131
rect 6837 4097 6871 4131
rect 12909 4097 12943 4131
rect 13369 4097 13403 4131
rect 14933 4097 14967 4131
rect 16129 4097 16163 4131
rect 16957 4097 16991 4131
rect 1685 4029 1719 4063
rect 2409 4029 2443 4063
rect 3157 4029 3191 4063
rect 5549 4029 5583 4063
rect 9505 4029 9539 4063
rect 10333 4029 10367 4063
rect 2145 3961 2179 3995
rect 7104 3961 7138 3995
rect 10600 3961 10634 3995
rect 13001 3961 13035 3995
rect 14473 3961 14507 3995
rect 14565 3961 14599 3995
rect 16221 3961 16255 3995
rect 2605 3893 2639 3927
rect 3341 3893 3375 3927
rect 3985 3893 4019 3927
rect 4353 3893 4387 3927
rect 5181 3893 5215 3927
rect 5641 3893 5675 3927
rect 8217 3893 8251 3927
rect 11713 3893 11747 3927
rect 2145 3689 2179 3723
rect 5457 3689 5491 3723
rect 7297 3689 7331 3723
rect 7757 3689 7791 3723
rect 15485 3689 15519 3723
rect 15853 3689 15887 3723
rect 16681 3689 16715 3723
rect 18061 3689 18095 3723
rect 6184 3621 6218 3655
rect 9137 3621 9171 3655
rect 11437 3621 11471 3655
rect 12357 3621 12391 3655
rect 12909 3621 12943 3655
rect 13001 3621 13035 3655
rect 1685 3553 1719 3587
rect 2881 3553 2915 3587
rect 4077 3553 4111 3587
rect 4344 3553 4378 3587
rect 5917 3553 5951 3587
rect 8401 3553 8435 3587
rect 8769 3553 8803 3587
rect 10425 3553 10459 3587
rect 14473 3553 14507 3587
rect 15945 3553 15979 3587
rect 17049 3553 17083 3587
rect 17141 3553 17175 3587
rect 17877 3553 17911 3587
rect 3065 3485 3099 3519
rect 10793 3485 10827 3519
rect 11345 3485 11379 3519
rect 13737 3485 13771 3519
rect 16129 3485 16163 3519
rect 17233 3485 17267 3519
rect 1869 3417 1903 3451
rect 10057 3417 10091 3451
rect 14657 3349 14691 3383
rect 5457 3145 5491 3179
rect 6193 3077 6227 3111
rect 7389 3077 7423 3111
rect 17463 3077 17497 3111
rect 8861 3009 8895 3043
rect 9781 3009 9815 3043
rect 10425 3009 10459 3043
rect 11253 3009 11287 3043
rect 13001 3009 13035 3043
rect 15301 3009 15335 3043
rect 15853 3009 15887 3043
rect 16865 3009 16899 3043
rect 1501 2941 1535 2975
rect 2421 2941 2455 2975
rect 3341 2941 3375 2975
rect 4261 2941 4295 2975
rect 5273 2941 5307 2975
rect 6009 2941 6043 2975
rect 6837 2941 6871 2975
rect 7205 2941 7239 2975
rect 8033 2941 8067 2975
rect 17360 2941 17394 2975
rect 1777 2873 1811 2907
rect 2697 2873 2731 2907
rect 3617 2873 3651 2907
rect 4537 2873 4571 2907
rect 8953 2873 8987 2907
rect 10517 2873 10551 2907
rect 12725 2873 12759 2907
rect 12817 2873 12851 2907
rect 14289 2873 14323 2907
rect 14381 2873 14415 2907
rect 15945 2873 15979 2907
rect 8217 2805 8251 2839
rect 2697 2601 2731 2635
rect 5549 2601 5583 2635
rect 11989 2601 12023 2635
rect 17693 2601 17727 2635
rect 10241 2533 10275 2567
rect 10333 2533 10367 2567
rect 11253 2533 11287 2567
rect 13369 2533 13403 2567
rect 14289 2533 14323 2567
rect 15669 2533 15703 2567
rect 1593 2465 1627 2499
rect 2513 2465 2547 2499
rect 3249 2465 3283 2499
rect 4077 2465 4111 2499
rect 5365 2465 5399 2499
rect 6101 2465 6135 2499
rect 7297 2465 7331 2499
rect 8493 2465 8527 2499
rect 11805 2465 11839 2499
rect 14816 2465 14850 2499
rect 17509 2465 17543 2499
rect 1777 2397 1811 2431
rect 7665 2397 7699 2431
rect 8125 2397 8159 2431
rect 8861 2397 8895 2431
rect 13277 2397 13311 2431
rect 15577 2397 15611 2431
rect 16497 2397 16531 2431
rect 6285 2329 6319 2363
rect 6929 2329 6963 2363
rect 14887 2329 14921 2363
rect 3433 2261 3467 2295
rect 4261 2261 4295 2295
<< metal1 >>
rect 3694 15240 3700 15292
rect 3752 15280 3758 15292
rect 5994 15280 6000 15292
rect 3752 15252 6000 15280
rect 3752 15240 3758 15252
rect 5994 15240 6000 15252
rect 6052 15240 6058 15292
rect 4062 15172 4068 15224
rect 4120 15212 4126 15224
rect 8110 15212 8116 15224
rect 4120 15184 8116 15212
rect 4120 15172 4126 15184
rect 8110 15172 8116 15184
rect 8168 15172 8174 15224
rect 12158 15172 12164 15224
rect 12216 15212 12222 15224
rect 15930 15212 15936 15224
rect 12216 15184 15936 15212
rect 12216 15172 12222 15184
rect 15930 15172 15936 15184
rect 15988 15172 15994 15224
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 934 14560 940 14612
rect 992 14600 998 14612
rect 1857 14603 1915 14609
rect 1857 14600 1869 14603
rect 992 14572 1869 14600
rect 992 14560 998 14572
rect 1857 14569 1869 14572
rect 1903 14569 1915 14603
rect 1857 14563 1915 14569
rect 2222 14560 2228 14612
rect 2280 14600 2286 14612
rect 2685 14603 2743 14609
rect 2685 14600 2697 14603
rect 2280 14572 2697 14600
rect 2280 14560 2286 14572
rect 2685 14569 2697 14572
rect 2731 14569 2743 14603
rect 2685 14563 2743 14569
rect 2774 14492 2780 14544
rect 2832 14532 2838 14544
rect 13630 14532 13636 14544
rect 2832 14504 13636 14532
rect 2832 14492 2838 14504
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14433 1731 14467
rect 1673 14427 1731 14433
rect 2501 14467 2559 14473
rect 2501 14433 2513 14467
rect 2547 14464 2559 14467
rect 15010 14464 15016 14476
rect 2547 14436 15016 14464
rect 2547 14433 2559 14436
rect 2501 14427 2559 14433
rect 1688 14396 1716 14427
rect 15010 14424 15016 14436
rect 15068 14424 15074 14476
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14464 15531 14467
rect 15746 14464 15752 14476
rect 15519 14436 15752 14464
rect 15519 14433 15531 14436
rect 15473 14427 15531 14433
rect 15746 14424 15752 14436
rect 15804 14464 15810 14476
rect 16298 14464 16304 14476
rect 15804 14436 16304 14464
rect 15804 14424 15810 14436
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 12250 14396 12256 14408
rect 1688 14368 12256 14396
rect 12250 14356 12256 14368
rect 12308 14396 12314 14408
rect 17678 14396 17684 14408
rect 12308 14368 17684 14396
rect 12308 14356 12314 14368
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 12710 14328 12716 14340
rect 4120 14300 12716 14328
rect 4120 14288 4126 14300
rect 12710 14288 12716 14300
rect 12768 14288 12774 14340
rect 13722 14288 13728 14340
rect 13780 14328 13786 14340
rect 15378 14328 15384 14340
rect 13780 14300 15384 14328
rect 13780 14288 13786 14300
rect 15378 14288 15384 14300
rect 15436 14288 15442 14340
rect 3050 14220 3056 14272
rect 3108 14260 3114 14272
rect 13446 14260 13452 14272
rect 3108 14232 13452 14260
rect 3108 14220 3114 14232
rect 13446 14220 13452 14232
rect 13504 14260 13510 14272
rect 13998 14260 14004 14272
rect 13504 14232 14004 14260
rect 13504 14220 13510 14232
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 15194 14220 15200 14272
rect 15252 14260 15258 14272
rect 15657 14263 15715 14269
rect 15657 14260 15669 14263
rect 15252 14232 15669 14260
rect 15252 14220 15258 14232
rect 15657 14229 15669 14232
rect 15703 14229 15715 14263
rect 15657 14223 15715 14229
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 1578 14016 1584 14068
rect 1636 14056 1642 14068
rect 2041 14059 2099 14065
rect 2041 14056 2053 14059
rect 1636 14028 2053 14056
rect 1636 14016 1642 14028
rect 2041 14025 2053 14028
rect 2087 14025 2099 14059
rect 2041 14019 2099 14025
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 3237 14059 3295 14065
rect 3237 14056 3249 14059
rect 2924 14028 3249 14056
rect 2924 14016 2930 14028
rect 3237 14025 3249 14028
rect 3283 14025 3295 14059
rect 3237 14019 3295 14025
rect 3694 14016 3700 14068
rect 3752 14056 3758 14068
rect 5718 14056 5724 14068
rect 3752 14028 5724 14056
rect 3752 14016 3758 14028
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 6181 14059 6239 14065
rect 6181 14025 6193 14059
rect 6227 14056 6239 14059
rect 6730 14056 6736 14068
rect 6227 14028 6736 14056
rect 6227 14025 6239 14028
rect 6181 14019 6239 14025
rect 6730 14016 6736 14028
rect 6788 14016 6794 14068
rect 13538 14016 13544 14068
rect 13596 14056 13602 14068
rect 14645 14059 14703 14065
rect 14645 14056 14657 14059
rect 13596 14028 14657 14056
rect 13596 14016 13602 14028
rect 14645 14025 14657 14028
rect 14691 14025 14703 14059
rect 14645 14019 14703 14025
rect 15562 14016 15568 14068
rect 15620 14056 15626 14068
rect 15841 14059 15899 14065
rect 15841 14056 15853 14059
rect 15620 14028 15853 14056
rect 15620 14016 15626 14028
rect 15841 14025 15853 14028
rect 15887 14025 15899 14059
rect 15841 14019 15899 14025
rect 5902 13948 5908 14000
rect 5960 13988 5966 14000
rect 7009 13991 7067 13997
rect 7009 13988 7021 13991
rect 5960 13960 7021 13988
rect 5960 13948 5966 13960
rect 7009 13957 7021 13960
rect 7055 13957 7067 13991
rect 7009 13951 7067 13957
rect 9398 13880 9404 13932
rect 9456 13920 9462 13932
rect 16206 13920 16212 13932
rect 9456 13892 16212 13920
rect 9456 13880 9462 13892
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13852 1915 13855
rect 2774 13852 2780 13864
rect 1903 13824 2780 13852
rect 1903 13821 1915 13824
rect 1857 13815 1915 13821
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 3050 13852 3056 13864
rect 3011 13824 3056 13852
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 5810 13812 5816 13864
rect 5868 13852 5874 13864
rect 5997 13855 6055 13861
rect 5997 13852 6009 13855
rect 5868 13824 6009 13852
rect 5868 13812 5874 13824
rect 5997 13821 6009 13824
rect 6043 13821 6055 13855
rect 5997 13815 6055 13821
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6144 13824 6837 13852
rect 6144 13812 6150 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 13633 13855 13691 13861
rect 13633 13821 13645 13855
rect 13679 13852 13691 13855
rect 14182 13852 14188 13864
rect 13679 13824 14188 13852
rect 13679 13821 13691 13824
rect 13633 13815 13691 13821
rect 14182 13812 14188 13824
rect 14240 13852 14246 13864
rect 14366 13852 14372 13864
rect 14240 13824 14372 13852
rect 14240 13812 14246 13824
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 14918 13852 14924 13864
rect 14507 13824 14924 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 14918 13812 14924 13824
rect 14976 13852 14982 13864
rect 15102 13852 15108 13864
rect 14976 13824 15108 13852
rect 14976 13812 14982 13824
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 15654 13852 15660 13864
rect 15615 13824 15660 13852
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 7374 13744 7380 13796
rect 7432 13784 7438 13796
rect 9214 13784 9220 13796
rect 7432 13756 9220 13784
rect 7432 13744 7438 13756
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 9306 13744 9312 13796
rect 9364 13784 9370 13796
rect 10226 13784 10232 13796
rect 9364 13756 10232 13784
rect 9364 13744 9370 13756
rect 10226 13744 10232 13756
rect 10284 13744 10290 13796
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 11974 13784 11980 13796
rect 11296 13756 11980 13784
rect 11296 13744 11302 13756
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 12084 13756 13860 13784
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 12084 13716 12112 13756
rect 13832 13725 13860 13756
rect 3568 13688 12112 13716
rect 13817 13719 13875 13725
rect 3568 13676 3574 13688
rect 13817 13685 13829 13719
rect 13863 13685 13875 13719
rect 13817 13679 13875 13685
rect 13998 13676 14004 13728
rect 14056 13716 14062 13728
rect 19610 13716 19616 13728
rect 14056 13688 19616 13716
rect 14056 13676 14062 13688
rect 19610 13676 19616 13688
rect 19668 13676 19674 13728
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 290 13472 296 13524
rect 348 13512 354 13524
rect 1765 13515 1823 13521
rect 1765 13512 1777 13515
rect 348 13484 1777 13512
rect 348 13472 354 13484
rect 1765 13481 1777 13484
rect 1811 13481 1823 13515
rect 1765 13475 1823 13481
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 13538 13512 13544 13524
rect 4304 13484 13544 13512
rect 4304 13472 4310 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 13630 13472 13636 13524
rect 13688 13512 13694 13524
rect 18322 13512 18328 13524
rect 13688 13484 18328 13512
rect 13688 13472 13694 13484
rect 18322 13472 18328 13484
rect 18380 13472 18386 13524
rect 1854 13404 1860 13456
rect 1912 13444 1918 13456
rect 2777 13447 2835 13453
rect 2777 13444 2789 13447
rect 1912 13416 2789 13444
rect 1912 13404 1918 13416
rect 2777 13413 2789 13416
rect 2823 13444 2835 13447
rect 3881 13447 3939 13453
rect 3881 13444 3893 13447
rect 2823 13416 3893 13444
rect 2823 13413 2835 13416
rect 2777 13407 2835 13413
rect 3881 13413 3893 13416
rect 3927 13413 3939 13447
rect 3881 13407 3939 13413
rect 5442 13404 5448 13456
rect 5500 13444 5506 13456
rect 15562 13444 15568 13456
rect 5500 13416 15568 13444
rect 5500 13404 5506 13416
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 1581 13379 1639 13385
rect 1581 13345 1593 13379
rect 1627 13345 1639 13379
rect 1581 13339 1639 13345
rect 2685 13379 2743 13385
rect 2685 13345 2697 13379
rect 2731 13376 2743 13379
rect 4065 13379 4123 13385
rect 4065 13376 4077 13379
rect 2731 13348 4077 13376
rect 2731 13345 2743 13348
rect 2685 13339 2743 13345
rect 4065 13345 4077 13348
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 1596 13308 1624 13339
rect 4798 13336 4804 13388
rect 4856 13376 4862 13388
rect 15194 13376 15200 13388
rect 4856 13348 15200 13376
rect 4856 13336 4862 13348
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 15448 13379 15506 13385
rect 15448 13345 15460 13379
rect 15494 13376 15506 13379
rect 16482 13376 16488 13388
rect 15494 13348 16488 13376
rect 15494 13345 15506 13348
rect 15448 13339 15506 13345
rect 16482 13336 16488 13348
rect 16540 13336 16546 13388
rect 17862 13376 17868 13388
rect 17823 13348 17868 13376
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 2958 13308 2964 13320
rect 1596 13280 2544 13308
rect 2919 13280 2964 13308
rect 1946 13132 1952 13184
rect 2004 13172 2010 13184
rect 2317 13175 2375 13181
rect 2317 13172 2329 13175
rect 2004 13144 2329 13172
rect 2004 13132 2010 13144
rect 2317 13141 2329 13144
rect 2363 13141 2375 13175
rect 2516 13172 2544 13280
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 9766 13308 9772 13320
rect 3620 13280 9772 13308
rect 3620 13172 3648 13280
rect 9766 13268 9772 13280
rect 9824 13308 9830 13320
rect 17034 13308 17040 13320
rect 9824 13280 17040 13308
rect 9824 13268 9830 13280
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 3881 13243 3939 13249
rect 3881 13209 3893 13243
rect 3927 13240 3939 13243
rect 7466 13240 7472 13252
rect 3927 13212 7472 13240
rect 3927 13209 3939 13212
rect 3881 13203 3939 13209
rect 7466 13200 7472 13212
rect 7524 13200 7530 13252
rect 15010 13200 15016 13252
rect 15068 13240 15074 13252
rect 18966 13240 18972 13252
rect 15068 13212 18972 13240
rect 15068 13200 15074 13212
rect 18966 13200 18972 13212
rect 19024 13200 19030 13252
rect 2516 13144 3648 13172
rect 2317 13135 2375 13141
rect 3694 13132 3700 13184
rect 3752 13172 3758 13184
rect 4706 13172 4712 13184
rect 3752 13144 4712 13172
rect 3752 13132 3758 13144
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 12710 13132 12716 13184
rect 12768 13172 12774 13184
rect 13170 13172 13176 13184
rect 12768 13144 13176 13172
rect 12768 13132 12774 13144
rect 13170 13132 13176 13144
rect 13228 13172 13234 13184
rect 15378 13172 15384 13184
rect 13228 13144 15384 13172
rect 13228 13132 13234 13144
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 15470 13132 15476 13184
rect 15528 13181 15534 13184
rect 15528 13175 15577 13181
rect 15528 13141 15531 13175
rect 15565 13141 15577 13175
rect 18046 13172 18052 13184
rect 18007 13144 18052 13172
rect 15528 13135 15577 13141
rect 15528 13132 15534 13135
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 4430 12968 4436 12980
rect 1627 12940 4436 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 4430 12928 4436 12940
rect 4488 12928 4494 12980
rect 15194 12900 15200 12912
rect 5920 12872 15200 12900
rect 2130 12832 2136 12844
rect 2091 12804 2136 12832
rect 2130 12792 2136 12804
rect 2188 12832 2194 12844
rect 2188 12804 2912 12832
rect 2188 12792 2194 12804
rect 1946 12764 1952 12776
rect 1907 12736 1952 12764
rect 1946 12724 1952 12736
rect 2004 12724 2010 12776
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12733 2835 12767
rect 2884 12764 2912 12804
rect 2884 12736 3832 12764
rect 2777 12727 2835 12733
rect 2792 12640 2820 12727
rect 2958 12656 2964 12708
rect 3016 12705 3022 12708
rect 3016 12699 3080 12705
rect 3016 12665 3034 12699
rect 3068 12665 3080 12699
rect 3016 12659 3080 12665
rect 3016 12656 3022 12659
rect 3804 12640 3832 12736
rect 4982 12724 4988 12776
rect 5040 12764 5046 12776
rect 5920 12773 5948 12872
rect 15194 12860 15200 12872
rect 15252 12860 15258 12912
rect 15378 12860 15384 12912
rect 15436 12900 15442 12912
rect 16669 12903 16727 12909
rect 15436 12872 15700 12900
rect 15436 12860 15442 12872
rect 6181 12835 6239 12841
rect 6181 12801 6193 12835
rect 6227 12832 6239 12835
rect 6638 12832 6644 12844
rect 6227 12804 6644 12832
rect 6227 12801 6239 12804
rect 6181 12795 6239 12801
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 11422 12792 11428 12844
rect 11480 12832 11486 12844
rect 15672 12832 15700 12872
rect 16669 12869 16681 12903
rect 16715 12900 16727 12903
rect 17954 12900 17960 12912
rect 16715 12872 17960 12900
rect 16715 12869 16727 12872
rect 16669 12863 16727 12869
rect 17954 12860 17960 12872
rect 18012 12860 18018 12912
rect 11480 12804 15608 12832
rect 15672 12804 17264 12832
rect 11480 12792 11486 12804
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 5040 12736 5457 12764
rect 5040 12724 5046 12736
rect 5445 12733 5457 12736
rect 5491 12764 5503 12767
rect 5905 12767 5963 12773
rect 5905 12764 5917 12767
rect 5491 12736 5917 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 5905 12733 5917 12736
rect 5951 12733 5963 12767
rect 5905 12727 5963 12733
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7892 12736 7941 12764
rect 7892 12724 7898 12736
rect 7929 12733 7941 12736
rect 7975 12764 7987 12767
rect 8018 12764 8024 12776
rect 7975 12736 8024 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 10870 12764 10876 12776
rect 8720 12736 10876 12764
rect 8720 12724 8726 12736
rect 10870 12724 10876 12736
rect 10928 12724 10934 12776
rect 12618 12724 12624 12776
rect 12676 12764 12682 12776
rect 12840 12767 12898 12773
rect 12840 12764 12852 12767
rect 12676 12736 12852 12764
rect 12676 12724 12682 12736
rect 12840 12733 12852 12736
rect 12886 12733 12898 12767
rect 12840 12727 12898 12733
rect 13998 12724 14004 12776
rect 14056 12764 14062 12776
rect 14220 12767 14278 12773
rect 14220 12764 14232 12767
rect 14056 12736 14232 12764
rect 14056 12724 14062 12736
rect 14220 12733 14232 12736
rect 14266 12733 14278 12767
rect 14220 12727 14278 12733
rect 14366 12724 14372 12776
rect 14424 12764 14430 12776
rect 15580 12773 15608 12804
rect 17236 12773 17264 12804
rect 14956 12767 15014 12773
rect 14956 12764 14968 12767
rect 14424 12736 14968 12764
rect 14424 12724 14430 12736
rect 14956 12733 14968 12736
rect 15002 12733 15014 12767
rect 14956 12727 15014 12733
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 16485 12767 16543 12773
rect 16485 12733 16497 12767
rect 16531 12733 16543 12767
rect 16485 12727 16543 12733
rect 17221 12767 17279 12773
rect 17221 12733 17233 12767
rect 17267 12733 17279 12767
rect 17221 12727 17279 12733
rect 8570 12696 8576 12708
rect 8531 12668 8576 12696
rect 8570 12656 8576 12668
rect 8628 12656 8634 12708
rect 8754 12656 8760 12708
rect 8812 12696 8818 12708
rect 13906 12696 13912 12708
rect 8812 12668 13912 12696
rect 8812 12656 8818 12668
rect 13906 12656 13912 12668
rect 13964 12656 13970 12708
rect 14734 12656 14740 12708
rect 14792 12696 14798 12708
rect 16500 12696 16528 12727
rect 14792 12668 16528 12696
rect 14792 12656 14798 12668
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 2774 12588 2780 12640
rect 2832 12588 2838 12640
rect 3786 12588 3792 12640
rect 3844 12628 3850 12640
rect 4157 12631 4215 12637
rect 4157 12628 4169 12631
rect 3844 12600 4169 12628
rect 3844 12588 3850 12600
rect 4157 12597 4169 12600
rect 4203 12597 4215 12631
rect 4614 12628 4620 12640
rect 4575 12600 4620 12628
rect 4157 12591 4215 12597
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 5534 12628 5540 12640
rect 5495 12600 5540 12628
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 5994 12628 6000 12640
rect 5955 12600 6000 12628
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 6825 12631 6883 12637
rect 6825 12597 6837 12631
rect 6871 12628 6883 12631
rect 7282 12628 7288 12640
rect 6871 12600 7288 12628
rect 6871 12597 6883 12600
rect 6825 12591 6883 12597
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 12943 12631 13001 12637
rect 12943 12597 12955 12631
rect 12989 12628 13001 12631
rect 13262 12628 13268 12640
rect 12989 12600 13268 12628
rect 12989 12597 13001 12600
rect 12943 12591 13001 12597
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 14323 12631 14381 12637
rect 14323 12597 14335 12631
rect 14369 12628 14381 12631
rect 14550 12628 14556 12640
rect 14369 12600 14556 12628
rect 14369 12597 14381 12600
rect 14323 12591 14381 12597
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 15010 12588 15016 12640
rect 15068 12637 15074 12640
rect 15068 12631 15117 12637
rect 15068 12597 15071 12631
rect 15105 12597 15117 12631
rect 15068 12591 15117 12597
rect 15749 12631 15807 12637
rect 15749 12597 15761 12631
rect 15795 12628 15807 12631
rect 16390 12628 16396 12640
rect 15795 12600 16396 12628
rect 15795 12597 15807 12600
rect 15749 12591 15807 12597
rect 15068 12588 15074 12591
rect 16390 12588 16396 12600
rect 16448 12588 16454 12640
rect 17402 12628 17408 12640
rect 17363 12600 17408 12628
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 2038 12384 2044 12436
rect 2096 12424 2102 12436
rect 2317 12427 2375 12433
rect 2317 12424 2329 12427
rect 2096 12396 2329 12424
rect 2096 12384 2102 12396
rect 2317 12393 2329 12396
rect 2363 12393 2375 12427
rect 2317 12387 2375 12393
rect 2590 12384 2596 12436
rect 2648 12424 2654 12436
rect 2685 12427 2743 12433
rect 2685 12424 2697 12427
rect 2648 12396 2697 12424
rect 2648 12384 2654 12396
rect 2685 12393 2697 12396
rect 2731 12424 2743 12427
rect 5626 12424 5632 12436
rect 2731 12396 5632 12424
rect 2731 12393 2743 12396
rect 2685 12387 2743 12393
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 9582 12424 9588 12436
rect 6196 12396 9588 12424
rect 6196 12368 6224 12396
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11112 12396 17172 12424
rect 11112 12384 11118 12396
rect 6178 12356 6184 12368
rect 1596 12328 6184 12356
rect 1596 12297 1624 12328
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 6638 12316 6644 12368
rect 6696 12365 6702 12368
rect 6696 12359 6760 12365
rect 6696 12325 6714 12359
rect 6748 12325 6760 12359
rect 6696 12319 6760 12325
rect 6696 12316 6702 12319
rect 6914 12316 6920 12368
rect 6972 12316 6978 12368
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 7524 12328 11192 12356
rect 7524 12316 7530 12328
rect 4890 12297 4896 12300
rect 1581 12291 1639 12297
rect 1581 12257 1593 12291
rect 1627 12257 1639 12291
rect 1581 12251 1639 12257
rect 4884 12251 4896 12297
rect 4948 12288 4954 12300
rect 6932 12288 6960 12316
rect 8662 12288 8668 12300
rect 4948 12260 4984 12288
rect 6472 12260 6960 12288
rect 8623 12260 8668 12288
rect 4890 12248 4896 12251
rect 4948 12248 4954 12260
rect 1670 12180 1676 12232
rect 1728 12220 1734 12232
rect 2777 12223 2835 12229
rect 2777 12220 2789 12223
rect 1728 12192 2789 12220
rect 1728 12180 1734 12192
rect 2777 12189 2789 12192
rect 2823 12189 2835 12223
rect 2958 12220 2964 12232
rect 2919 12192 2964 12220
rect 2777 12183 2835 12189
rect 2958 12180 2964 12192
rect 3016 12180 3022 12232
rect 4522 12180 4528 12232
rect 4580 12220 4586 12232
rect 6472 12229 6500 12260
rect 8662 12248 8668 12260
rect 8720 12248 8726 12300
rect 8754 12248 8760 12300
rect 8812 12288 8818 12300
rect 11164 12288 11192 12328
rect 11238 12316 11244 12368
rect 11296 12356 11302 12368
rect 11296 12328 14504 12356
rect 11296 12316 11302 12328
rect 11698 12288 11704 12300
rect 8812 12260 8857 12288
rect 11164 12260 11704 12288
rect 8812 12248 8818 12260
rect 11698 12248 11704 12260
rect 11756 12288 11762 12300
rect 12158 12288 12164 12300
rect 11756 12260 12164 12288
rect 11756 12248 11762 12260
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12472 12291 12530 12297
rect 12472 12288 12484 12291
rect 12268 12260 12484 12288
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 4580 12192 4629 12220
rect 4580 12180 4586 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 4617 12183 4675 12189
rect 5644 12192 6469 12220
rect 2498 12112 2504 12164
rect 2556 12152 2562 12164
rect 2976 12152 3004 12180
rect 2556 12124 3004 12152
rect 2556 12112 2562 12124
rect 1765 12087 1823 12093
rect 1765 12053 1777 12087
rect 1811 12084 1823 12087
rect 2866 12084 2872 12096
rect 1811 12056 2872 12084
rect 1811 12053 1823 12056
rect 1765 12047 1823 12053
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 4632 12084 4660 12183
rect 5644 12084 5672 12192
rect 6457 12189 6469 12192
rect 6503 12189 6515 12223
rect 6457 12183 6515 12189
rect 8941 12223 8999 12229
rect 8941 12189 8953 12223
rect 8987 12220 8999 12223
rect 9122 12220 9128 12232
rect 8987 12192 9128 12220
rect 8987 12189 8999 12192
rect 8941 12183 8999 12189
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 9582 12180 9588 12232
rect 9640 12180 9646 12232
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12268 12220 12296 12260
rect 12472 12257 12484 12260
rect 12518 12257 12530 12291
rect 12472 12251 12530 12257
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 14476 12297 14504 12328
rect 13392 12291 13450 12297
rect 13392 12288 13404 12291
rect 12768 12260 13404 12288
rect 12768 12248 12774 12260
rect 13392 12257 13404 12260
rect 13438 12257 13450 12291
rect 13392 12251 13450 12257
rect 14461 12291 14519 12297
rect 14461 12257 14473 12291
rect 14507 12257 14519 12291
rect 14461 12251 14519 12257
rect 15378 12248 15384 12300
rect 15436 12288 15442 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15436 12260 15669 12288
rect 15436 12248 15442 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 16393 12291 16451 12297
rect 16393 12257 16405 12291
rect 16439 12288 16451 12291
rect 16942 12288 16948 12300
rect 16439 12260 16948 12288
rect 16439 12257 16451 12260
rect 16393 12251 16451 12257
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17144 12297 17172 12396
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12257 17187 12291
rect 17865 12291 17923 12297
rect 17865 12288 17877 12291
rect 17129 12251 17187 12257
rect 17236 12260 17877 12288
rect 12124 12192 12296 12220
rect 12124 12180 12130 12192
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 17236 12220 17264 12260
rect 17865 12257 17877 12260
rect 17911 12257 17923 12291
rect 17865 12251 17923 12257
rect 13872 12192 17264 12220
rect 13872 12180 13878 12192
rect 9600 12152 9628 12180
rect 12342 12152 12348 12164
rect 9600 12124 12348 12152
rect 12342 12112 12348 12124
rect 12400 12112 12406 12164
rect 16577 12155 16635 12161
rect 16577 12121 16589 12155
rect 16623 12152 16635 12155
rect 19150 12152 19156 12164
rect 16623 12124 19156 12152
rect 16623 12121 16635 12124
rect 16577 12115 16635 12121
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 4632 12056 5672 12084
rect 5997 12087 6055 12093
rect 5997 12053 6009 12087
rect 6043 12084 6055 12087
rect 6454 12084 6460 12096
rect 6043 12056 6460 12084
rect 6043 12053 6055 12056
rect 5997 12047 6055 12053
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 7650 12084 7656 12096
rect 6788 12056 7656 12084
rect 6788 12044 6794 12056
rect 7650 12044 7656 12056
rect 7708 12084 7714 12096
rect 7837 12087 7895 12093
rect 7837 12084 7849 12087
rect 7708 12056 7849 12084
rect 7708 12044 7714 12056
rect 7837 12053 7849 12056
rect 7883 12053 7895 12087
rect 7837 12047 7895 12053
rect 8297 12087 8355 12093
rect 8297 12053 8309 12087
rect 8343 12084 8355 12087
rect 8386 12084 8392 12096
rect 8343 12056 8392 12084
rect 8343 12053 8355 12056
rect 8297 12047 8355 12053
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 12526 12044 12532 12096
rect 12584 12093 12590 12096
rect 12584 12087 12633 12093
rect 12584 12053 12587 12087
rect 12621 12053 12633 12087
rect 12584 12047 12633 12053
rect 12584 12044 12590 12047
rect 13446 12044 13452 12096
rect 13504 12093 13510 12096
rect 13504 12087 13553 12093
rect 13504 12053 13507 12087
rect 13541 12053 13553 12087
rect 13504 12047 13553 12053
rect 14645 12087 14703 12093
rect 14645 12053 14657 12087
rect 14691 12084 14703 12087
rect 14826 12084 14832 12096
rect 14691 12056 14832 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 13504 12044 13510 12047
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 15841 12087 15899 12093
rect 15841 12053 15853 12087
rect 15887 12084 15899 12087
rect 16114 12084 16120 12096
rect 15887 12056 16120 12084
rect 15887 12053 15899 12056
rect 15841 12047 15899 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 17313 12087 17371 12093
rect 17313 12053 17325 12087
rect 17359 12084 17371 12087
rect 17494 12084 17500 12096
rect 17359 12056 17500 12084
rect 17359 12053 17371 12056
rect 17313 12047 17371 12053
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 18049 12087 18107 12093
rect 18049 12053 18061 12087
rect 18095 12084 18107 12087
rect 18230 12084 18236 12096
rect 18095 12056 18236 12084
rect 18095 12053 18107 12056
rect 18049 12047 18107 12053
rect 18230 12044 18236 12056
rect 18288 12044 18294 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 4522 11880 4528 11892
rect 3620 11852 4528 11880
rect 2774 11772 2780 11824
rect 2832 11812 2838 11824
rect 3620 11812 3648 11852
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 4890 11840 4896 11892
rect 4948 11880 4954 11892
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4948 11852 4997 11880
rect 4948 11840 4954 11852
rect 4985 11849 4997 11852
rect 5031 11849 5043 11883
rect 4985 11843 5043 11849
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 11054 11880 11060 11892
rect 9640 11852 11060 11880
rect 9640 11840 9646 11852
rect 11054 11840 11060 11852
rect 11112 11840 11118 11892
rect 11606 11840 11612 11892
rect 11664 11880 11670 11892
rect 15197 11883 15255 11889
rect 11664 11852 14228 11880
rect 11664 11840 11670 11852
rect 2832 11784 3648 11812
rect 2832 11772 2838 11784
rect 2498 11704 2504 11756
rect 2556 11744 2562 11756
rect 3620 11753 3648 11784
rect 7834 11772 7840 11824
rect 7892 11812 7898 11824
rect 8665 11815 8723 11821
rect 8665 11812 8677 11815
rect 7892 11784 8677 11812
rect 7892 11772 7898 11784
rect 8665 11781 8677 11784
rect 8711 11781 8723 11815
rect 8665 11775 8723 11781
rect 2869 11747 2927 11753
rect 2869 11744 2881 11747
rect 2556 11716 2881 11744
rect 2556 11704 2562 11716
rect 2869 11713 2881 11716
rect 2915 11713 2927 11747
rect 2869 11707 2927 11713
rect 3605 11747 3663 11753
rect 3605 11713 3617 11747
rect 3651 11713 3663 11747
rect 3605 11707 3663 11713
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 5905 11747 5963 11753
rect 5905 11744 5917 11747
rect 5592 11716 5917 11744
rect 5592 11704 5598 11716
rect 5905 11713 5917 11716
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 6089 11747 6147 11753
rect 6089 11713 6101 11747
rect 6135 11744 6147 11747
rect 6730 11744 6736 11756
rect 6135 11716 6736 11744
rect 6135 11713 6147 11716
rect 6089 11707 6147 11713
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9217 11747 9275 11753
rect 9217 11744 9229 11747
rect 9180 11716 9229 11744
rect 9180 11704 9186 11716
rect 9217 11713 9229 11716
rect 9263 11713 9275 11747
rect 9217 11707 9275 11713
rect 12342 11704 12348 11756
rect 12400 11744 12406 11756
rect 13081 11747 13139 11753
rect 13081 11744 13093 11747
rect 12400 11716 13093 11744
rect 12400 11704 12406 11716
rect 13081 11713 13093 11716
rect 13127 11744 13139 11747
rect 13630 11744 13636 11756
rect 13127 11716 13636 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 14200 11753 14228 11852
rect 15197 11849 15209 11883
rect 15243 11880 15255 11883
rect 17586 11880 17592 11892
rect 15243 11852 17592 11880
rect 15243 11849 15255 11852
rect 15197 11843 15255 11849
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 16206 11772 16212 11824
rect 16264 11812 16270 11824
rect 19610 11812 19616 11824
rect 16264 11784 19616 11812
rect 16264 11772 16270 11784
rect 19610 11772 19616 11784
rect 19668 11772 19674 11824
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11713 14243 11747
rect 15930 11744 15936 11756
rect 14185 11707 14243 11713
rect 14936 11716 15936 11744
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11676 1639 11679
rect 1854 11676 1860 11688
rect 1627 11648 1860 11676
rect 1627 11645 1639 11648
rect 1581 11639 1639 11645
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 2682 11676 2688 11688
rect 2595 11648 2688 11676
rect 2682 11636 2688 11648
rect 2740 11676 2746 11688
rect 6362 11676 6368 11688
rect 2740 11648 6368 11676
rect 2740 11636 2746 11648
rect 6362 11636 6368 11648
rect 6420 11636 6426 11688
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 6914 11676 6920 11688
rect 6871 11648 6920 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 6914 11636 6920 11648
rect 6972 11676 6978 11688
rect 7466 11676 7472 11688
rect 6972 11648 7472 11676
rect 6972 11636 6978 11648
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 7558 11636 7564 11688
rect 7616 11676 7622 11688
rect 12158 11676 12164 11688
rect 7616 11648 12164 11676
rect 7616 11636 7622 11648
rect 12158 11636 12164 11648
rect 12216 11676 12222 11688
rect 14936 11676 14964 11716
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 17126 11744 17132 11756
rect 16316 11716 17132 11744
rect 12216 11648 14964 11676
rect 15013 11679 15071 11685
rect 12216 11636 12222 11648
rect 15013 11645 15025 11679
rect 15059 11676 15071 11679
rect 15102 11676 15108 11688
rect 15059 11648 15108 11676
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 15749 11679 15807 11685
rect 15749 11645 15761 11679
rect 15795 11676 15807 11679
rect 16316 11676 16344 11716
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 17862 11704 17868 11756
rect 17920 11744 17926 11756
rect 18322 11744 18328 11756
rect 17920 11716 18328 11744
rect 17920 11704 17926 11716
rect 18322 11704 18328 11716
rect 18380 11704 18386 11756
rect 16482 11676 16488 11688
rect 15795 11648 16344 11676
rect 16443 11648 16488 11676
rect 15795 11645 15807 11648
rect 15749 11639 15807 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 3786 11568 3792 11620
rect 3844 11617 3850 11620
rect 3844 11611 3908 11617
rect 3844 11577 3862 11611
rect 3896 11577 3908 11611
rect 3844 11571 3908 11577
rect 3844 11568 3850 11571
rect 6730 11568 6736 11620
rect 6788 11608 6794 11620
rect 7070 11611 7128 11617
rect 7070 11608 7082 11611
rect 6788 11580 7082 11608
rect 6788 11568 6794 11580
rect 7070 11577 7082 11580
rect 7116 11577 7128 11611
rect 12805 11611 12863 11617
rect 12805 11608 12817 11611
rect 7070 11571 7128 11577
rect 7208 11580 12817 11608
rect 1762 11540 1768 11552
rect 1723 11512 1768 11540
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 2317 11543 2375 11549
rect 2317 11540 2329 11543
rect 1912 11512 2329 11540
rect 1912 11500 1918 11512
rect 2317 11509 2329 11512
rect 2363 11509 2375 11543
rect 2317 11503 2375 11509
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 5442 11540 5448 11552
rect 2832 11512 2877 11540
rect 5403 11512 5448 11540
rect 2832 11500 2838 11512
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 5776 11512 5825 11540
rect 5776 11500 5782 11512
rect 5813 11509 5825 11512
rect 5859 11540 5871 11543
rect 5994 11540 6000 11552
rect 5859 11512 6000 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 7208 11540 7236 11580
rect 12805 11577 12817 11580
rect 12851 11608 12863 11611
rect 13538 11608 13544 11620
rect 12851 11580 13544 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 13538 11568 13544 11580
rect 13596 11568 13602 11620
rect 14001 11611 14059 11617
rect 14001 11577 14013 11611
rect 14047 11608 14059 11611
rect 14458 11608 14464 11620
rect 14047 11580 14464 11608
rect 14047 11577 14059 11580
rect 14001 11571 14059 11577
rect 14458 11568 14464 11580
rect 14516 11568 14522 11620
rect 14642 11568 14648 11620
rect 14700 11608 14706 11620
rect 17236 11608 17264 11639
rect 14700 11580 16344 11608
rect 14700 11568 14706 11580
rect 8202 11540 8208 11552
rect 6420 11512 7236 11540
rect 8163 11512 8208 11540
rect 6420 11500 6426 11512
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 9030 11540 9036 11552
rect 8991 11512 9036 11540
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9122 11500 9128 11552
rect 9180 11540 9186 11552
rect 9180 11512 9225 11540
rect 9180 11500 9186 11512
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12897 11543 12955 11549
rect 12492 11512 12537 11540
rect 12492 11500 12498 11512
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 13354 11540 13360 11552
rect 12943 11512 13360 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 14090 11500 14096 11552
rect 14148 11540 14154 11552
rect 14148 11512 14193 11540
rect 14148 11500 14154 11512
rect 14274 11500 14280 11552
rect 14332 11540 14338 11552
rect 15102 11540 15108 11552
rect 14332 11512 15108 11540
rect 14332 11500 14338 11512
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15933 11543 15991 11549
rect 15933 11509 15945 11543
rect 15979 11540 15991 11543
rect 16206 11540 16212 11552
rect 15979 11512 16212 11540
rect 15979 11509 15991 11512
rect 15933 11503 15991 11509
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16316 11540 16344 11580
rect 16500 11580 17264 11608
rect 16500 11540 16528 11580
rect 16316 11512 16528 11540
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 16669 11543 16727 11549
rect 16669 11540 16681 11543
rect 16632 11512 16681 11540
rect 16632 11500 16638 11512
rect 16669 11509 16681 11512
rect 16715 11509 16727 11543
rect 17402 11540 17408 11552
rect 17363 11512 17408 11540
rect 16669 11503 16727 11509
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 2685 11339 2743 11345
rect 2685 11305 2697 11339
rect 2731 11336 2743 11339
rect 2774 11336 2780 11348
rect 2731 11308 2780 11336
rect 2731 11305 2743 11308
rect 2685 11299 2743 11305
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 2958 11296 2964 11348
rect 3016 11336 3022 11348
rect 3145 11339 3203 11345
rect 3145 11336 3157 11339
rect 3016 11308 3157 11336
rect 3016 11296 3022 11308
rect 3145 11305 3157 11308
rect 3191 11305 3203 11339
rect 3145 11299 3203 11305
rect 3234 11296 3240 11348
rect 3292 11336 3298 11348
rect 3418 11336 3424 11348
rect 3292 11308 3424 11336
rect 3292 11296 3298 11308
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 3510 11296 3516 11348
rect 3568 11336 3574 11348
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 3568 11308 4077 11336
rect 3568 11296 3574 11308
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 4430 11336 4436 11348
rect 4391 11308 4436 11336
rect 4065 11299 4123 11305
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 6086 11296 6092 11348
rect 6144 11336 6150 11348
rect 6362 11336 6368 11348
rect 6144 11308 6368 11336
rect 6144 11296 6150 11308
rect 6362 11296 6368 11308
rect 6420 11336 6426 11348
rect 14642 11336 14648 11348
rect 6420 11308 14648 11336
rect 6420 11296 6426 11308
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 15194 11296 15200 11348
rect 15252 11336 15258 11348
rect 15562 11336 15568 11348
rect 15252 11308 15568 11336
rect 15252 11296 15258 11308
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 15657 11339 15715 11345
rect 15657 11305 15669 11339
rect 15703 11336 15715 11339
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 15703 11308 16497 11336
rect 15703 11305 15715 11308
rect 15657 11299 15715 11305
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 16485 11299 16543 11305
rect 2976 11200 3004 11296
rect 3053 11271 3111 11277
rect 3053 11237 3065 11271
rect 3099 11268 3111 11271
rect 5350 11268 5356 11280
rect 3099 11240 5356 11268
rect 3099 11237 3111 11240
rect 3053 11231 3111 11237
rect 5350 11228 5356 11240
rect 5408 11228 5414 11280
rect 6270 11228 6276 11280
rect 6328 11268 6334 11280
rect 7736 11271 7794 11277
rect 7736 11268 7748 11271
rect 6328 11240 6776 11268
rect 6328 11228 6334 11240
rect 5626 11200 5632 11212
rect 2976 11172 5632 11200
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5721 11203 5779 11209
rect 5721 11169 5733 11203
rect 5767 11200 5779 11203
rect 6638 11200 6644 11212
rect 5767 11172 6644 11200
rect 5767 11169 5779 11172
rect 5721 11163 5779 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 6748 11209 6776 11240
rect 6840 11240 7748 11268
rect 6733 11203 6791 11209
rect 6733 11169 6745 11203
rect 6779 11169 6791 11203
rect 6733 11163 6791 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 1949 11135 2007 11141
rect 1949 11132 1961 11135
rect 1636 11104 1961 11132
rect 1636 11092 1642 11104
rect 1949 11101 1961 11104
rect 1995 11101 2007 11135
rect 2130 11132 2136 11144
rect 2091 11104 2136 11132
rect 1949 11095 2007 11101
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 3326 11132 3332 11144
rect 3287 11104 3332 11132
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 4890 11132 4896 11144
rect 4755 11104 4896 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 1489 11067 1547 11073
rect 1489 11033 1501 11067
rect 1535 11064 1547 11067
rect 4540 11064 4568 11095
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 5810 11132 5816 11144
rect 5771 11104 5816 11132
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 5994 11132 6000 11144
rect 5907 11104 6000 11132
rect 5994 11092 6000 11104
rect 6052 11132 6058 11144
rect 6840 11132 6868 11240
rect 7736 11237 7748 11240
rect 7782 11268 7794 11271
rect 8202 11268 8208 11280
rect 7782 11240 8208 11268
rect 7782 11237 7794 11240
rect 7736 11231 7794 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 13078 11268 13084 11280
rect 10520 11240 13084 11268
rect 7466 11132 7472 11144
rect 6052 11104 6868 11132
rect 7427 11104 7472 11132
rect 6052 11092 6058 11104
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 8754 11092 8760 11144
rect 8812 11132 8818 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 8812 11104 9689 11132
rect 8812 11092 8818 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 10318 11092 10324 11144
rect 10376 11132 10382 11144
rect 10520 11141 10548 11240
rect 10772 11203 10830 11209
rect 10772 11169 10784 11203
rect 10818 11200 10830 11203
rect 11330 11200 11336 11212
rect 10818 11172 11336 11200
rect 10818 11169 10830 11172
rect 10772 11163 10830 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 12544 11209 12572 11240
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 13538 11228 13544 11280
rect 13596 11268 13602 11280
rect 13596 11240 17908 11268
rect 13596 11228 13602 11240
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11169 12587 11203
rect 12529 11163 12587 11169
rect 12796 11203 12854 11209
rect 12796 11169 12808 11203
rect 12842 11200 12854 11203
rect 12842 11172 13584 11200
rect 12842 11169 12854 11172
rect 12796 11163 12854 11169
rect 13556 11144 13584 11172
rect 14366 11160 14372 11212
rect 14424 11200 14430 11212
rect 14461 11203 14519 11209
rect 14461 11200 14473 11203
rect 14424 11172 14473 11200
rect 14424 11160 14430 11172
rect 14461 11169 14473 11172
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 15194 11160 15200 11212
rect 15252 11160 15258 11212
rect 16850 11200 16856 11212
rect 16811 11172 16856 11200
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 17880 11209 17908 11240
rect 17865 11203 17923 11209
rect 17865 11169 17877 11203
rect 17911 11169 17923 11203
rect 17865 11163 17923 11169
rect 10505 11135 10563 11141
rect 10505 11132 10517 11135
rect 10376 11104 10517 11132
rect 10376 11092 10382 11104
rect 10505 11101 10517 11104
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 13538 11092 13544 11144
rect 13596 11092 13602 11144
rect 13722 11092 13728 11144
rect 13780 11092 13786 11144
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 15212 11132 15240 11160
rect 13964 11104 15240 11132
rect 13964 11092 13970 11104
rect 15654 11092 15660 11144
rect 15712 11132 15718 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15712 11104 15761 11132
rect 15712 11092 15718 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 1535 11036 4568 11064
rect 5184 11036 5488 11064
rect 1535 11033 1547 11036
rect 1489 11027 1547 11033
rect 1670 10956 1676 11008
rect 1728 10996 1734 11008
rect 5184 10996 5212 11036
rect 5350 10996 5356 11008
rect 1728 10968 5212 10996
rect 5311 10968 5356 10996
rect 1728 10956 1734 10968
rect 5350 10956 5356 10968
rect 5408 10956 5414 11008
rect 5460 10996 5488 11036
rect 6546 11024 6552 11076
rect 6604 11064 6610 11076
rect 6917 11067 6975 11073
rect 6917 11064 6929 11067
rect 6604 11036 6929 11064
rect 6604 11024 6610 11036
rect 6917 11033 6929 11036
rect 6963 11033 6975 11067
rect 13740 11064 13768 11092
rect 6917 11027 6975 11033
rect 8680 11036 8984 11064
rect 13740 11036 13952 11064
rect 8680 10996 8708 11036
rect 8846 10996 8852 11008
rect 5460 10968 8708 10996
rect 8807 10968 8852 10996
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 8956 10996 8984 11036
rect 10410 10996 10416 11008
rect 8956 10968 10416 10996
rect 10410 10956 10416 10968
rect 10468 10956 10474 11008
rect 11790 10956 11796 11008
rect 11848 10996 11854 11008
rect 13924 11005 13952 11036
rect 15562 11024 15568 11076
rect 15620 11064 15626 11076
rect 15856 11064 15884 11095
rect 16206 11092 16212 11144
rect 16264 11132 16270 11144
rect 16390 11132 16396 11144
rect 16264 11104 16396 11132
rect 16264 11092 16270 11104
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 16758 11092 16764 11144
rect 16816 11132 16822 11144
rect 16945 11135 17003 11141
rect 16945 11132 16957 11135
rect 16816 11104 16957 11132
rect 16816 11092 16822 11104
rect 16945 11101 16957 11104
rect 16991 11101 17003 11135
rect 16945 11095 17003 11101
rect 17034 11092 17040 11144
rect 17092 11132 17098 11144
rect 17092 11104 17137 11132
rect 17092 11092 17098 11104
rect 15620 11036 15884 11064
rect 18049 11067 18107 11073
rect 15620 11024 15626 11036
rect 18049 11033 18061 11067
rect 18095 11064 18107 11067
rect 18138 11064 18144 11076
rect 18095 11036 18144 11064
rect 18095 11033 18107 11036
rect 18049 11027 18107 11033
rect 18138 11024 18144 11036
rect 18196 11024 18202 11076
rect 11885 10999 11943 11005
rect 11885 10996 11897 10999
rect 11848 10968 11897 10996
rect 11848 10956 11854 10968
rect 11885 10965 11897 10968
rect 11931 10965 11943 10999
rect 11885 10959 11943 10965
rect 13909 10999 13967 11005
rect 13909 10965 13921 10999
rect 13955 10965 13967 10999
rect 14642 10996 14648 11008
rect 14603 10968 14648 10996
rect 13909 10959 13967 10965
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 15102 10956 15108 11008
rect 15160 10996 15166 11008
rect 15289 10999 15347 11005
rect 15289 10996 15301 10999
rect 15160 10968 15301 10996
rect 15160 10956 15166 10968
rect 15289 10965 15301 10968
rect 15335 10965 15347 10999
rect 15289 10959 15347 10965
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 12250 10792 12256 10804
rect 1688 10764 12256 10792
rect 1688 10597 1716 10764
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 12986 10792 12992 10804
rect 12947 10764 12992 10792
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 13722 10792 13728 10804
rect 13556 10764 13728 10792
rect 3789 10727 3847 10733
rect 3789 10693 3801 10727
rect 3835 10693 3847 10727
rect 3789 10687 3847 10693
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10557 1731 10591
rect 2406 10588 2412 10600
rect 2367 10560 2412 10588
rect 1673 10551 1731 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 3804 10588 3832 10687
rect 4246 10684 4252 10736
rect 4304 10724 4310 10736
rect 4341 10727 4399 10733
rect 4341 10724 4353 10727
rect 4304 10696 4353 10724
rect 4304 10684 4310 10696
rect 4341 10693 4353 10696
rect 4387 10724 4399 10727
rect 4522 10724 4528 10736
rect 4387 10696 4528 10724
rect 4387 10693 4399 10696
rect 4341 10687 4399 10693
rect 4522 10684 4528 10696
rect 4580 10684 4586 10736
rect 5534 10724 5540 10736
rect 5184 10696 5540 10724
rect 5184 10656 5212 10696
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 6638 10684 6644 10736
rect 6696 10724 6702 10736
rect 6825 10727 6883 10733
rect 6825 10724 6837 10727
rect 6696 10696 6837 10724
rect 6696 10684 6702 10696
rect 6825 10693 6837 10696
rect 6871 10693 6883 10727
rect 8846 10724 8852 10736
rect 6825 10687 6883 10693
rect 7300 10696 8852 10724
rect 2556 10560 3832 10588
rect 4448 10628 5212 10656
rect 5261 10659 5319 10665
rect 2556 10548 2562 10560
rect 2676 10523 2734 10529
rect 2676 10489 2688 10523
rect 2722 10520 2734 10523
rect 3326 10520 3332 10532
rect 2722 10492 3332 10520
rect 2722 10489 2734 10492
rect 2676 10483 2734 10489
rect 3326 10480 3332 10492
rect 3384 10480 3390 10532
rect 1857 10455 1915 10461
rect 1857 10421 1869 10455
rect 1903 10452 1915 10455
rect 2774 10452 2780 10464
rect 1903 10424 2780 10452
rect 1903 10421 1915 10424
rect 1857 10415 1915 10421
rect 2774 10412 2780 10424
rect 2832 10412 2838 10464
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 4448 10452 4476 10628
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 7300 10656 7328 10696
rect 8846 10684 8852 10696
rect 8904 10684 8910 10736
rect 5307 10628 7328 10656
rect 7469 10659 7527 10665
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7650 10656 7656 10668
rect 7515 10628 7656 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 10410 10616 10416 10668
rect 10468 10656 10474 10668
rect 11146 10656 11152 10668
rect 10468 10628 11152 10656
rect 10468 10616 10474 10628
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 11388 10628 11652 10656
rect 11388 10616 11394 10628
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10557 4583 10591
rect 4525 10551 4583 10557
rect 4985 10591 5043 10597
rect 4985 10557 4997 10591
rect 5031 10588 5043 10591
rect 5350 10588 5356 10600
rect 5031 10560 5356 10588
rect 5031 10557 5043 10560
rect 4985 10551 5043 10557
rect 4540 10520 4568 10551
rect 5350 10548 5356 10560
rect 5408 10548 5414 10600
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10588 5871 10591
rect 6730 10588 6736 10600
rect 5859 10560 6736 10588
rect 5859 10557 5871 10560
rect 5813 10551 5871 10557
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10588 7251 10591
rect 7282 10588 7288 10600
rect 7239 10560 7288 10588
rect 7239 10557 7251 10560
rect 7193 10551 7251 10557
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 7926 10548 7932 10600
rect 7984 10588 7990 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 7984 10560 8033 10588
rect 7984 10548 7990 10560
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10588 8907 10591
rect 10318 10588 10324 10600
rect 8895 10560 10324 10588
rect 8895 10557 8907 10560
rect 8849 10551 8907 10557
rect 10318 10548 10324 10560
rect 10376 10588 10382 10600
rect 10778 10588 10784 10600
rect 10376 10560 10784 10588
rect 10376 10548 10382 10560
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 11054 10588 11060 10600
rect 11015 10560 11060 10588
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 5258 10520 5264 10532
rect 4540 10492 5264 10520
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 6089 10523 6147 10529
rect 6089 10489 6101 10523
rect 6135 10489 6147 10523
rect 6089 10483 6147 10489
rect 9116 10523 9174 10529
rect 9116 10489 9128 10523
rect 9162 10520 9174 10523
rect 11624 10520 11652 10628
rect 13078 10616 13084 10668
rect 13136 10656 13142 10668
rect 13556 10665 13584 10764
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 13136 10628 13553 10656
rect 13136 10616 13142 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 12250 10548 12256 10600
rect 12308 10588 12314 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12308 10560 12817 10588
rect 12308 10548 12314 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 13556 10588 13584 10619
rect 15381 10591 15439 10597
rect 15381 10588 15393 10591
rect 13556 10560 15393 10588
rect 12805 10551 12863 10557
rect 15381 10557 15393 10560
rect 15427 10557 15439 10591
rect 15381 10551 15439 10557
rect 16022 10548 16028 10600
rect 16080 10588 16086 10600
rect 16482 10588 16488 10600
rect 16080 10560 16488 10588
rect 16080 10548 16086 10560
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 17218 10588 17224 10600
rect 17179 10560 17224 10588
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 12342 10520 12348 10532
rect 9162 10492 11560 10520
rect 11624 10492 12348 10520
rect 9162 10489 9174 10492
rect 9116 10483 9174 10489
rect 3108 10424 4476 10452
rect 3108 10412 3114 10424
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 4617 10455 4675 10461
rect 4617 10452 4629 10455
rect 4580 10424 4629 10452
rect 4580 10412 4586 10424
rect 4617 10421 4629 10424
rect 4663 10421 4675 10455
rect 4617 10415 4675 10421
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 5132 10424 5177 10452
rect 5132 10412 5138 10424
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 6104 10452 6132 10483
rect 5408 10424 6132 10452
rect 5408 10412 5414 10424
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 6236 10424 7297 10452
rect 6236 10412 6242 10424
rect 7285 10421 7297 10424
rect 7331 10421 7343 10455
rect 7285 10415 7343 10421
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 7524 10424 8217 10452
rect 7524 10412 7530 10424
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8205 10415 8263 10421
rect 9490 10412 9496 10464
rect 9548 10452 9554 10464
rect 10134 10452 10140 10464
rect 9548 10424 10140 10452
rect 9548 10412 9554 10424
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 10229 10455 10287 10461
rect 10229 10421 10241 10455
rect 10275 10452 10287 10455
rect 10318 10452 10324 10464
rect 10275 10424 10324 10452
rect 10275 10421 10287 10424
rect 10229 10415 10287 10421
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 10686 10452 10692 10464
rect 10647 10424 10692 10452
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 11532 10452 11560 10492
rect 12342 10480 12348 10492
rect 12400 10480 12406 10532
rect 13808 10523 13866 10529
rect 13808 10489 13820 10523
rect 13854 10520 13866 10523
rect 15470 10520 15476 10532
rect 13854 10492 15476 10520
rect 13854 10489 13866 10492
rect 13808 10483 13866 10489
rect 15470 10480 15476 10492
rect 15528 10480 15534 10532
rect 15648 10523 15706 10529
rect 15648 10489 15660 10523
rect 15694 10489 15706 10523
rect 16666 10520 16672 10532
rect 15648 10483 15706 10489
rect 16408 10492 16672 10520
rect 11790 10452 11796 10464
rect 11532 10424 11796 10452
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 13596 10424 14933 10452
rect 13596 10412 13602 10424
rect 14921 10421 14933 10424
rect 14967 10421 14979 10455
rect 15663 10452 15691 10483
rect 16408 10452 16436 10492
rect 16666 10480 16672 10492
rect 16724 10480 16730 10532
rect 15663 10424 16436 10452
rect 14921 10415 14979 10421
rect 16482 10412 16488 10464
rect 16540 10452 16546 10464
rect 16761 10455 16819 10461
rect 16761 10452 16773 10455
rect 16540 10424 16773 10452
rect 16540 10412 16546 10424
rect 16761 10421 16773 10424
rect 16807 10452 16819 10455
rect 17034 10452 17040 10464
rect 16807 10424 17040 10452
rect 16807 10421 16819 10424
rect 16761 10415 16819 10421
rect 17034 10412 17040 10424
rect 17092 10412 17098 10464
rect 17310 10412 17316 10464
rect 17368 10452 17374 10464
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 17368 10424 17417 10452
rect 17368 10412 17374 10424
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 1995 10220 2789 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 2777 10211 2835 10217
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 3145 10251 3203 10257
rect 3145 10248 3157 10251
rect 3108 10220 3157 10248
rect 3108 10208 3114 10220
rect 3145 10217 3157 10220
rect 3191 10217 3203 10251
rect 3145 10211 3203 10217
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 4890 10248 4896 10260
rect 3752 10220 4896 10248
rect 3752 10208 3758 10220
rect 4890 10208 4896 10220
rect 4948 10208 4954 10260
rect 4985 10251 5043 10257
rect 4985 10217 4997 10251
rect 5031 10248 5043 10251
rect 5074 10248 5080 10260
rect 5031 10220 5080 10248
rect 5031 10217 5043 10220
rect 4985 10211 5043 10217
rect 5074 10208 5080 10220
rect 5132 10208 5138 10260
rect 5353 10251 5411 10257
rect 5353 10217 5365 10251
rect 5399 10248 5411 10251
rect 5442 10248 5448 10260
rect 5399 10220 5448 10248
rect 5399 10217 5411 10220
rect 5353 10211 5411 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 5868 10220 6193 10248
rect 5868 10208 5874 10220
rect 6181 10217 6193 10220
rect 6227 10217 6239 10251
rect 6181 10211 6239 10217
rect 6362 10208 6368 10260
rect 6420 10248 6426 10260
rect 6549 10251 6607 10257
rect 6549 10248 6561 10251
rect 6420 10220 6561 10248
rect 6420 10208 6426 10220
rect 6549 10217 6561 10220
rect 6595 10217 6607 10251
rect 6549 10211 6607 10217
rect 6730 10208 6736 10260
rect 6788 10248 6794 10260
rect 9769 10251 9827 10257
rect 9769 10248 9781 10251
rect 6788 10220 8432 10248
rect 6788 10208 6794 10220
rect 3786 10140 3792 10192
rect 3844 10180 3850 10192
rect 4341 10183 4399 10189
rect 4341 10180 4353 10183
rect 3844 10152 4353 10180
rect 3844 10140 3850 10152
rect 4341 10149 4353 10152
rect 4387 10149 4399 10183
rect 4341 10143 4399 10149
rect 5626 10140 5632 10192
rect 5684 10180 5690 10192
rect 6641 10183 6699 10189
rect 6641 10180 6653 10183
rect 5684 10152 6653 10180
rect 5684 10140 5690 10152
rect 6641 10149 6653 10152
rect 6687 10180 6699 10183
rect 7828 10183 7886 10189
rect 6687 10152 7779 10180
rect 6687 10149 6699 10152
rect 6641 10143 6699 10149
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 3050 10112 3056 10124
rect 2087 10084 3056 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 3988 10084 4077 10112
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2498 10044 2504 10056
rect 2271 10016 2504 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 2958 10004 2964 10056
rect 3016 10044 3022 10056
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 3016 10016 3249 10044
rect 3016 10004 3022 10016
rect 3237 10013 3249 10016
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3326 10004 3332 10056
rect 3384 10044 3390 10056
rect 3384 10016 3429 10044
rect 3384 10004 3390 10016
rect 3988 9908 4016 10084
rect 4065 10081 4077 10084
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 5810 10112 5816 10124
rect 4212 10084 5816 10112
rect 4212 10072 4218 10084
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 7558 10112 7564 10124
rect 7519 10084 7564 10112
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 7650 10072 7656 10124
rect 7708 10072 7714 10124
rect 7751 10112 7779 10152
rect 7828 10149 7840 10183
rect 7874 10180 7886 10183
rect 8294 10180 8300 10192
rect 7874 10152 8300 10180
rect 7874 10149 7886 10152
rect 7828 10143 7886 10149
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 8404 10180 8432 10220
rect 8496 10220 9781 10248
rect 8496 10180 8524 10220
rect 9769 10217 9781 10220
rect 9815 10217 9827 10251
rect 9769 10211 9827 10217
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10965 10251 11023 10257
rect 10965 10248 10977 10251
rect 10183 10220 10977 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10965 10217 10977 10220
rect 11011 10217 11023 10251
rect 10965 10211 11023 10217
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 12529 10251 12587 10257
rect 12529 10248 12541 10251
rect 12492 10220 12541 10248
rect 12492 10208 12498 10220
rect 12529 10217 12541 10220
rect 12575 10217 12587 10251
rect 13354 10248 13360 10260
rect 13315 10220 13360 10248
rect 12529 10211 12587 10217
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 13725 10251 13783 10257
rect 13725 10217 13737 10251
rect 13771 10248 13783 10251
rect 13906 10248 13912 10260
rect 13771 10220 13912 10248
rect 13771 10217 13783 10220
rect 13725 10211 13783 10217
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 15654 10208 15660 10260
rect 15712 10248 15718 10260
rect 15841 10251 15899 10257
rect 15841 10248 15853 10251
rect 15712 10220 15853 10248
rect 15712 10208 15718 10220
rect 15841 10217 15853 10220
rect 15887 10217 15899 10251
rect 15841 10211 15899 10217
rect 16850 10208 16856 10260
rect 16908 10248 16914 10260
rect 17221 10251 17279 10257
rect 17221 10248 17233 10251
rect 16908 10220 17233 10248
rect 16908 10208 16914 10220
rect 17221 10217 17233 10220
rect 17267 10217 17279 10251
rect 17221 10211 17279 10217
rect 17681 10251 17739 10257
rect 17681 10217 17693 10251
rect 17727 10248 17739 10251
rect 18414 10248 18420 10260
rect 17727 10220 18420 10248
rect 17727 10217 17739 10220
rect 17681 10211 17739 10217
rect 8404 10152 8524 10180
rect 8938 10140 8944 10192
rect 8996 10140 9002 10192
rect 10686 10140 10692 10192
rect 10744 10180 10750 10192
rect 11425 10183 11483 10189
rect 11425 10180 11437 10183
rect 10744 10152 11437 10180
rect 10744 10140 10750 10152
rect 11425 10149 11437 10152
rect 11471 10149 11483 10183
rect 11425 10143 11483 10149
rect 11532 10152 12839 10180
rect 8956 10112 8984 10140
rect 11330 10112 11336 10124
rect 7751 10084 8892 10112
rect 8956 10084 10548 10112
rect 11291 10084 11336 10112
rect 5442 10044 5448 10056
rect 5403 10016 5448 10044
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10044 5687 10047
rect 5994 10044 6000 10056
rect 5675 10016 6000 10044
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6362 10004 6368 10056
rect 6420 10044 6426 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6420 10016 6837 10044
rect 6420 10004 6426 10016
rect 6825 10013 6837 10016
rect 6871 10044 6883 10047
rect 7668 10044 7696 10072
rect 6871 10016 7696 10044
rect 8864 10044 8892 10084
rect 9398 10044 9404 10056
rect 8864 10016 9404 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 4430 9936 4436 9988
rect 4488 9976 4494 9988
rect 5350 9976 5356 9988
rect 4488 9948 5356 9976
rect 4488 9936 4494 9948
rect 5350 9936 5356 9948
rect 5408 9936 5414 9988
rect 5534 9936 5540 9988
rect 5592 9976 5598 9988
rect 7282 9976 7288 9988
rect 5592 9948 7288 9976
rect 5592 9936 5598 9948
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 9674 9976 9680 9988
rect 8496 9948 9680 9976
rect 8496 9908 8524 9948
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 10244 9976 10272 10007
rect 10318 10004 10324 10056
rect 10376 10044 10382 10056
rect 10520 10044 10548 10084
rect 11330 10072 11336 10084
rect 11388 10072 11394 10124
rect 11532 10112 11560 10152
rect 12811 10112 12839 10152
rect 14458 10140 14464 10192
rect 14516 10180 14522 10192
rect 15102 10180 15108 10192
rect 14516 10152 15108 10180
rect 14516 10140 14522 10152
rect 15102 10140 15108 10152
rect 15160 10140 15166 10192
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 17696 10180 17724 10211
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 15344 10152 17724 10180
rect 15344 10140 15350 10152
rect 14642 10121 14648 10124
rect 13817 10115 13875 10121
rect 13817 10112 13829 10115
rect 11440 10084 11560 10112
rect 11808 10084 12756 10112
rect 12811 10084 13829 10112
rect 11440 10044 11468 10084
rect 11808 10056 11836 10084
rect 10376 10016 10421 10044
rect 10520 10016 11468 10044
rect 11609 10047 11667 10053
rect 10376 10004 10382 10016
rect 11609 10013 11621 10047
rect 11655 10044 11667 10047
rect 11790 10044 11796 10056
rect 11655 10016 11796 10044
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12250 10004 12256 10056
rect 12308 10044 12314 10056
rect 12434 10044 12440 10056
rect 12308 10016 12440 10044
rect 12308 10004 12314 10016
rect 12434 10004 12440 10016
rect 12492 10004 12498 10056
rect 12618 10044 12624 10056
rect 12579 10016 12624 10044
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 12728 10053 12756 10084
rect 13817 10081 13829 10084
rect 13863 10081 13875 10115
rect 13817 10075 13875 10081
rect 14620 10115 14648 10121
rect 14620 10081 14632 10115
rect 14620 10075 14648 10081
rect 14642 10072 14648 10075
rect 14700 10072 14706 10124
rect 16209 10115 16267 10121
rect 16209 10081 16221 10115
rect 16255 10112 16267 10115
rect 17126 10112 17132 10124
rect 16255 10084 17132 10112
rect 16255 10081 16267 10084
rect 16209 10075 16267 10081
rect 17126 10072 17132 10084
rect 17184 10072 17190 10124
rect 17218 10072 17224 10124
rect 17276 10112 17282 10124
rect 17589 10115 17647 10121
rect 17589 10112 17601 10115
rect 17276 10084 17601 10112
rect 17276 10072 17282 10084
rect 17589 10081 17601 10084
rect 17635 10081 17647 10115
rect 17589 10075 17647 10081
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 13909 10047 13967 10053
rect 13909 10044 13921 10047
rect 13596 10016 13921 10044
rect 13596 10004 13602 10016
rect 13909 10013 13921 10016
rect 13955 10013 13967 10047
rect 16298 10044 16304 10056
rect 16259 10016 16304 10044
rect 13909 10007 13967 10013
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 16482 10044 16488 10056
rect 16443 10016 16488 10044
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 17770 10044 17776 10056
rect 17731 10016 17776 10044
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 12161 9979 12219 9985
rect 12161 9976 12173 9979
rect 10244 9948 12173 9976
rect 12161 9945 12173 9948
rect 12207 9945 12219 9979
rect 12161 9939 12219 9945
rect 12268 9948 15056 9976
rect 8938 9908 8944 9920
rect 3988 9880 8524 9908
rect 8899 9880 8944 9908
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 10686 9868 10692 9920
rect 10744 9908 10750 9920
rect 12268 9908 12296 9948
rect 10744 9880 12296 9908
rect 10744 9868 10750 9880
rect 13722 9868 13728 9920
rect 13780 9908 13786 9920
rect 14691 9911 14749 9917
rect 14691 9908 14703 9911
rect 13780 9880 14703 9908
rect 13780 9868 13786 9880
rect 14691 9877 14703 9880
rect 14737 9877 14749 9911
rect 15028 9908 15056 9948
rect 18506 9908 18512 9920
rect 15028 9880 18512 9908
rect 14691 9871 14749 9877
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 3050 9664 3056 9716
rect 3108 9704 3114 9716
rect 3697 9707 3755 9713
rect 3697 9704 3709 9707
rect 3108 9676 3709 9704
rect 3108 9664 3114 9676
rect 3697 9673 3709 9676
rect 3743 9673 3755 9707
rect 3697 9667 3755 9673
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 5442 9704 5448 9716
rect 4948 9676 5304 9704
rect 5403 9676 5448 9704
rect 4948 9664 4954 9676
rect 3237 9639 3295 9645
rect 3237 9605 3249 9639
rect 3283 9605 3295 9639
rect 5276 9636 5304 9676
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 7024 9676 9628 9704
rect 7024 9636 7052 9676
rect 5276 9608 7052 9636
rect 8849 9639 8907 9645
rect 3237 9599 3295 9605
rect 8849 9605 8861 9639
rect 8895 9636 8907 9639
rect 9122 9636 9128 9648
rect 8895 9608 9128 9636
rect 8895 9605 8907 9608
rect 8849 9599 8907 9605
rect 3252 9568 3280 9599
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 9600 9636 9628 9676
rect 10594 9664 10600 9716
rect 10652 9704 10658 9716
rect 10962 9704 10968 9716
rect 10652 9676 10968 9704
rect 10652 9664 10658 9676
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 12618 9704 12624 9716
rect 12483 9676 12624 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 12618 9664 12624 9676
rect 12676 9664 12682 9716
rect 15562 9664 15568 9716
rect 15620 9704 15626 9716
rect 15657 9707 15715 9713
rect 15657 9704 15669 9707
rect 15620 9676 15669 9704
rect 15620 9664 15626 9676
rect 15657 9673 15669 9676
rect 15703 9673 15715 9707
rect 15657 9667 15715 9673
rect 9674 9636 9680 9648
rect 9600 9608 9680 9636
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 9769 9639 9827 9645
rect 9769 9605 9781 9639
rect 9815 9605 9827 9639
rect 9769 9599 9827 9605
rect 10689 9639 10747 9645
rect 10689 9605 10701 9639
rect 10735 9636 10747 9639
rect 11330 9636 11336 9648
rect 10735 9608 11336 9636
rect 10735 9605 10747 9608
rect 10689 9599 10747 9605
rect 3326 9568 3332 9580
rect 3239 9540 3332 9568
rect 3326 9528 3332 9540
rect 3384 9568 3390 9580
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 3384 9540 4261 9568
rect 3384 9528 3390 9540
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9568 6147 9571
rect 6362 9568 6368 9580
rect 6135 9540 6368 9568
rect 6135 9537 6147 9540
rect 6089 9531 6147 9537
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 8938 9528 8944 9580
rect 8996 9568 9002 9580
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 8996 9540 9413 9568
rect 8996 9528 9002 9540
rect 9401 9537 9413 9540
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 1857 9503 1915 9509
rect 1857 9500 1869 9503
rect 1636 9472 1869 9500
rect 1636 9460 1642 9472
rect 1857 9469 1869 9472
rect 1903 9500 1915 9503
rect 2406 9500 2412 9512
rect 1903 9472 2412 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 2406 9460 2412 9472
rect 2464 9500 2470 9512
rect 4062 9500 4068 9512
rect 2464 9472 4068 9500
rect 2464 9460 2470 9472
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 5350 9500 5356 9512
rect 5311 9472 5356 9500
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 7009 9503 7067 9509
rect 5736 9472 6960 9500
rect 2124 9435 2182 9441
rect 2124 9401 2136 9435
rect 2170 9432 2182 9435
rect 2958 9432 2964 9444
rect 2170 9404 2964 9432
rect 2170 9401 2182 9404
rect 2124 9395 2182 9401
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 4154 9432 4160 9444
rect 4115 9404 4160 9432
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 5736 9432 5764 9472
rect 5092 9404 5764 9432
rect 5813 9435 5871 9441
rect 5092 9376 5120 9404
rect 5813 9401 5825 9435
rect 5859 9432 5871 9435
rect 6730 9432 6736 9444
rect 5859 9404 6736 9432
rect 5859 9401 5871 9404
rect 5813 9395 5871 9401
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9364 4123 9367
rect 5074 9364 5080 9376
rect 4111 9336 5080 9364
rect 4111 9333 4123 9336
rect 4065 9327 4123 9333
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5258 9364 5264 9376
rect 5215 9336 5264 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 5960 9336 6005 9364
rect 5960 9324 5966 9336
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6638 9364 6644 9376
rect 6236 9336 6644 9364
rect 6236 9324 6242 9336
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 6932 9364 6960 9472
rect 7009 9469 7021 9503
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 7276 9503 7334 9509
rect 7276 9469 7288 9503
rect 7322 9500 7334 9503
rect 8956 9500 8984 9528
rect 7322 9472 8984 9500
rect 9784 9500 9812 9599
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 11514 9596 11520 9648
rect 11572 9636 11578 9648
rect 11698 9636 11704 9648
rect 11572 9608 11704 9636
rect 11572 9596 11578 9608
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 12161 9639 12219 9645
rect 12161 9605 12173 9639
rect 12207 9636 12219 9639
rect 13630 9636 13636 9648
rect 12207 9608 13636 9636
rect 12207 9605 12219 9608
rect 12161 9599 12219 9605
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 16758 9636 16764 9648
rect 16719 9608 16764 9636
rect 16758 9596 16764 9608
rect 16816 9596 16822 9648
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 11146 9568 11152 9580
rect 10459 9540 11152 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 11146 9528 11152 9540
rect 11204 9528 11210 9580
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9568 11299 9571
rect 12342 9568 12348 9580
rect 11287 9540 12348 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 12342 9528 12348 9540
rect 12400 9568 12406 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12400 9540 13001 9568
rect 12400 9528 12406 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13814 9528 13820 9580
rect 13872 9568 13878 9580
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 13872 9540 14289 9568
rect 13872 9528 13878 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 17218 9568 17224 9580
rect 16163 9540 17224 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 17218 9528 17224 9540
rect 17276 9528 17282 9580
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9568 17371 9571
rect 17770 9568 17776 9580
rect 17359 9540 17776 9568
rect 17359 9537 17371 9540
rect 17313 9531 17371 9537
rect 11882 9500 11888 9512
rect 9784 9472 11888 9500
rect 7322 9469 7334 9472
rect 7276 9463 7334 9469
rect 7024 9432 7052 9463
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 12066 9500 12072 9512
rect 12027 9472 12072 9500
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 12802 9500 12808 9512
rect 12360 9472 12808 9500
rect 12360 9444 12388 9472
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 14544 9503 14602 9509
rect 14544 9469 14556 9503
rect 14590 9469 14602 9503
rect 16482 9500 16488 9512
rect 14544 9463 14602 9469
rect 15672 9472 16488 9500
rect 7558 9432 7564 9444
rect 7024 9404 7564 9432
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 9217 9435 9275 9441
rect 9217 9432 9229 9435
rect 7668 9404 9229 9432
rect 7668 9364 7696 9404
rect 9217 9401 9229 9404
rect 9263 9432 9275 9435
rect 9398 9432 9404 9444
rect 9263 9404 9404 9432
rect 9263 9401 9275 9404
rect 9217 9395 9275 9401
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 12158 9432 12164 9444
rect 12119 9404 12164 9432
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 12342 9392 12348 9444
rect 12400 9392 12406 9444
rect 12897 9435 12955 9441
rect 12897 9432 12909 9435
rect 12728 9404 12909 9432
rect 12728 9376 12756 9404
rect 12897 9401 12909 9404
rect 12943 9401 12955 9435
rect 12897 9395 12955 9401
rect 6932 9336 7696 9364
rect 8389 9367 8447 9373
rect 8389 9333 8401 9367
rect 8435 9364 8447 9367
rect 8478 9364 8484 9376
rect 8435 9336 8484 9364
rect 8435 9333 8447 9336
rect 8389 9327 8447 9333
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 9306 9364 9312 9376
rect 9267 9336 9312 9364
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 10134 9364 10140 9376
rect 10095 9336 10140 9364
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10229 9367 10287 9373
rect 10229 9333 10241 9367
rect 10275 9364 10287 9367
rect 10410 9364 10416 9376
rect 10275 9336 10416 9364
rect 10275 9333 10287 9336
rect 10229 9327 10287 9333
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 11054 9364 11060 9376
rect 11015 9336 11060 9364
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 11514 9364 11520 9376
rect 11195 9336 11520 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 11885 9367 11943 9373
rect 11885 9364 11897 9367
rect 11756 9336 11897 9364
rect 11756 9324 11762 9336
rect 11885 9333 11897 9336
rect 11931 9333 11943 9367
rect 11885 9327 11943 9333
rect 12710 9324 12716 9376
rect 12768 9324 12774 9376
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 13354 9364 13360 9376
rect 12851 9336 13360 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 13630 9364 13636 9376
rect 13591 9336 13636 9364
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 14559 9364 14587 9463
rect 15672 9364 15700 9472
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 17328 9500 17356 9531
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 16724 9472 17356 9500
rect 16724 9460 16730 9472
rect 16114 9392 16120 9444
rect 16172 9432 16178 9444
rect 17129 9435 17187 9441
rect 17129 9432 17141 9435
rect 16172 9404 17141 9432
rect 16172 9392 16178 9404
rect 17129 9401 17141 9404
rect 17175 9401 17187 9435
rect 17129 9395 17187 9401
rect 17218 9392 17224 9444
rect 17276 9432 17282 9444
rect 17276 9404 17321 9432
rect 17276 9392 17282 9404
rect 14559 9336 15700 9364
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 2958 9160 2964 9172
rect 2919 9132 2964 9160
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9129 5503 9163
rect 5902 9160 5908 9172
rect 5863 9132 5908 9160
rect 5445 9123 5503 9129
rect 1848 9095 1906 9101
rect 1848 9061 1860 9095
rect 1894 9092 1906 9095
rect 2130 9092 2136 9104
rect 1894 9064 2136 9092
rect 1894 9061 1906 9064
rect 1848 9055 1906 9061
rect 2130 9052 2136 9064
rect 2188 9092 2194 9104
rect 5460 9092 5488 9123
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 6362 9160 6368 9172
rect 6323 9132 6368 9160
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 7101 9163 7159 9169
rect 7101 9160 7113 9163
rect 6788 9132 7113 9160
rect 6788 9120 6794 9132
rect 7101 9129 7113 9132
rect 7147 9129 7159 9163
rect 7101 9123 7159 9129
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 7340 9132 8309 9160
rect 7340 9120 7346 9132
rect 8297 9129 8309 9132
rect 8343 9129 8355 9163
rect 8297 9123 8355 9129
rect 8389 9163 8447 9169
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 9030 9160 9036 9172
rect 8435 9132 9036 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 10505 9163 10563 9169
rect 10505 9129 10517 9163
rect 10551 9160 10563 9163
rect 11054 9160 11060 9172
rect 10551 9132 11060 9160
rect 10551 9129 10563 9132
rect 10505 9123 10563 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11146 9120 11152 9172
rect 11204 9160 11210 9172
rect 11330 9160 11336 9172
rect 11204 9132 11336 9160
rect 11204 9120 11210 9132
rect 11330 9120 11336 9132
rect 11388 9160 11394 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 11388 9132 12357 9160
rect 11388 9120 11394 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 12897 9163 12955 9169
rect 12897 9129 12909 9163
rect 12943 9160 12955 9163
rect 13354 9160 13360 9172
rect 12943 9132 13360 9160
rect 12943 9129 12955 9132
rect 12897 9123 12955 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 14093 9163 14151 9169
rect 14093 9160 14105 9163
rect 13872 9132 14105 9160
rect 13872 9120 13878 9132
rect 14093 9129 14105 9132
rect 14139 9160 14151 9163
rect 16666 9160 16672 9172
rect 14139 9132 15240 9160
rect 16627 9132 16672 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 2188 9064 5488 9092
rect 2188 9052 2194 9064
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 7561 9095 7619 9101
rect 7561 9092 7573 9095
rect 5868 9064 7573 9092
rect 5868 9052 5874 9064
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 4338 9033 4344 9036
rect 4332 9024 4344 9033
rect 4299 8996 4344 9024
rect 4332 8987 4344 8996
rect 4338 8984 4344 8987
rect 4396 8984 4402 9036
rect 5902 8984 5908 9036
rect 5960 9024 5966 9036
rect 6273 9027 6331 9033
rect 6273 9024 6285 9027
rect 5960 8996 6285 9024
rect 5960 8984 5966 8996
rect 6273 8993 6285 8996
rect 6319 8993 6331 9027
rect 6273 8987 6331 8993
rect 6656 8968 6684 9064
rect 7561 9061 7573 9064
rect 7607 9092 7619 9095
rect 11514 9092 11520 9104
rect 7607 9064 11520 9092
rect 7607 9061 7619 9064
rect 7561 9055 7619 9061
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 11698 9052 11704 9104
rect 11756 9092 11762 9104
rect 11756 9064 14320 9092
rect 11756 9052 11762 9064
rect 7469 9027 7527 9033
rect 7469 8993 7481 9027
rect 7515 9024 7527 9027
rect 8202 9024 8208 9036
rect 7515 8996 8208 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 9024 8355 9027
rect 8757 9027 8815 9033
rect 8757 9024 8769 9027
rect 8343 8996 8769 9024
rect 8343 8993 8355 8996
rect 8297 8987 8355 8993
rect 8757 8993 8769 8996
rect 8803 9024 8815 9027
rect 9030 9024 9036 9036
rect 8803 8996 9036 9024
rect 8803 8993 8815 8996
rect 8757 8987 8815 8993
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9180 8996 10057 9024
rect 9180 8984 9186 8996
rect 10045 8993 10057 8996
rect 10091 9024 10103 9027
rect 10686 9024 10692 9036
rect 10091 8996 10692 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 10836 8996 10977 9024
rect 10836 8984 10842 8996
rect 10965 8993 10977 8996
rect 11011 8993 11023 9027
rect 11232 9027 11290 9033
rect 11232 9024 11244 9027
rect 10965 8987 11023 8993
rect 11072 8996 11244 9024
rect 4062 8956 4068 8968
rect 4023 8928 4068 8956
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 6549 8959 6607 8965
rect 6549 8956 6561 8959
rect 6512 8928 6561 8956
rect 6512 8916 6518 8928
rect 6549 8925 6561 8928
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6564 8888 6592 8919
rect 6638 8916 6644 8968
rect 6696 8916 6702 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 8849 8959 8907 8965
rect 8849 8925 8861 8959
rect 8895 8925 8907 8959
rect 8849 8919 8907 8925
rect 7668 8888 7696 8919
rect 6564 8860 7696 8888
rect 8864 8888 8892 8919
rect 8938 8916 8944 8968
rect 8996 8956 9002 8968
rect 8996 8928 9041 8956
rect 8996 8916 9002 8928
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9732 8928 10149 8956
rect 9732 8916 9738 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 11072 8956 11100 8996
rect 11232 8993 11244 8996
rect 11278 9024 11290 9027
rect 11606 9024 11612 9036
rect 11278 8996 11612 9024
rect 11278 8993 11290 8996
rect 11232 8987 11290 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 13814 9024 13820 9036
rect 13311 8996 13820 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 14292 9033 14320 9064
rect 14277 9027 14335 9033
rect 14277 8993 14289 9027
rect 14323 8993 14335 9027
rect 14277 8987 14335 8993
rect 14461 9027 14519 9033
rect 14461 8993 14473 9027
rect 14507 8993 14519 9027
rect 15212 9024 15240 9132
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 17126 9160 17132 9172
rect 17087 9132 17132 9160
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 17497 9163 17555 9169
rect 17497 9160 17509 9163
rect 17276 9132 17509 9160
rect 17276 9120 17282 9132
rect 17497 9129 17509 9132
rect 17543 9129 17555 9163
rect 17497 9123 17555 9129
rect 15556 9095 15614 9101
rect 15556 9061 15568 9095
rect 15602 9092 15614 9095
rect 15654 9092 15660 9104
rect 15602 9064 15660 9092
rect 15602 9061 15614 9064
rect 15556 9055 15614 9061
rect 15654 9052 15660 9064
rect 15712 9052 15718 9104
rect 17586 9052 17592 9104
rect 17644 9052 17650 9104
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 15212 8996 15301 9024
rect 14461 8987 14519 8993
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 10367 8928 11100 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 10042 8888 10048 8900
rect 8864 8860 10048 8888
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 6454 8820 6460 8832
rect 5224 8792 6460 8820
rect 5224 8780 5230 8792
rect 6454 8780 6460 8792
rect 6512 8820 6518 8832
rect 8864 8820 8892 8860
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 10152 8888 10180 8919
rect 10980 8900 11008 8928
rect 13078 8916 13084 8968
rect 13136 8956 13142 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 13136 8928 13369 8956
rect 13136 8916 13142 8928
rect 10152 8860 10916 8888
rect 6512 8792 8892 8820
rect 9677 8823 9735 8829
rect 6512 8780 6518 8792
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 10778 8820 10784 8832
rect 9723 8792 10784 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 10888 8820 10916 8860
rect 10962 8848 10968 8900
rect 11020 8848 11026 8900
rect 12158 8820 12164 8832
rect 10888 8792 12164 8820
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 13280 8820 13308 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13538 8956 13544 8968
rect 13499 8928 13544 8956
rect 13357 8919 13415 8925
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 14476 8956 14504 8987
rect 15378 8984 15384 9036
rect 15436 8984 15442 9036
rect 17604 9024 17632 9052
rect 17604 8996 17908 9024
rect 15396 8956 15424 8984
rect 17586 8956 17592 8968
rect 14476 8928 15424 8956
rect 17547 8928 17592 8956
rect 17586 8916 17592 8928
rect 17644 8916 17650 8968
rect 17770 8956 17776 8968
rect 17731 8928 17776 8956
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 13814 8820 13820 8832
rect 13280 8792 13820 8820
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 14645 8823 14703 8829
rect 14645 8820 14657 8823
rect 14516 8792 14657 8820
rect 14516 8780 14522 8792
rect 14645 8789 14657 8792
rect 14691 8789 14703 8823
rect 14645 8783 14703 8789
rect 17770 8780 17776 8832
rect 17828 8820 17834 8832
rect 17880 8820 17908 8996
rect 17828 8792 17908 8820
rect 17828 8780 17834 8792
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 2096 8588 4261 8616
rect 2096 8576 2102 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 5408 8588 9873 8616
rect 5408 8576 5414 8588
rect 9861 8585 9873 8588
rect 9907 8616 9919 8619
rect 12066 8616 12072 8628
rect 9907 8588 12072 8616
rect 9907 8585 9919 8588
rect 9861 8579 9919 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 12897 8619 12955 8625
rect 12897 8616 12909 8619
rect 12768 8588 12909 8616
rect 12768 8576 12774 8588
rect 12897 8585 12909 8588
rect 12943 8585 12955 8619
rect 12897 8579 12955 8585
rect 15654 8576 15660 8628
rect 15712 8616 15718 8628
rect 15933 8619 15991 8625
rect 15933 8616 15945 8619
rect 15712 8588 15945 8616
rect 15712 8576 15718 8588
rect 15933 8585 15945 8588
rect 15979 8585 15991 8619
rect 15933 8579 15991 8585
rect 16206 8576 16212 8628
rect 16264 8576 16270 8628
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 16393 8619 16451 8625
rect 16393 8616 16405 8619
rect 16356 8588 16405 8616
rect 16356 8576 16362 8588
rect 16393 8585 16405 8588
rect 16439 8585 16451 8619
rect 16393 8579 16451 8585
rect 1578 8508 1584 8560
rect 1636 8548 1642 8560
rect 1857 8551 1915 8557
rect 1857 8548 1869 8551
rect 1636 8520 1869 8548
rect 1636 8508 1642 8520
rect 1857 8517 1869 8520
rect 1903 8517 1915 8551
rect 1857 8511 1915 8517
rect 4338 8508 4344 8560
rect 4396 8548 4402 8560
rect 7009 8551 7067 8557
rect 7009 8548 7021 8551
rect 4396 8520 7021 8548
rect 4396 8508 4402 8520
rect 7009 8517 7021 8520
rect 7055 8517 7067 8551
rect 7009 8511 7067 8517
rect 7377 8551 7435 8557
rect 7377 8517 7389 8551
rect 7423 8517 7435 8551
rect 7377 8511 7435 8517
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8480 2559 8483
rect 2958 8480 2964 8492
rect 2547 8452 2964 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 3384 8452 3709 8480
rect 3384 8440 3390 8452
rect 3697 8449 3709 8452
rect 3743 8480 3755 8483
rect 4246 8480 4252 8492
rect 3743 8452 4252 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 4246 8440 4252 8452
rect 4304 8480 4310 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4304 8452 4905 8480
rect 4304 8440 4310 8452
rect 4893 8449 4905 8452
rect 4939 8480 4951 8483
rect 5166 8480 5172 8492
rect 4939 8452 5172 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 5994 8440 6000 8492
rect 6052 8480 6058 8492
rect 6089 8483 6147 8489
rect 6089 8480 6101 8483
rect 6052 8452 6101 8480
rect 6052 8440 6058 8452
rect 6089 8449 6101 8452
rect 6135 8449 6147 8483
rect 6089 8443 6147 8449
rect 7392 8424 7420 8511
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 10042 8548 10048 8560
rect 9364 8520 10048 8548
rect 9364 8508 9370 8520
rect 10042 8508 10048 8520
rect 10100 8508 10106 8560
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 11664 8520 11805 8548
rect 11664 8508 11670 8520
rect 11793 8517 11805 8520
rect 11839 8517 11851 8551
rect 13998 8548 14004 8560
rect 11793 8511 11851 8517
rect 11900 8520 14004 8548
rect 7834 8480 7840 8492
rect 7795 8452 7840 8480
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 8018 8480 8024 8492
rect 7979 8452 8024 8480
rect 8018 8440 8024 8452
rect 8076 8440 8082 8492
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 10413 8483 10471 8489
rect 10413 8480 10425 8483
rect 9732 8452 10425 8480
rect 9732 8440 9738 8452
rect 10413 8449 10425 8452
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 11514 8440 11520 8492
rect 11572 8480 11578 8492
rect 11900 8480 11928 8520
rect 13998 8508 14004 8520
rect 14056 8508 14062 8560
rect 13538 8480 13544 8492
rect 11572 8452 11928 8480
rect 13499 8452 13544 8480
rect 11572 8440 11578 8452
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 13906 8440 13912 8492
rect 13964 8480 13970 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 13964 8452 14565 8480
rect 13964 8440 13970 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 16224 8424 16252 8576
rect 16666 8440 16672 8492
rect 16724 8480 16730 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16724 8452 16957 8480
rect 16724 8440 16730 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 3418 8412 3424 8424
rect 3379 8384 3424 8412
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 3513 8415 3571 8421
rect 3513 8381 3525 8415
rect 3559 8412 3571 8415
rect 3602 8412 3608 8424
rect 3559 8384 3608 8412
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 1486 8304 1492 8356
rect 1544 8344 1550 8356
rect 2317 8347 2375 8353
rect 2317 8344 2329 8347
rect 1544 8316 2329 8344
rect 1544 8304 1550 8316
rect 2317 8313 2329 8316
rect 2363 8313 2375 8347
rect 2317 8307 2375 8313
rect 2958 8304 2964 8356
rect 3016 8344 3022 8356
rect 3528 8344 3556 8375
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 4617 8415 4675 8421
rect 4617 8381 4629 8415
rect 4663 8412 4675 8415
rect 4706 8412 4712 8424
rect 4663 8384 4712 8412
rect 4663 8381 4675 8384
rect 4617 8375 4675 8381
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8412 6883 8415
rect 7282 8412 7288 8424
rect 6871 8384 7288 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 7374 8372 7380 8424
rect 7432 8372 7438 8424
rect 8570 8412 8576 8424
rect 7576 8384 7880 8412
rect 8531 8384 8576 8412
rect 3016 8316 3556 8344
rect 3016 8304 3022 8316
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 5902 8344 5908 8356
rect 4304 8316 5908 8344
rect 4304 8304 4310 8316
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 5997 8347 6055 8353
rect 5997 8313 6009 8347
rect 6043 8344 6055 8347
rect 6362 8344 6368 8356
rect 6043 8316 6368 8344
rect 6043 8313 6055 8316
rect 5997 8307 6055 8313
rect 6362 8304 6368 8316
rect 6420 8344 6426 8356
rect 7576 8344 7604 8384
rect 6420 8316 7604 8344
rect 6420 8304 6426 8316
rect 7650 8304 7656 8356
rect 7708 8344 7714 8356
rect 7745 8347 7803 8353
rect 7745 8344 7757 8347
rect 7708 8316 7757 8344
rect 7708 8304 7714 8316
rect 7745 8313 7757 8316
rect 7791 8313 7803 8347
rect 7852 8344 7880 8384
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 9398 8372 9404 8424
rect 9456 8412 9462 8424
rect 10686 8421 10692 8424
rect 10680 8412 10692 8421
rect 9456 8384 10548 8412
rect 10647 8384 10692 8412
rect 9456 8372 9462 8384
rect 10134 8344 10140 8356
rect 7852 8316 10140 8344
rect 7745 8307 7803 8313
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 10520 8344 10548 8384
rect 10680 8375 10692 8384
rect 10686 8372 10692 8375
rect 10744 8372 10750 8424
rect 12342 8372 12348 8424
rect 12400 8412 12406 8424
rect 12710 8412 12716 8424
rect 12400 8384 12716 8412
rect 12400 8372 12406 8384
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 15746 8412 15752 8424
rect 14660 8384 15752 8412
rect 13265 8347 13323 8353
rect 13265 8344 13277 8347
rect 10520 8316 13277 8344
rect 13265 8313 13277 8316
rect 13311 8344 13323 8347
rect 14660 8344 14688 8384
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 16206 8372 16212 8424
rect 16264 8372 16270 8424
rect 13311 8316 14688 8344
rect 14820 8347 14878 8353
rect 13311 8313 13323 8316
rect 13265 8307 13323 8313
rect 14820 8313 14832 8347
rect 14866 8344 14878 8347
rect 15102 8344 15108 8356
rect 14866 8316 15108 8344
rect 14866 8313 14878 8316
rect 14820 8307 14878 8313
rect 15102 8304 15108 8316
rect 15160 8304 15166 8356
rect 16666 8304 16672 8356
rect 16724 8344 16730 8356
rect 16853 8347 16911 8353
rect 16853 8344 16865 8347
rect 16724 8316 16865 8344
rect 16724 8304 16730 8316
rect 16853 8313 16865 8316
rect 16899 8313 16911 8347
rect 16853 8307 16911 8313
rect 2222 8276 2228 8288
rect 2183 8248 2228 8276
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 3050 8276 3056 8288
rect 3011 8248 3056 8276
rect 3050 8236 3056 8248
rect 3108 8236 3114 8288
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 5534 8276 5540 8288
rect 4764 8248 4809 8276
rect 5495 8248 5540 8276
rect 4764 8236 4770 8248
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 7558 8236 7564 8288
rect 7616 8276 7622 8288
rect 11606 8276 11612 8288
rect 7616 8248 11612 8276
rect 7616 8236 7622 8248
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 12066 8236 12072 8288
rect 12124 8276 12130 8288
rect 12250 8276 12256 8288
rect 12124 8248 12256 8276
rect 12124 8236 12130 8248
rect 12250 8236 12256 8248
rect 12308 8236 12314 8288
rect 13357 8279 13415 8285
rect 13357 8245 13369 8279
rect 13403 8276 13415 8279
rect 13538 8276 13544 8288
rect 13403 8248 13544 8276
rect 13403 8245 13415 8248
rect 13357 8239 13415 8245
rect 13538 8236 13544 8248
rect 13596 8276 13602 8288
rect 15378 8276 15384 8288
rect 13596 8248 15384 8276
rect 13596 8236 13602 8248
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 16758 8276 16764 8288
rect 16719 8248 16764 8276
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 4525 8075 4583 8081
rect 4525 8072 4537 8075
rect 1995 8044 4537 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 4525 8041 4537 8044
rect 4571 8041 4583 8075
rect 4525 8035 4583 8041
rect 4985 8075 5043 8081
rect 4985 8041 4997 8075
rect 5031 8072 5043 8075
rect 5534 8072 5540 8084
rect 5031 8044 5540 8072
rect 5031 8041 5043 8044
rect 4985 8035 5043 8041
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 7101 8075 7159 8081
rect 7101 8072 7113 8075
rect 5644 8044 7113 8072
rect 1857 8007 1915 8013
rect 1857 7973 1869 8007
rect 1903 8004 1915 8007
rect 2038 8004 2044 8016
rect 1903 7976 2044 8004
rect 1903 7973 1915 7976
rect 1857 7967 1915 7973
rect 2038 7964 2044 7976
rect 2096 7964 2102 8016
rect 3602 8004 3608 8016
rect 3252 7976 3608 8004
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 2130 7868 2136 7880
rect 2091 7840 2136 7868
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 3068 7800 3096 7899
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7868 3203 7871
rect 3252 7868 3280 7976
rect 3602 7964 3608 7976
rect 3660 7964 3666 8016
rect 4893 7939 4951 7945
rect 4893 7905 4905 7939
rect 4939 7936 4951 7939
rect 5442 7936 5448 7948
rect 4939 7908 5448 7936
rect 4939 7905 4951 7908
rect 4893 7899 4951 7905
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 3191 7840 3280 7868
rect 3191 7837 3203 7840
rect 3145 7831 3203 7837
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 5166 7868 5172 7880
rect 3384 7840 3429 7868
rect 5079 7840 5172 7868
rect 3384 7828 3390 7840
rect 5166 7828 5172 7840
rect 5224 7868 5230 7880
rect 5644 7868 5672 8044
rect 7101 8041 7113 8044
rect 7147 8041 7159 8075
rect 7101 8035 7159 8041
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7432 8044 8033 8072
rect 7432 8032 7438 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 8021 8035 8079 8041
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 6178 7964 6184 8016
rect 6236 8004 6242 8016
rect 8956 8004 8984 8035
rect 10134 8032 10140 8084
rect 10192 8072 10198 8084
rect 11514 8072 11520 8084
rect 10192 8044 11520 8072
rect 10192 8032 10198 8044
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 12161 8075 12219 8081
rect 12161 8072 12173 8075
rect 11940 8044 12173 8072
rect 11940 8032 11946 8044
rect 12161 8041 12173 8044
rect 12207 8041 12219 8075
rect 12161 8035 12219 8041
rect 15749 8075 15807 8081
rect 15749 8041 15761 8075
rect 15795 8072 15807 8075
rect 16758 8072 16764 8084
rect 15795 8044 16764 8072
rect 15795 8041 15807 8044
rect 15749 8035 15807 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 16945 8075 17003 8081
rect 16945 8041 16957 8075
rect 16991 8072 17003 8075
rect 17586 8072 17592 8084
rect 16991 8044 17592 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 11054 8004 11060 8016
rect 6236 7976 8984 8004
rect 9048 7976 11060 8004
rect 6236 7964 6242 7976
rect 5994 7945 6000 7948
rect 5988 7936 6000 7945
rect 5955 7908 6000 7936
rect 5988 7899 6000 7908
rect 6052 7936 6058 7948
rect 6362 7936 6368 7948
rect 6052 7908 6368 7936
rect 5994 7896 6000 7899
rect 6052 7896 6058 7908
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 7190 7896 7196 7948
rect 7248 7936 7254 7948
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 7248 7908 7941 7936
rect 7248 7896 7254 7908
rect 7929 7905 7941 7908
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 8478 7896 8484 7948
rect 8536 7936 8542 7948
rect 8757 7939 8815 7945
rect 8757 7936 8769 7939
rect 8536 7908 8769 7936
rect 8536 7896 8542 7908
rect 8757 7905 8769 7908
rect 8803 7936 8815 7939
rect 9048 7936 9076 7976
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 13078 7964 13084 8016
rect 13136 8004 13142 8016
rect 13357 8007 13415 8013
rect 13357 8004 13369 8007
rect 13136 7976 13369 8004
rect 13136 7964 13142 7976
rect 13357 7973 13369 7976
rect 13403 7973 13415 8007
rect 13357 7967 13415 7973
rect 15286 7964 15292 8016
rect 15344 8004 15350 8016
rect 15470 8004 15476 8016
rect 15344 7976 15476 8004
rect 15344 7964 15350 7976
rect 15470 7964 15476 7976
rect 15528 8004 15534 8016
rect 17313 8007 17371 8013
rect 15528 7976 16252 8004
rect 15528 7964 15534 7976
rect 8803 7908 9076 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 9933 7939 9991 7945
rect 9933 7936 9945 7939
rect 9640 7908 9945 7936
rect 9640 7896 9646 7908
rect 9933 7905 9945 7908
rect 9979 7905 9991 7939
rect 12066 7936 12072 7948
rect 12027 7908 12072 7936
rect 9933 7899 9991 7905
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 13004 7908 13277 7936
rect 5224 7840 5672 7868
rect 5721 7871 5779 7877
rect 5224 7828 5230 7840
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 9674 7868 9680 7880
rect 8251 7840 8432 7868
rect 9635 7840 9680 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 4614 7800 4620 7812
rect 3068 7772 4620 7800
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 5736 7800 5764 7831
rect 5460 7772 5764 7800
rect 5460 7744 5488 7772
rect 2590 7692 2596 7744
rect 2648 7732 2654 7744
rect 2685 7735 2743 7741
rect 2685 7732 2697 7735
rect 2648 7704 2697 7732
rect 2648 7692 2654 7704
rect 2685 7701 2697 7704
rect 2731 7701 2743 7735
rect 2685 7695 2743 7701
rect 5442 7692 5448 7744
rect 5500 7692 5506 7744
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 8404 7732 8432 7840
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 11330 7868 11336 7880
rect 11112 7840 11336 7868
rect 11112 7828 11118 7840
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 11606 7828 11612 7880
rect 11664 7868 11670 7880
rect 12342 7877 12348 7880
rect 12299 7871 12348 7877
rect 11664 7840 11827 7868
rect 11664 7828 11670 7840
rect 8478 7760 8484 7812
rect 8536 7800 8542 7812
rect 9122 7800 9128 7812
rect 8536 7772 9128 7800
rect 8536 7760 8542 7772
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 10686 7732 10692 7744
rect 8404 7704 10692 7732
rect 10686 7692 10692 7704
rect 10744 7732 10750 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10744 7704 11069 7732
rect 10744 7692 10750 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 11606 7692 11612 7744
rect 11664 7732 11670 7744
rect 11701 7735 11759 7741
rect 11701 7732 11713 7735
rect 11664 7704 11713 7732
rect 11664 7692 11670 7704
rect 11701 7701 11713 7704
rect 11747 7701 11759 7735
rect 11799 7732 11827 7840
rect 12299 7837 12311 7871
rect 12345 7837 12348 7871
rect 12299 7831 12348 7837
rect 12342 7828 12348 7831
rect 12400 7828 12406 7880
rect 12894 7800 12900 7812
rect 12855 7772 12900 7800
rect 12894 7760 12900 7772
rect 12952 7760 12958 7812
rect 13004 7732 13032 7908
rect 13265 7905 13277 7908
rect 13311 7936 13323 7939
rect 13311 7908 13584 7936
rect 13311 7905 13323 7908
rect 13265 7899 13323 7905
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 13096 7840 13461 7868
rect 13096 7744 13124 7840
rect 13449 7837 13461 7840
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 13556 7800 13584 7908
rect 13998 7896 14004 7948
rect 14056 7936 14062 7948
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 14056 7908 14473 7936
rect 14056 7896 14062 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 14476 7868 14504 7899
rect 15010 7896 15016 7948
rect 15068 7936 15074 7948
rect 16117 7939 16175 7945
rect 16117 7936 16129 7939
rect 15068 7908 16129 7936
rect 15068 7896 15074 7908
rect 16117 7905 16129 7908
rect 16163 7905 16175 7939
rect 16224 7936 16252 7976
rect 17313 7973 17325 8007
rect 17359 8004 17371 8007
rect 17862 8004 17868 8016
rect 17359 7976 17868 8004
rect 17359 7973 17371 7976
rect 17313 7967 17371 7973
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 17405 7939 17463 7945
rect 17405 7936 17417 7939
rect 16224 7908 17417 7936
rect 16117 7899 16175 7905
rect 17405 7905 17417 7908
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 16209 7871 16267 7877
rect 16209 7868 16221 7871
rect 14476 7840 16221 7868
rect 16209 7837 16221 7840
rect 16255 7837 16267 7871
rect 16209 7831 16267 7837
rect 16301 7871 16359 7877
rect 16301 7837 16313 7871
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 13556 7772 15424 7800
rect 11799 7704 13032 7732
rect 11701 7695 11759 7701
rect 13078 7692 13084 7744
rect 13136 7692 13142 7744
rect 14645 7735 14703 7741
rect 14645 7701 14657 7735
rect 14691 7732 14703 7735
rect 15286 7732 15292 7744
rect 14691 7704 15292 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 15396 7732 15424 7772
rect 15654 7760 15660 7812
rect 15712 7800 15718 7812
rect 16316 7800 16344 7831
rect 17218 7800 17224 7812
rect 15712 7772 17224 7800
rect 15712 7760 15718 7772
rect 17218 7760 17224 7772
rect 17276 7800 17282 7812
rect 17512 7800 17540 7831
rect 17276 7772 17540 7800
rect 17276 7760 17282 7772
rect 17862 7732 17868 7744
rect 15396 7704 17868 7732
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 2222 7528 2228 7540
rect 2183 7500 2228 7528
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 4246 7488 4252 7540
rect 4304 7488 4310 7540
rect 4341 7531 4399 7537
rect 4341 7497 4353 7531
rect 4387 7528 4399 7531
rect 4706 7528 4712 7540
rect 4387 7500 4712 7528
rect 4387 7497 4399 7500
rect 4341 7491 4399 7497
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 5534 7528 5540 7540
rect 5495 7500 5540 7528
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 7190 7528 7196 7540
rect 7151 7500 7196 7528
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 8018 7488 8024 7540
rect 8076 7528 8082 7540
rect 9582 7528 9588 7540
rect 8076 7500 9588 7528
rect 8076 7488 8082 7500
rect 9582 7488 9588 7500
rect 9640 7528 9646 7540
rect 9769 7531 9827 7537
rect 9769 7528 9781 7531
rect 9640 7500 9781 7528
rect 9640 7488 9646 7500
rect 9769 7497 9781 7500
rect 9815 7497 9827 7531
rect 11701 7531 11759 7537
rect 9769 7491 9827 7497
rect 10336 7500 11284 7528
rect 4264 7460 4292 7488
rect 6638 7460 6644 7472
rect 1504 7432 4292 7460
rect 6012 7432 6644 7460
rect 1504 7333 1532 7432
rect 2130 7352 2136 7404
rect 2188 7392 2194 7404
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2188 7364 2789 7392
rect 2188 7352 2194 7364
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 4890 7392 4896 7404
rect 4847 7364 4896 7392
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7392 5043 7395
rect 5074 7392 5080 7404
rect 5031 7364 5080 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 6012 7401 6040 7432
rect 6638 7420 6644 7432
rect 6696 7420 6702 7472
rect 8202 7460 8208 7472
rect 6748 7432 8208 7460
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 6181 7395 6239 7401
rect 6181 7361 6193 7395
rect 6227 7392 6239 7395
rect 6362 7392 6368 7404
rect 6227 7364 6368 7392
rect 6227 7361 6239 7364
rect 6181 7355 6239 7361
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7293 1547 7327
rect 2590 7324 2596 7336
rect 2551 7296 2596 7324
rect 1489 7287 1547 7293
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7324 2743 7327
rect 3050 7324 3056 7336
rect 2731 7296 3056 7324
rect 2731 7293 2743 7296
rect 2685 7287 2743 7293
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 3418 7324 3424 7336
rect 3379 7296 3424 7324
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 5810 7284 5816 7336
rect 5868 7324 5874 7336
rect 5905 7327 5963 7333
rect 5905 7324 5917 7327
rect 5868 7296 5917 7324
rect 5868 7284 5874 7296
rect 5905 7293 5917 7296
rect 5951 7324 5963 7327
rect 6748 7324 6776 7432
rect 8202 7420 8208 7432
rect 8260 7420 8266 7472
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8018 7392 8024 7404
rect 7883 7364 8024 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 10336 7392 10364 7500
rect 11256 7460 11284 7500
rect 11701 7497 11713 7531
rect 11747 7528 11759 7531
rect 12342 7528 12348 7540
rect 11747 7500 12348 7528
rect 11747 7497 11759 7500
rect 11701 7491 11759 7497
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 13906 7528 13912 7540
rect 13740 7500 13912 7528
rect 11256 7432 13676 7460
rect 10336 7364 10456 7392
rect 5951 7296 6776 7324
rect 7561 7327 7619 7333
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 7561 7293 7573 7327
rect 7607 7324 7619 7327
rect 8294 7324 8300 7336
rect 7607 7296 8300 7324
rect 7607 7293 7619 7296
rect 7561 7287 7619 7293
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7324 8447 7327
rect 9214 7324 9220 7336
rect 8435 7296 9220 7324
rect 8435 7293 8447 7296
rect 8389 7287 8447 7293
rect 9214 7284 9220 7296
rect 9272 7324 9278 7336
rect 9674 7324 9680 7336
rect 9272 7296 9680 7324
rect 9272 7284 9278 7296
rect 9674 7284 9680 7296
rect 9732 7324 9738 7336
rect 10321 7327 10379 7333
rect 10321 7324 10333 7327
rect 9732 7296 10333 7324
rect 9732 7284 9738 7296
rect 10321 7293 10333 7296
rect 10367 7293 10379 7327
rect 10321 7287 10379 7293
rect 4154 7216 4160 7268
rect 4212 7256 4218 7268
rect 7653 7259 7711 7265
rect 7653 7256 7665 7259
rect 4212 7228 7665 7256
rect 4212 7216 4218 7228
rect 7653 7225 7665 7228
rect 7699 7225 7711 7259
rect 8478 7256 8484 7268
rect 7653 7219 7711 7225
rect 8128 7228 8484 7256
rect 1673 7191 1731 7197
rect 1673 7157 1685 7191
rect 1719 7188 1731 7191
rect 3418 7188 3424 7200
rect 1719 7160 3424 7188
rect 1719 7157 1731 7160
rect 1673 7151 1731 7157
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 3602 7188 3608 7200
rect 3563 7160 3608 7188
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 4706 7188 4712 7200
rect 4667 7160 4712 7188
rect 4706 7148 4712 7160
rect 4764 7188 4770 7200
rect 8128 7188 8156 7228
rect 8478 7216 8484 7228
rect 8536 7216 8542 7268
rect 8570 7216 8576 7268
rect 8628 7265 8634 7268
rect 8628 7259 8692 7265
rect 8628 7225 8646 7259
rect 8680 7225 8692 7259
rect 8628 7219 8692 7225
rect 8628 7216 8634 7219
rect 4764 7160 8156 7188
rect 4764 7148 4770 7160
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 10428 7188 10456 7364
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12894 7392 12900 7404
rect 12124 7364 12900 7392
rect 12124 7352 12130 7364
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13078 7352 13084 7404
rect 13136 7392 13142 7404
rect 13136 7364 13308 7392
rect 13136 7352 13142 7364
rect 10588 7327 10646 7333
rect 10588 7293 10600 7327
rect 10634 7324 10646 7327
rect 11054 7324 11060 7336
rect 10634 7296 11060 7324
rect 10634 7293 10646 7296
rect 10588 7287 10646 7293
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 13170 7324 13176 7336
rect 12851 7296 13176 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 11072 7256 11100 7284
rect 12897 7259 12955 7265
rect 11072 7228 12848 7256
rect 8260 7160 10456 7188
rect 8260 7148 8266 7160
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12820 7188 12848 7228
rect 12897 7225 12909 7259
rect 12943 7256 12955 7259
rect 12986 7256 12992 7268
rect 12943 7228 12992 7256
rect 12943 7225 12955 7228
rect 12897 7219 12955 7225
rect 12986 7216 12992 7228
rect 13044 7216 13050 7268
rect 13170 7188 13176 7200
rect 12492 7160 12537 7188
rect 12820 7160 13176 7188
rect 12492 7148 12498 7160
rect 13170 7148 13176 7160
rect 13228 7188 13234 7200
rect 13280 7188 13308 7364
rect 13228 7160 13308 7188
rect 13648 7188 13676 7432
rect 13740 7333 13768 7500
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 15102 7528 15108 7540
rect 15063 7500 15108 7528
rect 15102 7488 15108 7500
rect 15160 7488 15166 7540
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 15565 7327 15623 7333
rect 15565 7324 15577 7327
rect 13771 7296 15577 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 15565 7293 15577 7296
rect 15611 7293 15623 7327
rect 15565 7287 15623 7293
rect 13992 7259 14050 7265
rect 13992 7225 14004 7259
rect 14038 7256 14050 7259
rect 15832 7259 15890 7265
rect 14038 7228 15792 7256
rect 14038 7225 14050 7228
rect 13992 7219 14050 7225
rect 15010 7188 15016 7200
rect 13648 7160 15016 7188
rect 13228 7148 13234 7160
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15764 7188 15792 7228
rect 15832 7225 15844 7259
rect 15878 7256 15890 7259
rect 16114 7256 16120 7268
rect 15878 7228 16120 7256
rect 15878 7225 15890 7228
rect 15832 7219 15890 7225
rect 16114 7216 16120 7228
rect 16172 7216 16178 7268
rect 16482 7188 16488 7200
rect 15764 7160 16488 7188
rect 16482 7148 16488 7160
rect 16540 7188 16546 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 16540 7160 16957 7188
rect 16540 7148 16546 7160
rect 16945 7157 16957 7160
rect 16991 7157 17003 7191
rect 16945 7151 17003 7157
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 2777 6987 2835 6993
rect 2777 6953 2789 6987
rect 2823 6984 2835 6987
rect 4154 6984 4160 6996
rect 2823 6956 4160 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 4154 6944 4160 6956
rect 4212 6944 4218 6996
rect 4706 6944 4712 6996
rect 4764 6984 4770 6996
rect 4982 6984 4988 6996
rect 4764 6956 4988 6984
rect 4764 6944 4770 6956
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 5445 6987 5503 6993
rect 5445 6984 5457 6987
rect 5132 6956 5457 6984
rect 5132 6944 5138 6956
rect 5445 6953 5457 6956
rect 5491 6984 5503 6987
rect 5994 6984 6000 6996
rect 5491 6956 6000 6984
rect 5491 6953 5503 6956
rect 5445 6947 5503 6953
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 6365 6987 6423 6993
rect 6365 6953 6377 6987
rect 6411 6984 6423 6987
rect 7101 6987 7159 6993
rect 7101 6984 7113 6987
rect 6411 6956 7113 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 7101 6953 7113 6956
rect 7147 6953 7159 6987
rect 7101 6947 7159 6953
rect 7469 6987 7527 6993
rect 7469 6953 7481 6987
rect 7515 6984 7527 6987
rect 8110 6984 8116 6996
rect 7515 6956 8116 6984
rect 7515 6953 7527 6956
rect 7469 6947 7527 6953
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 11977 6987 12035 6993
rect 8220 6956 10824 6984
rect 3142 6916 3148 6928
rect 3103 6888 3148 6916
rect 3142 6876 3148 6888
rect 3200 6876 3206 6928
rect 3712 6888 4476 6916
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 3712 6848 3740 6888
rect 1719 6820 3740 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 4321 6851 4379 6857
rect 4321 6848 4333 6851
rect 3844 6820 4333 6848
rect 3844 6808 3850 6820
rect 4321 6817 4333 6820
rect 4367 6817 4379 6851
rect 4448 6848 4476 6888
rect 5902 6876 5908 6928
rect 5960 6916 5966 6928
rect 8220 6916 8248 6956
rect 5960 6888 8248 6916
rect 8757 6919 8815 6925
rect 5960 6876 5966 6888
rect 8757 6885 8769 6919
rect 8803 6916 8815 6919
rect 9490 6916 9496 6928
rect 8803 6888 9496 6916
rect 8803 6885 8815 6888
rect 8757 6879 8815 6885
rect 9490 6876 9496 6888
rect 9548 6876 9554 6928
rect 10796 6925 10824 6956
rect 11977 6953 11989 6987
rect 12023 6984 12035 6987
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 12023 6956 12817 6984
rect 12023 6953 12035 6956
rect 11977 6947 12035 6953
rect 12805 6953 12817 6956
rect 12851 6953 12863 6987
rect 12805 6947 12863 6953
rect 13173 6987 13231 6993
rect 13173 6953 13185 6987
rect 13219 6984 13231 6987
rect 13630 6984 13636 6996
rect 13219 6956 13636 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 14369 6987 14427 6993
rect 14369 6984 14381 6987
rect 14148 6956 14381 6984
rect 14148 6944 14154 6956
rect 14369 6953 14381 6956
rect 14415 6953 14427 6987
rect 15654 6984 15660 6996
rect 15615 6956 15660 6984
rect 14369 6947 14427 6953
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 16574 6944 16580 6996
rect 16632 6984 16638 6996
rect 17037 6987 17095 6993
rect 17037 6984 17049 6987
rect 16632 6956 17049 6984
rect 16632 6944 16638 6956
rect 17037 6953 17049 6956
rect 17083 6953 17095 6987
rect 17037 6947 17095 6953
rect 10781 6919 10839 6925
rect 10781 6885 10793 6919
rect 10827 6916 10839 6919
rect 16592 6916 16620 6944
rect 10827 6888 16620 6916
rect 10827 6885 10839 6888
rect 10781 6879 10839 6885
rect 16850 6876 16856 6928
rect 16908 6916 16914 6928
rect 17129 6919 17187 6925
rect 17129 6916 17141 6919
rect 16908 6888 17141 6916
rect 16908 6876 16914 6888
rect 17129 6885 17141 6888
rect 17175 6885 17187 6919
rect 17129 6879 17187 6885
rect 5810 6848 5816 6860
rect 4448 6820 5816 6848
rect 4321 6811 4379 6817
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 6270 6848 6276 6860
rect 6231 6820 6276 6848
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 7561 6851 7619 6857
rect 7561 6817 7573 6851
rect 7607 6848 7619 6851
rect 8018 6848 8024 6860
rect 7607 6820 8024 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 8018 6808 8024 6820
rect 8076 6848 8082 6860
rect 9677 6851 9735 6857
rect 8076 6820 9168 6848
rect 8076 6808 8082 6820
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 3237 6783 3295 6789
rect 3237 6780 3249 6783
rect 3108 6752 3249 6780
rect 3108 6740 3114 6752
rect 3237 6749 3249 6752
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3878 6780 3884 6792
rect 3467 6752 3884 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 6549 6783 6607 6789
rect 6549 6780 6561 6783
rect 4065 6743 4123 6749
rect 6472 6752 6561 6780
rect 2406 6672 2412 6724
rect 2464 6712 2470 6724
rect 4080 6712 4108 6743
rect 2464 6684 4108 6712
rect 2464 6672 2470 6684
rect 1857 6647 1915 6653
rect 1857 6613 1869 6647
rect 1903 6644 1915 6647
rect 2958 6644 2964 6656
rect 1903 6616 2964 6644
rect 1903 6613 1915 6616
rect 1857 6607 1915 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 4080 6644 4108 6684
rect 4246 6644 4252 6656
rect 4080 6616 4252 6644
rect 4246 6604 4252 6616
rect 4304 6644 4310 6656
rect 5442 6644 5448 6656
rect 4304 6616 5448 6644
rect 4304 6604 4310 6616
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5902 6644 5908 6656
rect 5863 6616 5908 6644
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 6472 6644 6500 6752
rect 6549 6749 6561 6752
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 8846 6780 8852 6792
rect 7708 6752 7753 6780
rect 8807 6752 8852 6780
rect 7708 6740 7714 6752
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 8938 6740 8944 6792
rect 8996 6780 9002 6792
rect 9140 6780 9168 6820
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 10502 6848 10508 6860
rect 9723 6820 10508 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 10873 6851 10931 6857
rect 10873 6817 10885 6851
rect 10919 6848 10931 6851
rect 11514 6848 11520 6860
rect 10919 6820 11520 6848
rect 10919 6817 10931 6820
rect 10873 6811 10931 6817
rect 11514 6808 11520 6820
rect 11572 6848 11578 6860
rect 12069 6851 12127 6857
rect 11572 6820 12020 6848
rect 11572 6808 11578 6820
rect 10686 6780 10692 6792
rect 8996 6752 9041 6780
rect 9140 6752 10692 6780
rect 8996 6740 9002 6752
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 10962 6740 10968 6792
rect 11020 6780 11026 6792
rect 11992 6780 12020 6820
rect 12069 6817 12081 6851
rect 12115 6848 12127 6851
rect 12434 6848 12440 6860
rect 12115 6820 12440 6848
rect 12115 6817 12127 6820
rect 12069 6811 12127 6817
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 13170 6808 13176 6860
rect 13228 6848 13234 6860
rect 16868 6848 16896 6876
rect 13228 6820 13400 6848
rect 13228 6808 13234 6820
rect 12250 6780 12256 6792
rect 11020 6752 11065 6780
rect 11992 6752 12112 6780
rect 12211 6752 12256 6780
rect 11020 6740 11026 6752
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 10410 6712 10416 6724
rect 8168 6684 10272 6712
rect 10371 6684 10416 6712
rect 8168 6672 8174 6684
rect 6052 6616 6500 6644
rect 8389 6647 8447 6653
rect 6052 6604 6058 6616
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8478 6644 8484 6656
rect 8435 6616 8484 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 9861 6647 9919 6653
rect 9861 6644 9873 6647
rect 9732 6616 9873 6644
rect 9732 6604 9738 6616
rect 9861 6613 9873 6616
rect 9907 6613 9919 6647
rect 10244 6644 10272 6684
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 12084 6712 12112 6752
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13372 6789 13400 6820
rect 13648 6820 16896 6848
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 13136 6752 13277 6780
rect 13136 6740 13142 6752
rect 13265 6749 13277 6752
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 13648 6712 13676 6820
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 17460 6820 17877 6848
rect 17460 6808 17466 6820
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 13872 6752 14473 6780
rect 13872 6740 13878 6752
rect 14461 6749 14473 6752
rect 14507 6749 14519 6783
rect 14642 6780 14648 6792
rect 14603 6752 14648 6780
rect 14461 6743 14519 6749
rect 14642 6740 14648 6752
rect 14700 6740 14706 6792
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 15528 6752 15761 6780
rect 15528 6740 15534 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 11440 6684 12020 6712
rect 12084 6684 13676 6712
rect 13832 6684 14136 6712
rect 11440 6644 11468 6684
rect 10244 6616 11468 6644
rect 9861 6607 9919 6613
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 11609 6647 11667 6653
rect 11609 6644 11621 6647
rect 11572 6616 11621 6644
rect 11572 6604 11578 6616
rect 11609 6613 11621 6616
rect 11655 6613 11667 6647
rect 11992 6644 12020 6684
rect 13832 6644 13860 6684
rect 13998 6644 14004 6656
rect 11992 6616 13860 6644
rect 13959 6616 14004 6644
rect 11609 6607 11667 6613
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 14108 6644 14136 6684
rect 15102 6672 15108 6724
rect 15160 6712 15166 6724
rect 15856 6712 15884 6743
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17276 6752 17321 6780
rect 17276 6740 17282 6752
rect 16666 6712 16672 6724
rect 15160 6684 15884 6712
rect 16627 6684 16672 6712
rect 15160 6672 15166 6684
rect 16666 6672 16672 6684
rect 16724 6672 16730 6724
rect 15289 6647 15347 6653
rect 15289 6644 15301 6647
rect 14108 6616 15301 6644
rect 15289 6613 15301 6616
rect 15335 6613 15347 6647
rect 15289 6607 15347 6613
rect 18049 6647 18107 6653
rect 18049 6613 18061 6647
rect 18095 6644 18107 6647
rect 18969 6647 19027 6653
rect 18969 6644 18981 6647
rect 18095 6616 18981 6644
rect 18095 6613 18107 6616
rect 18049 6607 18107 6613
rect 18969 6613 18981 6616
rect 19015 6613 19027 6647
rect 18969 6607 19027 6613
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 3786 6440 3792 6452
rect 1688 6412 3648 6440
rect 3747 6412 3792 6440
rect 1688 6245 1716 6412
rect 2406 6304 2412 6316
rect 2367 6276 2412 6304
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 3620 6304 3648 6412
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 5258 6400 5264 6452
rect 5316 6440 5322 6452
rect 5316 6412 5580 6440
rect 5316 6400 5322 6412
rect 5552 6372 5580 6412
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 6328 6412 6837 6440
rect 6328 6400 6334 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 7800 6412 8033 6440
rect 7800 6400 7806 6412
rect 8021 6409 8033 6412
rect 8067 6409 8079 6443
rect 8021 6403 8079 6409
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 11149 6443 11207 6449
rect 11149 6440 11161 6443
rect 8352 6412 11161 6440
rect 8352 6400 8358 6412
rect 11149 6409 11161 6412
rect 11195 6409 11207 6443
rect 11149 6403 11207 6409
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 12710 6440 12716 6452
rect 12216 6412 12716 6440
rect 12216 6400 12222 6412
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 14734 6440 14740 6452
rect 13924 6412 14740 6440
rect 5552 6344 6684 6372
rect 4430 6304 4436 6316
rect 3620 6276 4436 6304
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6205 1731 6239
rect 1673 6199 1731 6205
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 4617 6239 4675 6245
rect 4617 6236 4629 6239
rect 4304 6208 4629 6236
rect 4304 6196 4310 6208
rect 4617 6205 4629 6208
rect 4663 6205 4675 6239
rect 4617 6199 4675 6205
rect 4706 6196 4712 6248
rect 4764 6236 4770 6248
rect 4884 6239 4942 6245
rect 4884 6236 4896 6239
rect 4764 6208 4896 6236
rect 4764 6196 4770 6208
rect 4884 6205 4896 6208
rect 4930 6236 4942 6239
rect 6270 6236 6276 6248
rect 4930 6208 6276 6236
rect 4930 6205 4942 6208
rect 4884 6199 4942 6205
rect 6270 6196 6276 6208
rect 6328 6196 6334 6248
rect 6656 6245 6684 6344
rect 10962 6332 10968 6384
rect 11020 6372 11026 6384
rect 13630 6372 13636 6384
rect 11020 6344 13636 6372
rect 11020 6332 11026 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 6840 6276 7481 6304
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 2590 6128 2596 6180
rect 2648 6177 2654 6180
rect 2648 6171 2712 6177
rect 2648 6137 2666 6171
rect 2700 6137 2712 6171
rect 2648 6131 2712 6137
rect 2648 6128 2654 6131
rect 1854 6100 1860 6112
rect 1815 6072 1860 6100
rect 1854 6060 1860 6072
rect 1912 6060 1918 6112
rect 5994 6060 6000 6112
rect 6052 6100 6058 6112
rect 6052 6072 6097 6100
rect 6052 6060 6058 6072
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 6236 6072 6469 6100
rect 6236 6060 6242 6072
rect 6457 6069 6469 6072
rect 6503 6069 6515 6103
rect 6457 6063 6515 6069
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 6840 6100 6868 6276
rect 7469 6273 7481 6276
rect 7515 6304 7527 6307
rect 7650 6304 7656 6316
rect 7515 6276 7656 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 8478 6304 8484 6316
rect 8439 6276 8484 6304
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 9214 6304 9220 6316
rect 8628 6276 8673 6304
rect 9175 6276 9220 6304
rect 8628 6264 8634 6276
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 11606 6304 11612 6316
rect 11567 6276 11612 6304
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 11790 6304 11796 6316
rect 11751 6276 11796 6304
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 11882 6264 11888 6316
rect 11940 6304 11946 6316
rect 12529 6307 12587 6313
rect 12529 6304 12541 6307
rect 11940 6276 12541 6304
rect 11940 6264 11946 6276
rect 12529 6273 12541 6276
rect 12575 6273 12587 6307
rect 12529 6267 12587 6273
rect 13541 6307 13599 6313
rect 13541 6273 13553 6307
rect 13587 6304 13599 6307
rect 13924 6304 13952 6412
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 15933 6443 15991 6449
rect 15933 6440 15945 6443
rect 15712 6412 15945 6440
rect 15712 6400 15718 6412
rect 15933 6409 15945 6412
rect 15979 6409 15991 6443
rect 15933 6403 15991 6409
rect 15473 6375 15531 6381
rect 15473 6341 15485 6375
rect 15519 6372 15531 6375
rect 16114 6372 16120 6384
rect 15519 6344 16120 6372
rect 15519 6341 15531 6344
rect 15473 6335 15531 6341
rect 16114 6332 16120 6344
rect 16172 6332 16178 6384
rect 17126 6332 17132 6384
rect 17184 6332 17190 6384
rect 13587 6276 13952 6304
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 13998 6264 14004 6316
rect 14056 6304 14062 6316
rect 16482 6304 16488 6316
rect 14056 6276 14228 6304
rect 16443 6276 16488 6304
rect 14056 6264 14062 6276
rect 7193 6239 7251 6245
rect 7193 6205 7205 6239
rect 7239 6236 7251 6239
rect 8754 6236 8760 6248
rect 7239 6208 8760 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 9484 6239 9542 6245
rect 9484 6205 9496 6239
rect 9530 6236 9542 6239
rect 10318 6236 10324 6248
rect 9530 6208 10324 6236
rect 9530 6205 9542 6208
rect 9484 6199 9542 6205
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 11514 6236 11520 6248
rect 11475 6208 11520 6236
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 14090 6236 14096 6248
rect 14051 6208 14096 6236
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 14200 6236 14228 6276
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 16850 6264 16856 6316
rect 16908 6304 16914 6316
rect 17034 6304 17040 6316
rect 16908 6276 17040 6304
rect 16908 6264 16914 6276
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 17144 6304 17172 6332
rect 17144 6276 17264 6304
rect 17126 6236 17132 6248
rect 14200 6208 17132 6236
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 17236 6245 17264 6276
rect 17221 6239 17279 6245
rect 17221 6205 17233 6239
rect 17267 6205 17279 6239
rect 17221 6199 17279 6205
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 7432 6140 8524 6168
rect 7432 6128 7438 6140
rect 7282 6100 7288 6112
rect 6788 6072 6868 6100
rect 7243 6072 7288 6100
rect 6788 6060 6794 6072
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 8386 6100 8392 6112
rect 8347 6072 8392 6100
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8496 6100 8524 6140
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 12621 6171 12679 6177
rect 12621 6168 12633 6171
rect 9180 6140 12633 6168
rect 9180 6128 9186 6140
rect 12621 6137 12633 6140
rect 12667 6168 12679 6171
rect 13170 6168 13176 6180
rect 12667 6140 13176 6168
rect 12667 6137 12679 6140
rect 12621 6131 12679 6137
rect 13170 6128 13176 6140
rect 13228 6128 13234 6180
rect 14360 6171 14418 6177
rect 14360 6137 14372 6171
rect 14406 6168 14418 6171
rect 14642 6168 14648 6180
rect 14406 6140 14648 6168
rect 14406 6137 14418 6140
rect 14360 6131 14418 6137
rect 14642 6128 14648 6140
rect 14700 6168 14706 6180
rect 15194 6168 15200 6180
rect 14700 6140 15200 6168
rect 14700 6128 14706 6140
rect 15194 6128 15200 6140
rect 15252 6128 15258 6180
rect 16301 6171 16359 6177
rect 16301 6137 16313 6171
rect 16347 6168 16359 6171
rect 16666 6168 16672 6180
rect 16347 6140 16672 6168
rect 16347 6137 16359 6140
rect 16301 6131 16359 6137
rect 16666 6128 16672 6140
rect 16724 6128 16730 6180
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 8496 6072 10609 6100
rect 10597 6069 10609 6072
rect 10643 6069 10655 6103
rect 10597 6063 10655 6069
rect 16393 6103 16451 6109
rect 16393 6069 16405 6103
rect 16439 6100 16451 6103
rect 17310 6100 17316 6112
rect 16439 6072 17316 6100
rect 16439 6069 16451 6072
rect 16393 6063 16451 6069
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 17402 6060 17408 6112
rect 17460 6100 17466 6112
rect 17460 6072 17505 6100
rect 17460 6060 17466 6072
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3283 5868 4077 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 5626 5896 5632 5908
rect 4488 5868 5632 5896
rect 4488 5856 4494 5868
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 6730 5896 6736 5908
rect 6328 5868 6736 5896
rect 6328 5856 6334 5868
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 7340 5868 9260 5896
rect 7340 5856 7346 5868
rect 3145 5831 3203 5837
rect 3145 5797 3157 5831
rect 3191 5828 3203 5831
rect 5902 5828 5908 5840
rect 3191 5800 4108 5828
rect 3191 5797 3203 5800
rect 3145 5791 3203 5797
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 1688 5624 1716 5723
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1820 5664 1869 5692
rect 1820 5652 1826 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 3786 5692 3792 5704
rect 3467 5664 3792 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4080 5692 4108 5800
rect 4264 5800 5908 5828
rect 4264 5692 4292 5800
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 6540 5831 6598 5837
rect 6540 5797 6552 5831
rect 6586 5828 6598 5831
rect 7374 5828 7380 5840
rect 6586 5800 7380 5828
rect 6586 5797 6598 5800
rect 6540 5791 6598 5797
rect 7374 5788 7380 5800
rect 7432 5788 7438 5840
rect 9122 5828 9128 5840
rect 8312 5800 9128 5828
rect 4430 5760 4436 5772
rect 4391 5732 4436 5760
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5760 5595 5763
rect 8312 5760 8340 5800
rect 9122 5788 9128 5800
rect 9180 5788 9186 5840
rect 9232 5828 9260 5868
rect 9306 5856 9312 5908
rect 9364 5896 9370 5908
rect 10962 5896 10968 5908
rect 9364 5868 10968 5896
rect 9364 5856 9370 5868
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 11790 5856 11796 5908
rect 11848 5896 11854 5908
rect 12897 5899 12955 5905
rect 12897 5896 12909 5899
rect 11848 5868 12909 5896
rect 11848 5856 11854 5868
rect 12897 5865 12909 5868
rect 12943 5896 12955 5899
rect 16485 5899 16543 5905
rect 12943 5868 13216 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 12158 5828 12164 5840
rect 9232 5800 12164 5828
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 13188 5828 13216 5868
rect 16485 5865 16497 5899
rect 16531 5896 16543 5899
rect 16758 5896 16764 5908
rect 16531 5868 16764 5896
rect 16531 5865 16543 5868
rect 16485 5859 16543 5865
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 17310 5896 17316 5908
rect 17271 5868 17316 5896
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 17678 5896 17684 5908
rect 17639 5868 17684 5896
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 13602 5831 13660 5837
rect 13602 5828 13614 5831
rect 13188 5800 13614 5828
rect 13602 5797 13614 5800
rect 13648 5797 13660 5831
rect 13602 5791 13660 5797
rect 16114 5788 16120 5840
rect 16172 5828 16178 5840
rect 16172 5800 16620 5828
rect 16172 5788 16178 5800
rect 5583 5732 8340 5760
rect 8757 5763 8815 5769
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 8757 5729 8769 5763
rect 8803 5760 8815 5763
rect 9490 5760 9496 5772
rect 8803 5732 9496 5760
rect 8803 5729 8815 5732
rect 8757 5723 8815 5729
rect 9490 5720 9496 5732
rect 9548 5760 9554 5772
rect 9933 5763 9991 5769
rect 9933 5760 9945 5763
rect 9548 5732 9945 5760
rect 9548 5720 9554 5732
rect 9933 5729 9945 5732
rect 9979 5729 9991 5763
rect 9933 5723 9991 5729
rect 11784 5763 11842 5769
rect 11784 5729 11796 5763
rect 11830 5760 11842 5763
rect 12250 5760 12256 5772
rect 11830 5732 12256 5760
rect 11830 5729 11842 5732
rect 11784 5723 11842 5729
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 13357 5763 13415 5769
rect 13357 5729 13369 5763
rect 13403 5760 13415 5763
rect 14090 5760 14096 5772
rect 13403 5732 14096 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 4080 5664 4292 5692
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 2777 5627 2835 5633
rect 2777 5624 2789 5627
rect 1688 5596 2789 5624
rect 2777 5593 2789 5596
rect 2823 5593 2835 5627
rect 2777 5587 2835 5593
rect 3786 5516 3792 5568
rect 3844 5556 3850 5568
rect 4540 5556 4568 5655
rect 4614 5652 4620 5704
rect 4672 5692 4678 5704
rect 4672 5664 4717 5692
rect 4672 5652 4678 5664
rect 6178 5652 6184 5704
rect 6236 5692 6242 5704
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 6236 5664 6285 5692
rect 6236 5652 6242 5664
rect 6273 5661 6285 5664
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 9030 5692 9036 5704
rect 8435 5664 9036 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9214 5652 9220 5704
rect 9272 5692 9278 5704
rect 9582 5692 9588 5704
rect 9272 5664 9588 5692
rect 9272 5652 9278 5664
rect 9582 5652 9588 5664
rect 9640 5692 9646 5704
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9640 5664 9689 5692
rect 9640 5652 9646 5664
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 10962 5652 10968 5704
rect 11020 5692 11026 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11020 5664 11529 5692
rect 11020 5652 11026 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 7392 5596 8340 5624
rect 3844 5528 4568 5556
rect 5721 5559 5779 5565
rect 3844 5516 3850 5528
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 7392 5556 7420 5596
rect 7650 5556 7656 5568
rect 5767 5528 7420 5556
rect 7611 5528 7656 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 8312 5556 8340 5596
rect 8478 5584 8484 5636
rect 8536 5624 8542 5636
rect 9306 5624 9312 5636
rect 8536 5596 9312 5624
rect 8536 5584 8542 5596
rect 9306 5584 9312 5596
rect 9364 5584 9370 5636
rect 9122 5556 9128 5568
rect 8312 5528 9128 5556
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 10468 5528 11069 5556
rect 10468 5516 10474 5528
rect 11057 5525 11069 5528
rect 11103 5525 11115 5559
rect 11532 5556 11560 5655
rect 13372 5556 13400 5723
rect 14090 5720 14096 5732
rect 14148 5720 14154 5772
rect 15381 5763 15439 5769
rect 15381 5729 15393 5763
rect 15427 5760 15439 5763
rect 15654 5760 15660 5772
rect 15427 5732 15660 5760
rect 15427 5729 15439 5732
rect 15381 5723 15439 5729
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 16592 5760 16620 5800
rect 17494 5788 17500 5840
rect 17552 5828 17558 5840
rect 17773 5831 17831 5837
rect 17773 5828 17785 5831
rect 17552 5800 17785 5828
rect 17552 5788 17558 5800
rect 17773 5797 17785 5800
rect 17819 5828 17831 5831
rect 18322 5828 18328 5840
rect 17819 5800 18328 5828
rect 17819 5797 17831 5800
rect 17773 5791 17831 5797
rect 18322 5788 18328 5800
rect 18380 5788 18386 5840
rect 16592 5732 16712 5760
rect 16574 5692 16580 5704
rect 16535 5664 16580 5692
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 16684 5701 16712 5732
rect 16669 5695 16727 5701
rect 16669 5661 16681 5695
rect 16715 5692 16727 5695
rect 17034 5692 17040 5704
rect 16715 5664 17040 5692
rect 16715 5661 16727 5664
rect 16669 5655 16727 5661
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 17865 5695 17923 5701
rect 17865 5661 17877 5695
rect 17911 5661 17923 5695
rect 18966 5692 18972 5704
rect 18927 5664 18972 5692
rect 17865 5655 17923 5661
rect 17052 5624 17080 5652
rect 17880 5624 17908 5655
rect 18966 5652 18972 5664
rect 19024 5652 19030 5704
rect 17052 5596 17908 5624
rect 11532 5528 13400 5556
rect 14737 5559 14795 5565
rect 11057 5519 11115 5525
rect 14737 5525 14749 5559
rect 14783 5556 14795 5559
rect 15194 5556 15200 5568
rect 14783 5528 15200 5556
rect 14783 5525 14795 5528
rect 14737 5519 14795 5525
rect 15194 5516 15200 5528
rect 15252 5516 15258 5568
rect 15565 5559 15623 5565
rect 15565 5525 15577 5559
rect 15611 5556 15623 5559
rect 15654 5556 15660 5568
rect 15611 5528 15660 5556
rect 15611 5525 15623 5528
rect 15565 5519 15623 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 16114 5556 16120 5568
rect 16075 5528 16120 5556
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 1854 5352 1860 5364
rect 1815 5324 1860 5352
rect 1854 5312 1860 5324
rect 1912 5312 1918 5364
rect 3697 5355 3755 5361
rect 3697 5321 3709 5355
rect 3743 5352 3755 5355
rect 4430 5352 4436 5364
rect 3743 5324 4436 5352
rect 3743 5321 3755 5324
rect 3697 5315 3755 5321
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 8294 5352 8300 5364
rect 4908 5324 8300 5352
rect 4908 5284 4936 5324
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 9490 5352 9496 5364
rect 9451 5324 9496 5352
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 9582 5312 9588 5364
rect 9640 5352 9646 5364
rect 9953 5355 10011 5361
rect 9953 5352 9965 5355
rect 9640 5324 9965 5352
rect 9640 5312 9646 5324
rect 9953 5321 9965 5324
rect 9999 5321 10011 5355
rect 11698 5352 11704 5364
rect 9953 5315 10011 5321
rect 10152 5324 11704 5352
rect 6270 5284 6276 5296
rect 2608 5256 4936 5284
rect 6231 5256 6276 5284
rect 1670 5148 1676 5160
rect 1631 5120 1676 5148
rect 1670 5108 1676 5120
rect 1728 5108 1734 5160
rect 2608 5157 2636 5256
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 6362 5244 6368 5296
rect 6420 5284 6426 5296
rect 7285 5287 7343 5293
rect 7285 5284 7297 5287
rect 6420 5256 7297 5284
rect 6420 5244 6426 5256
rect 7285 5253 7297 5256
rect 7331 5253 7343 5287
rect 7285 5247 7343 5253
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 3234 5216 3240 5228
rect 2924 5188 3240 5216
rect 2924 5176 2930 5188
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4706 5216 4712 5228
rect 4387 5188 4712 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 7300 5216 7328 5247
rect 7300 5188 8248 5216
rect 2593 5151 2651 5157
rect 2593 5117 2605 5151
rect 2639 5117 2651 5151
rect 2593 5111 2651 5117
rect 3326 5108 3332 5160
rect 3384 5148 3390 5160
rect 4065 5151 4123 5157
rect 4065 5148 4077 5151
rect 3384 5120 4077 5148
rect 3384 5108 3390 5120
rect 4065 5117 4077 5120
rect 4111 5117 4123 5151
rect 4065 5111 4123 5117
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 4304 5120 4905 5148
rect 4304 5108 4310 5120
rect 4893 5117 4905 5120
rect 4939 5148 4951 5151
rect 6178 5148 6184 5160
rect 4939 5120 6184 5148
rect 4939 5117 4951 5120
rect 4893 5111 4951 5117
rect 6178 5108 6184 5120
rect 6236 5108 6242 5160
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6788 5120 6837 5148
rect 6788 5108 6794 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5148 7251 5151
rect 7374 5148 7380 5160
rect 7239 5120 7380 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 7742 5108 7748 5160
rect 7800 5148 7806 5160
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 7800 5120 8125 5148
rect 7800 5108 7806 5120
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8220 5148 8248 5188
rect 9858 5148 9864 5160
rect 8220 5120 9864 5148
rect 8113 5111 8171 5117
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 2866 5080 2872 5092
rect 2827 5052 2872 5080
rect 2866 5040 2872 5052
rect 2924 5040 2930 5092
rect 5074 5040 5080 5092
rect 5132 5089 5138 5092
rect 5132 5083 5196 5089
rect 5132 5049 5150 5083
rect 5184 5049 5196 5083
rect 5132 5043 5196 5049
rect 8380 5083 8438 5089
rect 8380 5049 8392 5083
rect 8426 5080 8438 5083
rect 9030 5080 9036 5092
rect 8426 5052 9036 5080
rect 8426 5049 8438 5052
rect 8380 5043 8438 5049
rect 5132 5040 5138 5043
rect 9030 5040 9036 5052
rect 9088 5040 9094 5092
rect 9968 5080 9996 5315
rect 10152 5157 10180 5324
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 13538 5312 13544 5364
rect 13596 5352 13602 5364
rect 13814 5352 13820 5364
rect 13596 5324 13820 5352
rect 13596 5312 13602 5324
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 15470 5352 15476 5364
rect 15431 5324 15476 5352
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 16666 5352 16672 5364
rect 16627 5324 16672 5352
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 12713 5287 12771 5293
rect 12713 5253 12725 5287
rect 12759 5284 12771 5287
rect 16298 5284 16304 5296
rect 12759 5256 16304 5284
rect 12759 5253 12771 5256
rect 12713 5247 12771 5253
rect 16298 5244 16304 5256
rect 16356 5244 16362 5296
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5216 13415 5219
rect 13630 5216 13636 5228
rect 13403 5188 13636 5216
rect 13403 5185 13415 5188
rect 13357 5179 13415 5185
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 14182 5216 14188 5228
rect 14143 5188 14188 5216
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5216 16083 5219
rect 16482 5216 16488 5228
rect 16071 5188 16488 5216
rect 16071 5185 16083 5188
rect 16025 5179 16083 5185
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 17034 5176 17040 5228
rect 17092 5216 17098 5228
rect 17221 5219 17279 5225
rect 17221 5216 17233 5219
rect 17092 5188 17233 5216
rect 17092 5176 17098 5188
rect 17221 5185 17233 5188
rect 17267 5185 17279 5219
rect 17221 5179 17279 5185
rect 10137 5151 10195 5157
rect 10137 5117 10149 5151
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 10229 5151 10287 5157
rect 10229 5117 10241 5151
rect 10275 5148 10287 5151
rect 10962 5148 10968 5160
rect 10275 5120 10968 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 10244 5080 10272 5111
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 12529 5151 12587 5157
rect 12529 5117 12541 5151
rect 12575 5148 12587 5151
rect 12710 5148 12716 5160
rect 12575 5120 12716 5148
rect 12575 5117 12587 5120
rect 12529 5111 12587 5117
rect 12710 5108 12716 5120
rect 12768 5108 12774 5160
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 16114 5148 16120 5160
rect 15887 5120 16120 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 16114 5108 16120 5120
rect 16172 5108 16178 5160
rect 17129 5151 17187 5157
rect 17129 5117 17141 5151
rect 17175 5148 17187 5151
rect 17310 5148 17316 5160
rect 17175 5120 17316 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 17310 5108 17316 5120
rect 17368 5108 17374 5160
rect 9968 5052 10272 5080
rect 10410 5040 10416 5092
rect 10468 5089 10474 5092
rect 10468 5083 10532 5089
rect 10468 5049 10486 5083
rect 10520 5049 10532 5083
rect 10468 5043 10532 5049
rect 10468 5040 10474 5043
rect 11146 5040 11152 5092
rect 11204 5080 11210 5092
rect 11698 5080 11704 5092
rect 11204 5052 11704 5080
rect 11204 5040 11210 5052
rect 11698 5040 11704 5052
rect 11756 5040 11762 5092
rect 13354 5040 13360 5092
rect 13412 5080 13418 5092
rect 13449 5083 13507 5089
rect 13449 5080 13461 5083
rect 13412 5052 13461 5080
rect 13412 5040 13418 5052
rect 13449 5049 13461 5052
rect 13495 5049 13507 5083
rect 13449 5043 13507 5049
rect 14829 5083 14887 5089
rect 14829 5049 14841 5083
rect 14875 5080 14887 5083
rect 17037 5083 17095 5089
rect 17037 5080 17049 5083
rect 14875 5052 17049 5080
rect 14875 5049 14887 5052
rect 14829 5043 14887 5049
rect 17037 5049 17049 5052
rect 17083 5049 17095 5083
rect 17037 5043 17095 5049
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 5012 4215 5015
rect 5626 5012 5632 5024
rect 4203 4984 5632 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 9398 5012 9404 5024
rect 6052 4984 9404 5012
rect 6052 4972 6058 4984
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 10836 4984 11621 5012
rect 10836 4972 10842 4984
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 15930 5012 15936 5024
rect 15891 4984 15936 5012
rect 11609 4975 11667 4981
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 1854 4808 1860 4820
rect 1815 4780 1860 4808
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2593 4811 2651 4817
rect 2593 4777 2605 4811
rect 2639 4808 2651 4811
rect 2774 4808 2780 4820
rect 2639 4780 2780 4808
rect 2639 4777 2651 4780
rect 2593 4771 2651 4777
rect 2774 4768 2780 4780
rect 2832 4768 2838 4820
rect 4798 4768 4804 4820
rect 4856 4768 4862 4820
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4808 4951 4811
rect 5350 4808 5356 4820
rect 4939 4780 5356 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 5626 4808 5632 4820
rect 5587 4780 5632 4808
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 8846 4808 8852 4820
rect 5920 4780 8852 4808
rect 3234 4740 3240 4752
rect 1688 4712 3240 4740
rect 1688 4681 1716 4712
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 4816 4740 4844 4768
rect 4816 4712 5396 4740
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4641 1731 4675
rect 2406 4672 2412 4684
rect 2367 4644 2412 4672
rect 1673 4635 1731 4641
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4672 3203 4675
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 3191 4644 4813 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 4801 4641 4813 4644
rect 4847 4672 4859 4675
rect 5166 4672 5172 4684
rect 4847 4644 5172 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5074 4604 5080 4616
rect 5035 4576 5080 4604
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5368 4604 5396 4712
rect 5920 4604 5948 4780
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 9030 4808 9036 4820
rect 8991 4780 9036 4808
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 11112 4780 15608 4808
rect 11112 4768 11118 4780
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 11146 4740 11152 4752
rect 6052 4712 6097 4740
rect 6932 4712 11152 4740
rect 6052 4700 6058 4712
rect 6932 4681 6960 4712
rect 11146 4700 11152 4712
rect 11204 4700 11210 4752
rect 11974 4740 11980 4752
rect 11935 4712 11980 4740
rect 11974 4700 11980 4712
rect 12032 4700 12038 4752
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 12124 4712 12169 4740
rect 12124 4700 12130 4712
rect 12434 4700 12440 4752
rect 12492 4740 12498 4752
rect 13725 4743 13783 4749
rect 13725 4740 13737 4743
rect 12492 4712 13737 4740
rect 12492 4700 12498 4712
rect 13725 4709 13737 4712
rect 13771 4709 13783 4743
rect 13725 4703 13783 4709
rect 13814 4700 13820 4752
rect 13872 4740 13878 4752
rect 13872 4712 13917 4740
rect 13872 4700 13878 4712
rect 15102 4700 15108 4752
rect 15160 4740 15166 4752
rect 15473 4743 15531 4749
rect 15473 4740 15485 4743
rect 15160 4712 15485 4740
rect 15160 4700 15166 4712
rect 15473 4709 15485 4712
rect 15519 4709 15531 4743
rect 15580 4740 15608 4780
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 16853 4811 16911 4817
rect 16853 4808 16865 4811
rect 15988 4780 16865 4808
rect 15988 4768 15994 4780
rect 16853 4777 16865 4780
rect 16899 4777 16911 4811
rect 16853 4771 16911 4777
rect 17126 4768 17132 4820
rect 17184 4808 17190 4820
rect 17221 4811 17279 4817
rect 17221 4808 17233 4811
rect 17184 4780 17233 4808
rect 17184 4768 17190 4780
rect 17221 4777 17233 4780
rect 17267 4777 17279 4811
rect 17221 4771 17279 4777
rect 16390 4740 16396 4752
rect 15580 4712 16252 4740
rect 16351 4712 16396 4740
rect 15473 4703 15531 4709
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4641 6975 4675
rect 7742 4672 7748 4684
rect 6917 4635 6975 4641
rect 7668 4644 7748 4672
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 5368 4576 6101 4604
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 5092 4536 5120 4564
rect 5442 4536 5448 4548
rect 5092 4508 5448 4536
rect 5442 4496 5448 4508
rect 5500 4536 5506 4548
rect 6196 4536 6224 4567
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 7668 4613 7696 4644
rect 7742 4632 7748 4644
rect 7800 4632 7806 4684
rect 7920 4675 7978 4681
rect 7920 4641 7932 4675
rect 7966 4672 7978 4675
rect 8478 4672 8484 4684
rect 7966 4644 8484 4672
rect 7966 4641 7978 4644
rect 7920 4635 7978 4641
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 8904 4644 9689 4672
rect 8904 4632 8910 4644
rect 9677 4641 9689 4644
rect 9723 4641 9735 4675
rect 10778 4672 10784 4684
rect 10739 4644 10784 4672
rect 9677 4635 9735 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 16224 4672 16252 4712
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 16758 4672 16764 4684
rect 16224 4644 16764 4672
rect 16758 4632 16764 4644
rect 16816 4632 16822 4684
rect 17034 4632 17040 4684
rect 17092 4672 17098 4684
rect 17092 4644 17448 4672
rect 17092 4632 17098 4644
rect 7653 4607 7711 4613
rect 7653 4604 7665 4607
rect 6328 4576 7665 4604
rect 6328 4564 6334 4576
rect 7653 4573 7665 4576
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 9858 4564 9864 4616
rect 9916 4604 9922 4616
rect 10502 4604 10508 4616
rect 9916 4576 10508 4604
rect 9916 4564 9922 4576
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4573 13047 4607
rect 14366 4604 14372 4616
rect 14327 4576 14372 4604
rect 12989 4567 13047 4573
rect 5500 4508 6224 4536
rect 5500 4496 5506 4508
rect 8938 4496 8944 4548
rect 8996 4536 9002 4548
rect 10413 4539 10471 4545
rect 10413 4536 10425 4539
rect 8996 4508 10425 4536
rect 8996 4496 9002 4508
rect 10413 4505 10425 4508
rect 10459 4505 10471 4539
rect 13004 4536 13032 4567
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 15378 4604 15384 4616
rect 15339 4576 15384 4604
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 17310 4604 17316 4616
rect 17271 4576 17316 4604
rect 17310 4564 17316 4576
rect 17368 4564 17374 4616
rect 17420 4613 17448 4644
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 14274 4536 14280 4548
rect 13004 4508 14280 4536
rect 10413 4499 10471 4505
rect 14274 4496 14280 4508
rect 14332 4496 14338 4548
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 3329 4471 3387 4477
rect 3329 4468 3341 4471
rect 3292 4440 3341 4468
rect 3292 4428 3298 4440
rect 3329 4437 3341 4440
rect 3375 4437 3387 4471
rect 4430 4468 4436 4480
rect 4391 4440 4436 4468
rect 3329 4431 3387 4437
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 7101 4471 7159 4477
rect 7101 4437 7113 4471
rect 7147 4468 7159 4471
rect 9582 4468 9588 4480
rect 7147 4440 9588 4468
rect 7147 4437 7159 4440
rect 7101 4431 7159 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 9861 4471 9919 4477
rect 9861 4437 9873 4471
rect 9907 4468 9919 4471
rect 11790 4468 11796 4480
rect 9907 4440 11796 4468
rect 9907 4437 9919 4440
rect 9861 4431 9919 4437
rect 11790 4428 11796 4440
rect 11848 4428 11854 4480
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 1854 4264 1860 4276
rect 1815 4236 1860 4264
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 3326 4224 3332 4276
rect 3384 4264 3390 4276
rect 3384 4236 4936 4264
rect 3384 4224 3390 4236
rect 4706 4196 4712 4208
rect 4632 4168 4712 4196
rect 4430 4128 4436 4140
rect 4391 4100 4436 4128
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 4632 4137 4660 4168
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 4908 4196 4936 4236
rect 4982 4224 4988 4276
rect 5040 4264 5046 4276
rect 5994 4264 6000 4276
rect 5040 4236 6000 4264
rect 5040 4224 5046 4236
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 11054 4264 11060 4276
rect 6840 4236 11060 4264
rect 4908 4168 5396 4196
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 5368 4128 5396 4168
rect 5442 4156 5448 4208
rect 5500 4196 5506 4208
rect 6840 4196 6868 4236
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 5500 4168 5764 4196
rect 5500 4156 5506 4168
rect 5736 4137 5764 4168
rect 5828 4168 6868 4196
rect 5721 4131 5779 4137
rect 5368 4100 5672 4128
rect 4617 4091 4675 4097
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4029 1731 4063
rect 2397 4063 2455 4069
rect 2397 4060 2409 4063
rect 1673 4023 1731 4029
rect 2332 4032 2409 4060
rect 1688 3992 1716 4023
rect 2130 3992 2136 4004
rect 1688 3964 2136 3992
rect 2130 3952 2136 3964
rect 2188 3952 2194 4004
rect 2332 3992 2360 4032
rect 2397 4029 2409 4032
rect 2443 4029 2455 4063
rect 2397 4023 2455 4029
rect 3145 4063 3203 4069
rect 3145 4029 3157 4063
rect 3191 4060 3203 4063
rect 4706 4060 4712 4072
rect 3191 4032 4712 4060
rect 3191 4029 3203 4032
rect 3145 4023 3203 4029
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 4798 4020 4804 4072
rect 4856 4060 4862 4072
rect 5350 4060 5356 4072
rect 4856 4032 5356 4060
rect 4856 4020 4862 4032
rect 5350 4020 5356 4032
rect 5408 4060 5414 4072
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 5408 4032 5549 4060
rect 5408 4020 5414 4032
rect 5537 4029 5549 4032
rect 5583 4029 5595 4063
rect 5644 4060 5672 4100
rect 5721 4097 5733 4131
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 5828 4060 5856 4168
rect 8386 4156 8392 4208
rect 8444 4196 8450 4208
rect 8938 4196 8944 4208
rect 8444 4168 8944 4196
rect 8444 4156 8450 4168
rect 8938 4156 8944 4168
rect 8996 4196 9002 4208
rect 9125 4199 9183 4205
rect 9125 4196 9137 4199
rect 8996 4168 9137 4196
rect 8996 4156 9002 4168
rect 9125 4165 9137 4168
rect 9171 4165 9183 4199
rect 9125 4159 9183 4165
rect 9677 4199 9735 4205
rect 9677 4165 9689 4199
rect 9723 4196 9735 4199
rect 10318 4196 10324 4208
rect 9723 4168 10324 4196
rect 9723 4165 9735 4168
rect 9677 4159 9735 4165
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6328 4100 6837 4128
rect 6328 4088 6334 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 9140 4128 9168 4159
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 12897 4131 12955 4137
rect 9140 4100 9812 4128
rect 6825 4091 6883 4097
rect 7834 4060 7840 4072
rect 5644 4032 5856 4060
rect 7024 4032 7840 4060
rect 5537 4023 5595 4029
rect 3050 3992 3056 4004
rect 2332 3964 3056 3992
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 3878 3952 3884 4004
rect 3936 3992 3942 4004
rect 7024 3992 7052 4032
rect 7834 4020 7840 4032
rect 7892 4020 7898 4072
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4029 9551 4063
rect 9784 4060 9812 4100
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13170 4128 13176 4140
rect 12943 4100 13176 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 13354 4128 13360 4140
rect 13315 4100 13360 4128
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 14918 4128 14924 4140
rect 14879 4100 14924 4128
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15988 4100 16129 4128
rect 15988 4088 15994 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 16942 4128 16948 4140
rect 16903 4100 16948 4128
rect 16117 4091 16175 4097
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 10042 4060 10048 4072
rect 9784 4032 10048 4060
rect 9493 4023 9551 4029
rect 3936 3964 7052 3992
rect 7092 3995 7150 4001
rect 3936 3952 3942 3964
rect 7092 3961 7104 3995
rect 7138 3992 7150 3995
rect 7282 3992 7288 4004
rect 7138 3964 7288 3992
rect 7138 3961 7150 3964
rect 7092 3955 7150 3961
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 9508 3992 9536 4023
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 10321 4063 10379 4069
rect 10321 4029 10333 4063
rect 10367 4060 10379 4063
rect 10962 4060 10968 4072
rect 10367 4032 10968 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 10410 3992 10416 4004
rect 9508 3964 10416 3992
rect 10410 3952 10416 3964
rect 10468 3952 10474 4004
rect 10588 3995 10646 4001
rect 10588 3961 10600 3995
rect 10634 3992 10646 3995
rect 10778 3992 10784 4004
rect 10634 3964 10784 3992
rect 10634 3961 10646 3964
rect 10588 3955 10646 3961
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 12526 3952 12532 4004
rect 12584 3992 12590 4004
rect 12989 3995 13047 4001
rect 12989 3992 13001 3995
rect 12584 3964 13001 3992
rect 12584 3952 12590 3964
rect 12989 3961 13001 3964
rect 13035 3961 13047 3995
rect 12989 3955 13047 3961
rect 14090 3952 14096 4004
rect 14148 3992 14154 4004
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 14148 3964 14473 3992
rect 14148 3952 14154 3964
rect 14461 3961 14473 3964
rect 14507 3961 14519 3995
rect 14461 3955 14519 3961
rect 14550 3952 14556 4004
rect 14608 3992 14614 4004
rect 14608 3964 14653 3992
rect 14608 3952 14614 3964
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 16209 3995 16267 4001
rect 16209 3992 16221 3995
rect 15988 3964 16221 3992
rect 15988 3952 15994 3964
rect 16209 3961 16221 3964
rect 16255 3961 16267 3995
rect 16209 3955 16267 3961
rect 2593 3927 2651 3933
rect 2593 3893 2605 3927
rect 2639 3924 2651 3927
rect 2774 3924 2780 3936
rect 2639 3896 2780 3924
rect 2639 3893 2651 3896
rect 2593 3887 2651 3893
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 3326 3924 3332 3936
rect 3287 3896 3332 3924
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 3973 3927 4031 3933
rect 3973 3924 3985 3927
rect 3844 3896 3985 3924
rect 3844 3884 3850 3896
rect 3973 3893 3985 3896
rect 4019 3893 4031 3927
rect 3973 3887 4031 3893
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3924 4399 3927
rect 5169 3927 5227 3933
rect 5169 3924 5181 3927
rect 4387 3896 5181 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 5169 3893 5181 3896
rect 5215 3893 5227 3927
rect 5169 3887 5227 3893
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5629 3927 5687 3933
rect 5629 3924 5641 3927
rect 5316 3896 5641 3924
rect 5316 3884 5322 3896
rect 5629 3893 5641 3896
rect 5675 3924 5687 3927
rect 6454 3924 6460 3936
rect 5675 3896 6460 3924
rect 5675 3893 5687 3896
rect 5629 3887 5687 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 8205 3927 8263 3933
rect 8205 3893 8217 3927
rect 8251 3924 8263 3927
rect 8478 3924 8484 3936
rect 8251 3896 8484 3924
rect 8251 3893 8263 3896
rect 8205 3887 8263 3893
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11020 3896 11713 3924
rect 11020 3884 11026 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 15746 3924 15752 3936
rect 15252 3896 15752 3924
rect 15252 3884 15258 3896
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 4890 3720 4896 3732
rect 2179 3692 4896 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 2148 3584 2176 3683
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 5442 3720 5448 3732
rect 5403 3692 5448 3720
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 6270 3720 6276 3732
rect 5920 3692 6276 3720
rect 4246 3652 4252 3664
rect 4080 3624 4252 3652
rect 1719 3556 2176 3584
rect 2869 3587 2927 3593
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 2869 3553 2881 3587
rect 2915 3584 2927 3587
rect 3878 3584 3884 3596
rect 2915 3556 3884 3584
rect 2915 3553 2927 3556
rect 2869 3547 2927 3553
rect 3878 3544 3884 3556
rect 3936 3544 3942 3596
rect 4080 3593 4108 3624
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 4430 3612 4436 3664
rect 4488 3652 4494 3664
rect 5074 3652 5080 3664
rect 4488 3624 5080 3652
rect 4488 3612 4494 3624
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 4332 3587 4390 3593
rect 4332 3553 4344 3587
rect 4378 3584 4390 3587
rect 4614 3584 4620 3596
rect 4378 3556 4620 3584
rect 4378 3553 4390 3556
rect 4332 3547 4390 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 5920 3593 5948 3692
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 7282 3720 7288 3732
rect 7243 3692 7288 3720
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 8662 3720 8668 3732
rect 7791 3692 8668 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 8864 3692 14412 3720
rect 6172 3655 6230 3661
rect 6172 3621 6184 3655
rect 6218 3652 6230 3655
rect 7374 3652 7380 3664
rect 6218 3624 7380 3652
rect 6218 3621 6230 3624
rect 6172 3615 6230 3621
rect 7374 3612 7380 3624
rect 7432 3652 7438 3664
rect 7650 3652 7656 3664
rect 7432 3624 7656 3652
rect 7432 3612 7438 3624
rect 7650 3612 7656 3624
rect 7708 3612 7714 3664
rect 8864 3652 8892 3692
rect 7760 3624 8892 3652
rect 5905 3587 5963 3593
rect 5905 3553 5917 3587
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 7760 3584 7788 3624
rect 8938 3612 8944 3664
rect 8996 3652 9002 3664
rect 9125 3655 9183 3661
rect 9125 3652 9137 3655
rect 8996 3624 9137 3652
rect 8996 3612 9002 3624
rect 9125 3621 9137 3624
rect 9171 3652 9183 3655
rect 9214 3652 9220 3664
rect 9171 3624 9220 3652
rect 9171 3621 9183 3624
rect 9125 3615 9183 3621
rect 9214 3612 9220 3624
rect 9272 3612 9278 3664
rect 10594 3612 10600 3664
rect 10652 3652 10658 3664
rect 10778 3652 10784 3664
rect 10652 3624 10784 3652
rect 10652 3612 10658 3624
rect 10778 3612 10784 3624
rect 10836 3612 10842 3664
rect 11422 3652 11428 3664
rect 11383 3624 11428 3652
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 12342 3652 12348 3664
rect 12303 3624 12348 3652
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 12897 3655 12955 3661
rect 12897 3652 12909 3655
rect 12636 3624 12909 3652
rect 8386 3584 8392 3596
rect 6512 3556 7788 3584
rect 8347 3556 8392 3584
rect 6512 3544 6518 3556
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3584 8815 3587
rect 9030 3584 9036 3596
rect 8803 3556 9036 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 10318 3584 10324 3596
rect 9640 3556 10324 3584
rect 9640 3544 9646 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 10410 3544 10416 3596
rect 10468 3584 10474 3596
rect 10962 3584 10968 3596
rect 10468 3556 10968 3584
rect 10468 3544 10474 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 12308 3556 12388 3584
rect 12308 3544 12314 3556
rect 3050 3516 3056 3528
rect 3011 3488 3056 3516
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 7190 3476 7196 3528
rect 7248 3516 7254 3528
rect 10781 3519 10839 3525
rect 10781 3516 10793 3519
rect 7248 3488 10793 3516
rect 7248 3476 7254 3488
rect 10781 3485 10793 3488
rect 10827 3516 10839 3519
rect 11054 3516 11060 3528
rect 10827 3488 11060 3516
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 11606 3516 11612 3528
rect 11379 3488 11612 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 12360 3516 12388 3556
rect 12636 3516 12664 3624
rect 12897 3621 12909 3624
rect 12943 3621 12955 3655
rect 12897 3615 12955 3621
rect 12989 3655 13047 3661
rect 12989 3621 13001 3655
rect 13035 3652 13047 3655
rect 13538 3652 13544 3664
rect 13035 3624 13544 3652
rect 13035 3621 13047 3624
rect 12989 3615 13047 3621
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 14384 3652 14412 3692
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 15378 3720 15384 3732
rect 14700 3692 15384 3720
rect 14700 3680 14706 3692
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 15473 3723 15531 3729
rect 15473 3689 15485 3723
rect 15519 3689 15531 3723
rect 15838 3720 15844 3732
rect 15799 3692 15844 3720
rect 15473 3683 15531 3689
rect 15488 3652 15516 3683
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16632 3692 16681 3720
rect 16632 3680 16638 3692
rect 16669 3689 16681 3692
rect 16715 3689 16727 3723
rect 16669 3683 16727 3689
rect 16758 3680 16764 3732
rect 16816 3720 16822 3732
rect 16816 3692 17448 3720
rect 16816 3680 16822 3692
rect 17310 3652 17316 3664
rect 14384 3624 15424 3652
rect 15488 3624 17316 3652
rect 15396 3596 15424 3624
rect 17310 3612 17316 3624
rect 17368 3612 17374 3664
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 14461 3587 14519 3593
rect 14461 3584 14473 3587
rect 13872 3556 14473 3584
rect 13872 3544 13878 3556
rect 14461 3553 14473 3556
rect 14507 3553 14519 3587
rect 14461 3547 14519 3553
rect 15378 3544 15384 3596
rect 15436 3544 15442 3596
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 15933 3587 15991 3593
rect 15933 3584 15945 3587
rect 15528 3556 15945 3584
rect 15528 3544 15534 3556
rect 15933 3553 15945 3556
rect 15979 3553 15991 3587
rect 17034 3584 17040 3596
rect 16995 3556 17040 3584
rect 15933 3547 15991 3553
rect 17034 3544 17040 3556
rect 17092 3544 17098 3596
rect 17129 3587 17187 3593
rect 17129 3553 17141 3587
rect 17175 3584 17187 3587
rect 17420 3584 17448 3692
rect 17862 3680 17868 3732
rect 17920 3720 17926 3732
rect 18049 3723 18107 3729
rect 18049 3720 18061 3723
rect 17920 3692 18061 3720
rect 17920 3680 17926 3692
rect 18049 3689 18061 3692
rect 18095 3689 18107 3723
rect 18049 3683 18107 3689
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17175 3556 17356 3584
rect 17420 3556 17877 3584
rect 17175 3553 17187 3556
rect 17129 3547 17187 3553
rect 13722 3516 13728 3528
rect 12360 3488 12664 3516
rect 13683 3488 13728 3516
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 15746 3476 15752 3528
rect 15804 3516 15810 3528
rect 16117 3519 16175 3525
rect 16117 3516 16129 3519
rect 15804 3488 16129 3516
rect 15804 3476 15810 3488
rect 16117 3485 16129 3488
rect 16163 3516 16175 3519
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 16163 3488 17233 3516
rect 16163 3485 16175 3488
rect 16117 3479 16175 3485
rect 17221 3485 17233 3488
rect 17267 3485 17279 3519
rect 17221 3479 17279 3485
rect 1854 3448 1860 3460
rect 1815 3420 1860 3448
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 7742 3408 7748 3460
rect 7800 3448 7806 3460
rect 9950 3448 9956 3460
rect 7800 3420 9956 3448
rect 7800 3408 7806 3420
rect 9950 3408 9956 3420
rect 10008 3408 10014 3460
rect 10042 3408 10048 3460
rect 10100 3448 10106 3460
rect 10100 3420 10145 3448
rect 10100 3408 10106 3420
rect 12618 3408 12624 3460
rect 12676 3448 12682 3460
rect 14366 3448 14372 3460
rect 12676 3420 14372 3448
rect 12676 3408 12682 3420
rect 14366 3408 14372 3420
rect 14424 3408 14430 3460
rect 17328 3448 17356 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 14568 3420 17356 3448
rect 5166 3340 5172 3392
rect 5224 3380 5230 3392
rect 10410 3380 10416 3392
rect 5224 3352 10416 3380
rect 5224 3340 5230 3352
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 14568 3380 14596 3420
rect 11756 3352 14596 3380
rect 14645 3383 14703 3389
rect 11756 3340 11762 3352
rect 14645 3349 14657 3383
rect 14691 3380 14703 3383
rect 15194 3380 15200 3392
rect 14691 3352 15200 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 15194 3340 15200 3352
rect 15252 3340 15258 3392
rect 15378 3340 15384 3392
rect 15436 3380 15442 3392
rect 16390 3380 16396 3392
rect 15436 3352 16396 3380
rect 15436 3340 15442 3352
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 5445 3179 5503 3185
rect 5445 3145 5457 3179
rect 5491 3176 5503 3179
rect 7650 3176 7656 3188
rect 5491 3148 7656 3176
rect 5491 3145 5503 3148
rect 5445 3139 5503 3145
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 12250 3176 12256 3188
rect 8312 3148 12256 3176
rect 6181 3111 6239 3117
rect 2424 3080 5212 3108
rect 198 3000 204 3052
rect 256 3040 262 3052
rect 1762 3040 1768 3052
rect 256 3012 1768 3040
rect 256 3000 262 3012
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 1489 2975 1547 2981
rect 1489 2941 1501 2975
rect 1535 2972 1547 2975
rect 1578 2972 1584 2984
rect 1535 2944 1584 2972
rect 1535 2941 1547 2944
rect 1489 2935 1547 2941
rect 1578 2932 1584 2944
rect 1636 2932 1642 2984
rect 2424 2981 2452 3080
rect 4522 3040 4528 3052
rect 4264 3012 4528 3040
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2941 2467 2975
rect 2409 2935 2467 2941
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2972 3387 2975
rect 3786 2972 3792 2984
rect 3375 2944 3792 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 4264 2981 4292 3012
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 4249 2975 4307 2981
rect 4249 2941 4261 2975
rect 4295 2941 4307 2975
rect 4249 2935 4307 2941
rect 658 2864 664 2916
rect 716 2904 722 2916
rect 1765 2907 1823 2913
rect 1765 2904 1777 2907
rect 716 2876 1777 2904
rect 716 2864 722 2876
rect 1765 2873 1777 2876
rect 1811 2873 1823 2907
rect 1765 2867 1823 2873
rect 2130 2864 2136 2916
rect 2188 2904 2194 2916
rect 2685 2907 2743 2913
rect 2685 2904 2697 2907
rect 2188 2876 2697 2904
rect 2188 2864 2194 2876
rect 2685 2873 2697 2876
rect 2731 2873 2743 2907
rect 2685 2867 2743 2873
rect 3142 2864 3148 2916
rect 3200 2904 3206 2916
rect 3605 2907 3663 2913
rect 3605 2904 3617 2907
rect 3200 2876 3617 2904
rect 3200 2864 3206 2876
rect 3605 2873 3617 2876
rect 3651 2873 3663 2907
rect 3605 2867 3663 2873
rect 4525 2907 4583 2913
rect 4525 2873 4537 2907
rect 4571 2873 4583 2907
rect 5184 2904 5212 3080
rect 6181 3077 6193 3111
rect 6227 3108 6239 3111
rect 6454 3108 6460 3120
rect 6227 3080 6460 3108
rect 6227 3077 6239 3080
rect 6181 3071 6239 3077
rect 6454 3068 6460 3080
rect 6512 3068 6518 3120
rect 7377 3111 7435 3117
rect 7377 3077 7389 3111
rect 7423 3108 7435 3111
rect 8312 3108 8340 3148
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 17034 3176 17040 3188
rect 12400 3148 17040 3176
rect 12400 3136 12406 3148
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 11146 3108 11152 3120
rect 7423 3080 8340 3108
rect 8864 3080 11152 3108
rect 7423 3077 7435 3080
rect 7377 3071 7435 3077
rect 7392 3040 7420 3071
rect 5276 3012 7420 3040
rect 5276 2981 5304 3012
rect 7558 3000 7564 3052
rect 7616 3000 7622 3052
rect 8864 3049 8892 3080
rect 11146 3068 11152 3080
rect 11204 3068 11210 3120
rect 11422 3068 11428 3120
rect 11480 3108 11486 3120
rect 17451 3111 17509 3117
rect 17451 3108 17463 3111
rect 11480 3080 17463 3108
rect 11480 3068 11486 3080
rect 17451 3077 17463 3080
rect 17497 3077 17509 3111
rect 17451 3071 17509 3077
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3009 8907 3043
rect 9766 3040 9772 3052
rect 9727 3012 9772 3040
rect 8849 3003 8907 3009
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 10413 3043 10471 3049
rect 10413 3009 10425 3043
rect 10459 3040 10471 3043
rect 10870 3040 10876 3052
rect 10459 3012 10876 3040
rect 10459 3009 10471 3012
rect 10413 3003 10471 3009
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11238 3040 11244 3052
rect 11199 3012 11244 3040
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 12986 3040 12992 3052
rect 12947 3012 12992 3040
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 14550 3040 14556 3052
rect 13136 3012 14556 3040
rect 13136 3000 13142 3012
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 14734 3000 14740 3052
rect 14792 3040 14798 3052
rect 15289 3043 15347 3049
rect 14792 3012 15240 3040
rect 14792 3000 14798 3012
rect 5261 2975 5319 2981
rect 5261 2941 5273 2975
rect 5307 2941 5319 2975
rect 5261 2935 5319 2941
rect 5350 2932 5356 2984
rect 5408 2972 5414 2984
rect 5997 2975 6055 2981
rect 5997 2972 6009 2975
rect 5408 2944 6009 2972
rect 5408 2932 5414 2944
rect 5997 2941 6009 2944
rect 6043 2941 6055 2975
rect 5997 2935 6055 2941
rect 6730 2932 6736 2984
rect 6788 2972 6794 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6788 2944 6837 2972
rect 6788 2932 6794 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 7282 2972 7288 2984
rect 7239 2944 7288 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7576 2972 7604 3000
rect 7392 2944 7604 2972
rect 8021 2975 8079 2981
rect 7392 2904 7420 2944
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8662 2972 8668 2984
rect 8067 2944 8668 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 15212 2972 15240 3012
rect 15289 3009 15301 3043
rect 15335 3040 15347 3043
rect 15562 3040 15568 3052
rect 15335 3012 15568 3040
rect 15335 3009 15347 3012
rect 15289 3003 15347 3009
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 15841 3043 15899 3049
rect 15841 3040 15853 3043
rect 15672 3012 15853 3040
rect 15672 2972 15700 3012
rect 15841 3009 15853 3012
rect 15887 3009 15899 3043
rect 16850 3040 16856 3052
rect 16811 3012 16856 3040
rect 15841 3003 15899 3009
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 17348 2975 17406 2981
rect 17348 2972 17360 2975
rect 15212 2944 15700 2972
rect 16684 2944 17360 2972
rect 5184 2876 7420 2904
rect 4525 2867 4583 2873
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 4540 2836 4568 2867
rect 7558 2864 7564 2916
rect 7616 2904 7622 2916
rect 8941 2907 8999 2913
rect 7616 2876 8800 2904
rect 7616 2864 7622 2876
rect 1728 2808 4568 2836
rect 1728 2796 1734 2808
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 7742 2836 7748 2848
rect 4764 2808 7748 2836
rect 4764 2796 4770 2808
rect 7742 2796 7748 2808
rect 7800 2796 7806 2848
rect 8205 2839 8263 2845
rect 8205 2805 8217 2839
rect 8251 2836 8263 2839
rect 8662 2836 8668 2848
rect 8251 2808 8668 2836
rect 8251 2805 8263 2808
rect 8205 2799 8263 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 8772 2836 8800 2876
rect 8941 2873 8953 2907
rect 8987 2904 8999 2907
rect 9766 2904 9772 2916
rect 8987 2876 9772 2904
rect 8987 2873 8999 2876
rect 8941 2867 8999 2873
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 10502 2904 10508 2916
rect 10463 2876 10508 2904
rect 10502 2864 10508 2876
rect 10560 2864 10566 2916
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 12713 2907 12771 2913
rect 12713 2904 12725 2907
rect 10836 2876 12725 2904
rect 10836 2864 10842 2876
rect 12713 2873 12725 2876
rect 12759 2873 12771 2907
rect 12713 2867 12771 2873
rect 12805 2907 12863 2913
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 13078 2904 13084 2916
rect 12851 2876 13084 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 13078 2864 13084 2876
rect 13136 2864 13142 2916
rect 14277 2907 14335 2913
rect 14277 2904 14289 2907
rect 14108 2876 14289 2904
rect 10594 2836 10600 2848
rect 8772 2808 10600 2836
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 10686 2796 10692 2848
rect 10744 2836 10750 2848
rect 14108 2836 14136 2876
rect 14277 2873 14289 2876
rect 14323 2873 14335 2907
rect 14277 2867 14335 2873
rect 14366 2864 14372 2916
rect 14424 2904 14430 2916
rect 14424 2876 14469 2904
rect 14424 2864 14430 2876
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 15654 2904 15660 2916
rect 14884 2876 15660 2904
rect 14884 2864 14890 2876
rect 15654 2864 15660 2876
rect 15712 2864 15718 2916
rect 15930 2904 15936 2916
rect 15891 2876 15936 2904
rect 15930 2864 15936 2876
rect 15988 2864 15994 2916
rect 10744 2808 14136 2836
rect 10744 2796 10750 2808
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 16684 2836 16712 2944
rect 17348 2941 17360 2944
rect 17394 2941 17406 2975
rect 17348 2935 17406 2941
rect 14608 2808 16712 2836
rect 14608 2796 14614 2808
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 2685 2635 2743 2641
rect 2685 2601 2697 2635
rect 2731 2632 2743 2635
rect 2774 2632 2780 2644
rect 2731 2604 2780 2632
rect 2731 2601 2743 2604
rect 2685 2595 2743 2601
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 5537 2635 5595 2641
rect 5537 2601 5549 2635
rect 5583 2632 5595 2635
rect 8110 2632 8116 2644
rect 5583 2604 8116 2632
rect 5583 2601 5595 2604
rect 5537 2595 5595 2601
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 11977 2635 12035 2641
rect 11977 2601 11989 2635
rect 12023 2632 12035 2635
rect 15194 2632 15200 2644
rect 12023 2604 15200 2632
rect 12023 2601 12035 2604
rect 11977 2595 12035 2601
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 17678 2632 17684 2644
rect 17639 2604 17684 2632
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 3510 2564 3516 2576
rect 1596 2536 3516 2564
rect 1596 2505 1624 2536
rect 3510 2524 3516 2536
rect 3568 2524 3574 2576
rect 10226 2564 10232 2576
rect 6012 2536 8892 2564
rect 10187 2536 10232 2564
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2465 1639 2499
rect 1581 2459 1639 2465
rect 2501 2499 2559 2505
rect 2501 2465 2513 2499
rect 2547 2465 2559 2499
rect 2501 2459 2559 2465
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2465 3295 2499
rect 3237 2459 3295 2465
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4798 2496 4804 2508
rect 4111 2468 4804 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 1118 2388 1124 2440
rect 1176 2428 1182 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 1176 2400 1777 2428
rect 1176 2388 1182 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2516 2360 2544 2459
rect 3252 2428 3280 2459
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 5353 2499 5411 2505
rect 5353 2465 5365 2499
rect 5399 2496 5411 2499
rect 6012 2496 6040 2536
rect 5399 2468 6040 2496
rect 6089 2499 6147 2505
rect 5399 2465 5411 2468
rect 5353 2459 5411 2465
rect 6089 2465 6101 2499
rect 6135 2496 6147 2499
rect 7190 2496 7196 2508
rect 6135 2468 7196 2496
rect 6135 2465 6147 2468
rect 6089 2459 6147 2465
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 7374 2496 7380 2508
rect 7331 2468 7380 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 4982 2428 4988 2440
rect 3252 2400 4988 2428
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 7558 2428 7564 2440
rect 6288 2400 7564 2428
rect 4430 2360 4436 2372
rect 2516 2332 4436 2360
rect 4430 2320 4436 2332
rect 4488 2320 4494 2372
rect 6288 2369 6316 2400
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 7926 2428 7932 2440
rect 7699 2400 7932 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2428 8171 2431
rect 8386 2428 8392 2440
rect 8159 2400 8392 2428
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 6273 2363 6331 2369
rect 6273 2329 6285 2363
rect 6319 2329 6331 2363
rect 6273 2323 6331 2329
rect 6730 2320 6736 2372
rect 6788 2360 6794 2372
rect 6917 2363 6975 2369
rect 6917 2360 6929 2363
rect 6788 2332 6929 2360
rect 6788 2320 6794 2332
rect 6917 2329 6929 2332
rect 6963 2360 6975 2363
rect 8128 2360 8156 2391
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 8864 2437 8892 2536
rect 10226 2524 10232 2536
rect 10284 2524 10290 2576
rect 10321 2567 10379 2573
rect 10321 2533 10333 2567
rect 10367 2564 10379 2567
rect 10410 2564 10416 2576
rect 10367 2536 10416 2564
rect 10367 2533 10379 2536
rect 10321 2527 10379 2533
rect 10410 2524 10416 2536
rect 10468 2524 10474 2576
rect 11241 2567 11299 2573
rect 11241 2533 11253 2567
rect 11287 2564 11299 2567
rect 11330 2564 11336 2576
rect 11287 2536 11336 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 11330 2524 11336 2536
rect 11388 2524 11394 2576
rect 13357 2567 13415 2573
rect 13357 2533 13369 2567
rect 13403 2564 13415 2567
rect 13446 2564 13452 2576
rect 13403 2536 13452 2564
rect 13403 2533 13415 2536
rect 13357 2527 13415 2533
rect 13446 2524 13452 2536
rect 13504 2524 13510 2576
rect 14274 2564 14280 2576
rect 14235 2536 14280 2564
rect 14274 2524 14280 2536
rect 14332 2524 14338 2576
rect 15010 2524 15016 2576
rect 15068 2564 15074 2576
rect 15657 2567 15715 2573
rect 15657 2564 15669 2567
rect 15068 2536 15669 2564
rect 15068 2524 15074 2536
rect 15657 2533 15669 2536
rect 15703 2533 15715 2567
rect 15657 2527 15715 2533
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11756 2468 11805 2496
rect 11756 2456 11762 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 14804 2499 14862 2505
rect 14804 2465 14816 2499
rect 14850 2496 14862 2499
rect 17497 2499 17555 2505
rect 14850 2468 15056 2496
rect 14850 2465 14862 2468
rect 14804 2459 14862 2465
rect 8849 2431 8907 2437
rect 8849 2397 8861 2431
rect 8895 2428 8907 2431
rect 12526 2428 12532 2440
rect 8895 2400 12532 2428
rect 8895 2397 8907 2400
rect 8849 2391 8907 2397
rect 12526 2388 12532 2400
rect 12584 2388 12590 2440
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 12676 2400 13277 2428
rect 12676 2388 12682 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 6963 2332 8156 2360
rect 6963 2329 6975 2332
rect 6917 2323 6975 2329
rect 9766 2320 9772 2372
rect 9824 2360 9830 2372
rect 14875 2363 14933 2369
rect 14875 2360 14887 2363
rect 9824 2332 14887 2360
rect 9824 2320 9830 2332
rect 14875 2329 14887 2332
rect 14921 2329 14933 2363
rect 14875 2323 14933 2329
rect 3418 2292 3424 2304
rect 3379 2264 3424 2292
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 4249 2295 4307 2301
rect 4249 2292 4261 2295
rect 3568 2264 4261 2292
rect 3568 2252 3574 2264
rect 4249 2261 4261 2264
rect 4295 2261 4307 2295
rect 4249 2255 4307 2261
rect 10502 2252 10508 2304
rect 10560 2292 10566 2304
rect 15028 2292 15056 2468
rect 17497 2465 17509 2499
rect 17543 2496 17555 2499
rect 17770 2496 17776 2508
rect 17543 2468 17776 2496
rect 17543 2465 17555 2468
rect 17497 2459 17555 2465
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 15102 2388 15108 2440
rect 15160 2428 15166 2440
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 15160 2400 15577 2428
rect 15160 2388 15166 2400
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 16482 2428 16488 2440
rect 16443 2400 16488 2428
rect 15565 2391 15623 2397
rect 16482 2388 16488 2400
rect 16540 2388 16546 2440
rect 10560 2264 15056 2292
rect 10560 2252 10566 2264
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 7926 1980 7932 2032
rect 7984 2020 7990 2032
rect 10410 2020 10416 2032
rect 7984 1992 10416 2020
rect 7984 1980 7990 1992
rect 10410 1980 10416 1992
rect 10468 2020 10474 2032
rect 14550 2020 14556 2032
rect 10468 1992 14556 2020
rect 10468 1980 10474 1992
rect 14550 1980 14556 1992
rect 14608 1980 14614 2032
rect 13906 1368 13912 1420
rect 13964 1408 13970 1420
rect 16666 1408 16672 1420
rect 13964 1380 16672 1408
rect 13964 1368 13970 1380
rect 16666 1368 16672 1380
rect 16724 1368 16730 1420
<< via1 >>
rect 3700 15240 3752 15292
rect 6000 15240 6052 15292
rect 4068 15172 4120 15224
rect 8116 15172 8168 15224
rect 12164 15172 12216 15224
rect 15936 15172 15988 15224
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 940 14560 992 14612
rect 2228 14560 2280 14612
rect 2780 14492 2832 14544
rect 13636 14492 13688 14544
rect 15016 14424 15068 14476
rect 15752 14424 15804 14476
rect 16304 14424 16356 14476
rect 12256 14356 12308 14408
rect 17684 14356 17736 14408
rect 4068 14288 4120 14340
rect 12716 14288 12768 14340
rect 13728 14288 13780 14340
rect 15384 14288 15436 14340
rect 3056 14220 3108 14272
rect 13452 14220 13504 14272
rect 14004 14220 14056 14272
rect 15200 14220 15252 14272
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 1584 14016 1636 14068
rect 2872 14016 2924 14068
rect 3700 14016 3752 14068
rect 5724 14016 5776 14068
rect 6736 14016 6788 14068
rect 13544 14016 13596 14068
rect 15568 14016 15620 14068
rect 5908 13948 5960 14000
rect 9404 13880 9456 13932
rect 16212 13880 16264 13932
rect 2780 13812 2832 13864
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 5816 13812 5868 13864
rect 6092 13812 6144 13864
rect 14188 13812 14240 13864
rect 14372 13812 14424 13864
rect 14924 13812 14976 13864
rect 15108 13812 15160 13864
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 7380 13744 7432 13796
rect 9220 13744 9272 13796
rect 9312 13744 9364 13796
rect 10232 13744 10284 13796
rect 11244 13744 11296 13796
rect 11980 13744 12032 13796
rect 3516 13676 3568 13728
rect 14004 13676 14056 13728
rect 19616 13676 19668 13728
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 296 13472 348 13524
rect 4252 13472 4304 13524
rect 13544 13472 13596 13524
rect 13636 13472 13688 13524
rect 18328 13472 18380 13524
rect 1860 13404 1912 13456
rect 5448 13404 5500 13456
rect 15568 13404 15620 13456
rect 4804 13336 4856 13388
rect 15200 13336 15252 13388
rect 16488 13336 16540 13388
rect 17868 13379 17920 13388
rect 17868 13345 17877 13379
rect 17877 13345 17911 13379
rect 17911 13345 17920 13379
rect 17868 13336 17920 13345
rect 2964 13311 3016 13320
rect 1952 13132 2004 13184
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 9772 13268 9824 13320
rect 17040 13268 17092 13320
rect 7472 13200 7524 13252
rect 15016 13200 15068 13252
rect 18972 13200 19024 13252
rect 3700 13132 3752 13184
rect 4712 13132 4764 13184
rect 12716 13132 12768 13184
rect 13176 13132 13228 13184
rect 15384 13132 15436 13184
rect 15476 13132 15528 13184
rect 18052 13175 18104 13184
rect 18052 13141 18061 13175
rect 18061 13141 18095 13175
rect 18095 13141 18104 13175
rect 18052 13132 18104 13141
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 4436 12928 4488 12980
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 1952 12767 2004 12776
rect 1952 12733 1961 12767
rect 1961 12733 1995 12767
rect 1995 12733 2004 12767
rect 1952 12724 2004 12733
rect 2964 12656 3016 12708
rect 4988 12724 5040 12776
rect 15200 12860 15252 12912
rect 15384 12860 15436 12912
rect 6644 12792 6696 12844
rect 11428 12792 11480 12844
rect 17960 12860 18012 12912
rect 7840 12724 7892 12776
rect 8024 12724 8076 12776
rect 8668 12724 8720 12776
rect 10876 12724 10928 12776
rect 12624 12724 12676 12776
rect 14004 12724 14056 12776
rect 14372 12724 14424 12776
rect 8576 12699 8628 12708
rect 8576 12665 8585 12699
rect 8585 12665 8619 12699
rect 8619 12665 8628 12699
rect 8576 12656 8628 12665
rect 8760 12656 8812 12708
rect 13912 12656 13964 12708
rect 14740 12656 14792 12708
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 2780 12588 2832 12640
rect 3792 12588 3844 12640
rect 4620 12631 4672 12640
rect 4620 12597 4629 12631
rect 4629 12597 4663 12631
rect 4663 12597 4672 12631
rect 4620 12588 4672 12597
rect 5540 12631 5592 12640
rect 5540 12597 5549 12631
rect 5549 12597 5583 12631
rect 5583 12597 5592 12631
rect 5540 12588 5592 12597
rect 6000 12631 6052 12640
rect 6000 12597 6009 12631
rect 6009 12597 6043 12631
rect 6043 12597 6052 12631
rect 6000 12588 6052 12597
rect 7288 12588 7340 12640
rect 13268 12588 13320 12640
rect 14556 12588 14608 12640
rect 15016 12588 15068 12640
rect 16396 12588 16448 12640
rect 17408 12631 17460 12640
rect 17408 12597 17417 12631
rect 17417 12597 17451 12631
rect 17451 12597 17460 12631
rect 17408 12588 17460 12597
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 2044 12384 2096 12436
rect 2596 12384 2648 12436
rect 5632 12384 5684 12436
rect 9588 12384 9640 12436
rect 11060 12384 11112 12436
rect 6184 12316 6236 12368
rect 6644 12316 6696 12368
rect 6920 12316 6972 12368
rect 7472 12316 7524 12368
rect 4896 12291 4948 12300
rect 4896 12257 4930 12291
rect 4930 12257 4948 12291
rect 8668 12291 8720 12300
rect 4896 12248 4948 12257
rect 1676 12180 1728 12232
rect 2964 12223 3016 12232
rect 2964 12189 2973 12223
rect 2973 12189 3007 12223
rect 3007 12189 3016 12223
rect 2964 12180 3016 12189
rect 4528 12180 4580 12232
rect 8668 12257 8677 12291
rect 8677 12257 8711 12291
rect 8711 12257 8720 12291
rect 8668 12248 8720 12257
rect 8760 12291 8812 12300
rect 8760 12257 8769 12291
rect 8769 12257 8803 12291
rect 8803 12257 8812 12291
rect 11244 12316 11296 12368
rect 8760 12248 8812 12257
rect 11704 12248 11756 12300
rect 12164 12248 12216 12300
rect 2504 12112 2556 12164
rect 2872 12044 2924 12096
rect 9128 12180 9180 12232
rect 9588 12180 9640 12232
rect 12072 12180 12124 12232
rect 12716 12248 12768 12300
rect 15384 12248 15436 12300
rect 16948 12248 17000 12300
rect 13820 12180 13872 12232
rect 12348 12112 12400 12164
rect 19156 12112 19208 12164
rect 6460 12044 6512 12096
rect 6736 12044 6788 12096
rect 7656 12044 7708 12096
rect 8392 12044 8444 12096
rect 12532 12044 12584 12096
rect 13452 12044 13504 12096
rect 14832 12044 14884 12096
rect 16120 12044 16172 12096
rect 17500 12044 17552 12096
rect 18236 12044 18288 12096
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 2780 11772 2832 11824
rect 4528 11840 4580 11892
rect 4896 11840 4948 11892
rect 9588 11840 9640 11892
rect 11060 11840 11112 11892
rect 11612 11840 11664 11892
rect 2504 11704 2556 11756
rect 7840 11772 7892 11824
rect 5540 11704 5592 11756
rect 6736 11704 6788 11756
rect 9128 11704 9180 11756
rect 12348 11704 12400 11756
rect 13636 11704 13688 11756
rect 17592 11840 17644 11892
rect 16212 11772 16264 11824
rect 19616 11772 19668 11824
rect 1860 11636 1912 11688
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 6368 11636 6420 11688
rect 6920 11636 6972 11688
rect 7472 11636 7524 11688
rect 7564 11636 7616 11688
rect 12164 11636 12216 11688
rect 15936 11704 15988 11756
rect 15108 11636 15160 11688
rect 17132 11704 17184 11756
rect 17868 11704 17920 11756
rect 18328 11704 18380 11756
rect 16488 11679 16540 11688
rect 16488 11645 16497 11679
rect 16497 11645 16531 11679
rect 16531 11645 16540 11679
rect 16488 11636 16540 11645
rect 3792 11568 3844 11620
rect 6736 11568 6788 11620
rect 1768 11543 1820 11552
rect 1768 11509 1777 11543
rect 1777 11509 1811 11543
rect 1811 11509 1820 11543
rect 1768 11500 1820 11509
rect 1860 11500 1912 11552
rect 2780 11543 2832 11552
rect 2780 11509 2789 11543
rect 2789 11509 2823 11543
rect 2823 11509 2832 11543
rect 5448 11543 5500 11552
rect 2780 11500 2832 11509
rect 5448 11509 5457 11543
rect 5457 11509 5491 11543
rect 5491 11509 5500 11543
rect 5448 11500 5500 11509
rect 5724 11500 5776 11552
rect 6000 11500 6052 11552
rect 6368 11500 6420 11552
rect 13544 11568 13596 11620
rect 14464 11568 14516 11620
rect 14648 11568 14700 11620
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 9036 11543 9088 11552
rect 9036 11509 9045 11543
rect 9045 11509 9079 11543
rect 9079 11509 9088 11543
rect 9036 11500 9088 11509
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 12440 11543 12492 11552
rect 12440 11509 12449 11543
rect 12449 11509 12483 11543
rect 12483 11509 12492 11543
rect 12440 11500 12492 11509
rect 13360 11500 13412 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 14096 11543 14148 11552
rect 14096 11509 14105 11543
rect 14105 11509 14139 11543
rect 14139 11509 14148 11543
rect 14096 11500 14148 11509
rect 14280 11500 14332 11552
rect 15108 11500 15160 11552
rect 16212 11500 16264 11552
rect 16580 11500 16632 11552
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 2780 11296 2832 11348
rect 2964 11296 3016 11348
rect 3240 11296 3292 11348
rect 3424 11296 3476 11348
rect 3516 11296 3568 11348
rect 4436 11339 4488 11348
rect 4436 11305 4445 11339
rect 4445 11305 4479 11339
rect 4479 11305 4488 11339
rect 4436 11296 4488 11305
rect 6092 11296 6144 11348
rect 6368 11296 6420 11348
rect 14648 11296 14700 11348
rect 15200 11296 15252 11348
rect 15568 11296 15620 11348
rect 5356 11228 5408 11280
rect 6276 11228 6328 11280
rect 5632 11160 5684 11212
rect 6644 11160 6696 11212
rect 1584 11092 1636 11144
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 3332 11135 3384 11144
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 3332 11092 3384 11101
rect 4896 11092 4948 11144
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 6000 11135 6052 11144
rect 6000 11101 6009 11135
rect 6009 11101 6043 11135
rect 6043 11101 6052 11135
rect 8208 11228 8260 11280
rect 7472 11135 7524 11144
rect 6000 11092 6052 11101
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 8760 11092 8812 11144
rect 10324 11092 10376 11144
rect 11336 11160 11388 11212
rect 13084 11228 13136 11280
rect 13544 11228 13596 11280
rect 14372 11160 14424 11212
rect 15200 11160 15252 11212
rect 16856 11203 16908 11212
rect 16856 11169 16865 11203
rect 16865 11169 16899 11203
rect 16899 11169 16908 11203
rect 16856 11160 16908 11169
rect 13544 11092 13596 11144
rect 13728 11092 13780 11144
rect 13912 11092 13964 11144
rect 15660 11092 15712 11144
rect 1676 10956 1728 11008
rect 5356 10999 5408 11008
rect 5356 10965 5365 10999
rect 5365 10965 5399 10999
rect 5399 10965 5408 10999
rect 5356 10956 5408 10965
rect 6552 11024 6604 11076
rect 8852 10999 8904 11008
rect 8852 10965 8861 10999
rect 8861 10965 8895 10999
rect 8895 10965 8904 10999
rect 8852 10956 8904 10965
rect 10416 10956 10468 11008
rect 11796 10956 11848 11008
rect 15568 11024 15620 11076
rect 16212 11092 16264 11144
rect 16396 11092 16448 11144
rect 16764 11092 16816 11144
rect 17040 11135 17092 11144
rect 17040 11101 17049 11135
rect 17049 11101 17083 11135
rect 17083 11101 17092 11135
rect 17040 11092 17092 11101
rect 18144 11024 18196 11076
rect 14648 10999 14700 11008
rect 14648 10965 14657 10999
rect 14657 10965 14691 10999
rect 14691 10965 14700 10999
rect 14648 10956 14700 10965
rect 15108 10956 15160 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 12256 10752 12308 10804
rect 12992 10795 13044 10804
rect 12992 10761 13001 10795
rect 13001 10761 13035 10795
rect 13035 10761 13044 10795
rect 12992 10752 13044 10761
rect 2412 10591 2464 10600
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 2504 10548 2556 10600
rect 4252 10684 4304 10736
rect 4528 10684 4580 10736
rect 5540 10684 5592 10736
rect 6644 10684 6696 10736
rect 3332 10480 3384 10532
rect 2780 10412 2832 10464
rect 3056 10412 3108 10464
rect 8852 10684 8904 10736
rect 7656 10616 7708 10668
rect 10416 10616 10468 10668
rect 11152 10659 11204 10668
rect 11152 10625 11161 10659
rect 11161 10625 11195 10659
rect 11195 10625 11204 10659
rect 11152 10616 11204 10625
rect 11336 10659 11388 10668
rect 11336 10625 11345 10659
rect 11345 10625 11379 10659
rect 11379 10625 11388 10659
rect 11336 10616 11388 10625
rect 5356 10548 5408 10600
rect 6736 10548 6788 10600
rect 7288 10548 7340 10600
rect 7932 10548 7984 10600
rect 10324 10548 10376 10600
rect 10784 10548 10836 10600
rect 11060 10591 11112 10600
rect 11060 10557 11069 10591
rect 11069 10557 11103 10591
rect 11103 10557 11112 10591
rect 11060 10548 11112 10557
rect 5264 10480 5316 10532
rect 13084 10616 13136 10668
rect 13728 10752 13780 10804
rect 12256 10548 12308 10600
rect 16028 10548 16080 10600
rect 16488 10548 16540 10600
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 4528 10412 4580 10464
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 5356 10412 5408 10464
rect 6184 10412 6236 10464
rect 7472 10412 7524 10464
rect 9496 10412 9548 10464
rect 10140 10412 10192 10464
rect 10324 10412 10376 10464
rect 10692 10455 10744 10464
rect 10692 10421 10701 10455
rect 10701 10421 10735 10455
rect 10735 10421 10744 10455
rect 10692 10412 10744 10421
rect 12348 10480 12400 10532
rect 15476 10480 15528 10532
rect 11796 10412 11848 10464
rect 13544 10412 13596 10464
rect 16672 10480 16724 10532
rect 16488 10412 16540 10464
rect 17040 10412 17092 10464
rect 17316 10412 17368 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 3056 10208 3108 10260
rect 3700 10208 3752 10260
rect 4896 10208 4948 10260
rect 5080 10208 5132 10260
rect 5448 10208 5500 10260
rect 5816 10208 5868 10260
rect 6368 10208 6420 10260
rect 6736 10208 6788 10260
rect 3792 10140 3844 10192
rect 5632 10140 5684 10192
rect 3056 10072 3108 10124
rect 2504 10004 2556 10056
rect 2964 10004 3016 10056
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 4160 10072 4212 10124
rect 5816 10072 5868 10124
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 7656 10072 7708 10124
rect 8300 10140 8352 10192
rect 12440 10208 12492 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 13912 10208 13964 10260
rect 15660 10208 15712 10260
rect 16856 10208 16908 10260
rect 8944 10140 8996 10192
rect 10692 10140 10744 10192
rect 11336 10115 11388 10124
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 5448 10004 5500 10013
rect 6000 10004 6052 10056
rect 6368 10004 6420 10056
rect 9404 10004 9456 10056
rect 4436 9936 4488 9988
rect 5356 9936 5408 9988
rect 5540 9936 5592 9988
rect 7288 9936 7340 9988
rect 9680 9936 9732 9988
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 14464 10140 14516 10192
rect 15108 10140 15160 10192
rect 15292 10140 15344 10192
rect 18420 10208 18472 10260
rect 10324 10004 10376 10013
rect 11796 10004 11848 10056
rect 12256 10004 12308 10056
rect 12440 10004 12492 10056
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 14648 10115 14700 10124
rect 14648 10081 14666 10115
rect 14666 10081 14700 10115
rect 14648 10072 14700 10081
rect 17132 10072 17184 10124
rect 17224 10072 17276 10124
rect 13544 10004 13596 10056
rect 16304 10047 16356 10056
rect 16304 10013 16313 10047
rect 16313 10013 16347 10047
rect 16347 10013 16356 10047
rect 16304 10004 16356 10013
rect 16488 10047 16540 10056
rect 16488 10013 16497 10047
rect 16497 10013 16531 10047
rect 16531 10013 16540 10047
rect 16488 10004 16540 10013
rect 17776 10047 17828 10056
rect 17776 10013 17785 10047
rect 17785 10013 17819 10047
rect 17819 10013 17828 10047
rect 17776 10004 17828 10013
rect 8944 9911 8996 9920
rect 8944 9877 8953 9911
rect 8953 9877 8987 9911
rect 8987 9877 8996 9911
rect 8944 9868 8996 9877
rect 10692 9868 10744 9920
rect 13728 9868 13780 9920
rect 18512 9868 18564 9920
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 3056 9664 3108 9716
rect 4896 9664 4948 9716
rect 5448 9707 5500 9716
rect 5448 9673 5457 9707
rect 5457 9673 5491 9707
rect 5491 9673 5500 9707
rect 5448 9664 5500 9673
rect 9128 9596 9180 9648
rect 10600 9664 10652 9716
rect 10968 9664 11020 9716
rect 12624 9664 12676 9716
rect 15568 9664 15620 9716
rect 9680 9596 9732 9648
rect 3332 9528 3384 9580
rect 6368 9528 6420 9580
rect 8944 9528 8996 9580
rect 1584 9460 1636 9512
rect 2412 9460 2464 9512
rect 4068 9460 4120 9512
rect 5356 9503 5408 9512
rect 5356 9469 5365 9503
rect 5365 9469 5399 9503
rect 5399 9469 5408 9503
rect 5356 9460 5408 9469
rect 2964 9392 3016 9444
rect 4160 9435 4212 9444
rect 4160 9401 4169 9435
rect 4169 9401 4203 9435
rect 4203 9401 4212 9435
rect 4160 9392 4212 9401
rect 6736 9392 6788 9444
rect 5080 9324 5132 9376
rect 5264 9324 5316 9376
rect 5908 9367 5960 9376
rect 5908 9333 5917 9367
rect 5917 9333 5951 9367
rect 5951 9333 5960 9367
rect 5908 9324 5960 9333
rect 6184 9324 6236 9376
rect 6644 9324 6696 9376
rect 11336 9596 11388 9648
rect 11520 9596 11572 9648
rect 11704 9596 11756 9648
rect 13636 9596 13688 9648
rect 16764 9639 16816 9648
rect 16764 9605 16773 9639
rect 16773 9605 16807 9639
rect 16807 9605 16816 9639
rect 16764 9596 16816 9605
rect 11152 9528 11204 9580
rect 12348 9528 12400 9580
rect 13820 9528 13872 9580
rect 17224 9528 17276 9580
rect 11888 9460 11940 9512
rect 12072 9503 12124 9512
rect 12072 9469 12081 9503
rect 12081 9469 12115 9503
rect 12115 9469 12124 9503
rect 12072 9460 12124 9469
rect 12808 9460 12860 9512
rect 7564 9392 7616 9444
rect 9404 9392 9456 9444
rect 12164 9435 12216 9444
rect 12164 9401 12173 9435
rect 12173 9401 12207 9435
rect 12207 9401 12216 9435
rect 12164 9392 12216 9401
rect 12348 9392 12400 9444
rect 8484 9324 8536 9376
rect 9312 9367 9364 9376
rect 9312 9333 9321 9367
rect 9321 9333 9355 9367
rect 9355 9333 9364 9367
rect 9312 9324 9364 9333
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 10416 9324 10468 9376
rect 11060 9367 11112 9376
rect 11060 9333 11069 9367
rect 11069 9333 11103 9367
rect 11103 9333 11112 9367
rect 11060 9324 11112 9333
rect 11520 9324 11572 9376
rect 11704 9324 11756 9376
rect 12716 9324 12768 9376
rect 13360 9324 13412 9376
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 16488 9460 16540 9512
rect 16672 9460 16724 9512
rect 17776 9528 17828 9580
rect 16120 9392 16172 9444
rect 17224 9435 17276 9444
rect 17224 9401 17233 9435
rect 17233 9401 17267 9435
rect 17267 9401 17276 9435
rect 17224 9392 17276 9401
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 5908 9163 5960 9172
rect 2136 9052 2188 9104
rect 5908 9129 5917 9163
rect 5917 9129 5951 9163
rect 5951 9129 5960 9163
rect 5908 9120 5960 9129
rect 6368 9163 6420 9172
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 6736 9120 6788 9172
rect 7288 9120 7340 9172
rect 9036 9120 9088 9172
rect 11060 9120 11112 9172
rect 11152 9120 11204 9172
rect 11336 9120 11388 9172
rect 13360 9120 13412 9172
rect 13820 9120 13872 9172
rect 16672 9163 16724 9172
rect 5816 9052 5868 9104
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 4344 9027 4396 9036
rect 4344 8993 4378 9027
rect 4378 8993 4396 9027
rect 4344 8984 4396 8993
rect 5908 8984 5960 9036
rect 11520 9052 11572 9104
rect 11704 9052 11756 9104
rect 8208 8984 8260 9036
rect 9036 8984 9088 9036
rect 9128 8984 9180 9036
rect 10692 8984 10744 9036
rect 10784 8984 10836 9036
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 6460 8916 6512 8968
rect 6644 8916 6696 8968
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 9680 8916 9732 8968
rect 11612 8984 11664 9036
rect 13820 8984 13872 9036
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 17132 9163 17184 9172
rect 17132 9129 17141 9163
rect 17141 9129 17175 9163
rect 17175 9129 17184 9163
rect 17132 9120 17184 9129
rect 17224 9120 17276 9172
rect 15660 9052 15712 9104
rect 17592 9052 17644 9104
rect 5172 8780 5224 8832
rect 6460 8780 6512 8832
rect 10048 8848 10100 8900
rect 13084 8916 13136 8968
rect 10784 8780 10836 8832
rect 10968 8848 11020 8900
rect 12164 8780 12216 8832
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 15384 8984 15436 9036
rect 17592 8959 17644 8968
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 17776 8959 17828 8968
rect 17776 8925 17785 8959
rect 17785 8925 17819 8959
rect 17819 8925 17828 8959
rect 17776 8916 17828 8925
rect 13820 8780 13872 8832
rect 14464 8780 14516 8832
rect 17776 8780 17828 8832
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 2044 8576 2096 8628
rect 5356 8576 5408 8628
rect 12072 8576 12124 8628
rect 12716 8576 12768 8628
rect 15660 8576 15712 8628
rect 16212 8576 16264 8628
rect 16304 8576 16356 8628
rect 1584 8508 1636 8560
rect 4344 8508 4396 8560
rect 2964 8440 3016 8492
rect 3332 8440 3384 8492
rect 4252 8440 4304 8492
rect 5172 8440 5224 8492
rect 6000 8440 6052 8492
rect 9312 8508 9364 8560
rect 10048 8508 10100 8560
rect 11612 8508 11664 8560
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 9680 8440 9732 8492
rect 11520 8440 11572 8492
rect 14004 8508 14056 8560
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 13912 8440 13964 8492
rect 16672 8440 16724 8492
rect 3424 8415 3476 8424
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 1492 8304 1544 8356
rect 2964 8304 3016 8356
rect 3608 8372 3660 8424
rect 4712 8372 4764 8424
rect 7288 8372 7340 8424
rect 7380 8372 7432 8424
rect 8576 8415 8628 8424
rect 4252 8304 4304 8356
rect 5908 8347 5960 8356
rect 5908 8313 5917 8347
rect 5917 8313 5951 8347
rect 5951 8313 5960 8347
rect 5908 8304 5960 8313
rect 6368 8304 6420 8356
rect 7656 8304 7708 8356
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 9404 8372 9456 8424
rect 10692 8415 10744 8424
rect 10140 8304 10192 8356
rect 10692 8381 10726 8415
rect 10726 8381 10744 8415
rect 10692 8372 10744 8381
rect 12348 8372 12400 8424
rect 12716 8372 12768 8424
rect 15752 8372 15804 8424
rect 16212 8372 16264 8424
rect 15108 8304 15160 8356
rect 16672 8304 16724 8356
rect 2228 8279 2280 8288
rect 2228 8245 2237 8279
rect 2237 8245 2271 8279
rect 2271 8245 2280 8279
rect 2228 8236 2280 8245
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 4712 8279 4764 8288
rect 4712 8245 4721 8279
rect 4721 8245 4755 8279
rect 4755 8245 4764 8279
rect 5540 8279 5592 8288
rect 4712 8236 4764 8245
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 5540 8236 5592 8245
rect 7564 8236 7616 8288
rect 11612 8236 11664 8288
rect 12072 8236 12124 8288
rect 12256 8236 12308 8288
rect 13544 8236 13596 8288
rect 15384 8236 15436 8288
rect 16764 8279 16816 8288
rect 16764 8245 16773 8279
rect 16773 8245 16807 8279
rect 16807 8245 16816 8279
rect 16764 8236 16816 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 5540 8032 5592 8084
rect 2044 7964 2096 8016
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 3608 7964 3660 8016
rect 5448 7896 5500 7948
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 5172 7871 5224 7880
rect 3332 7828 3384 7837
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 7380 8032 7432 8084
rect 6184 7964 6236 8016
rect 10140 8032 10192 8084
rect 11520 8032 11572 8084
rect 11888 8032 11940 8084
rect 16764 8032 16816 8084
rect 17592 8032 17644 8084
rect 6000 7939 6052 7948
rect 6000 7905 6034 7939
rect 6034 7905 6052 7939
rect 6000 7896 6052 7905
rect 6368 7896 6420 7948
rect 7196 7896 7248 7948
rect 8484 7896 8536 7948
rect 11060 7964 11112 8016
rect 13084 7964 13136 8016
rect 15292 7964 15344 8016
rect 15476 7964 15528 8016
rect 9588 7896 9640 7948
rect 12072 7939 12124 7948
rect 12072 7905 12081 7939
rect 12081 7905 12115 7939
rect 12115 7905 12124 7939
rect 12072 7896 12124 7905
rect 5172 7828 5224 7837
rect 9680 7871 9732 7880
rect 4620 7760 4672 7812
rect 2596 7692 2648 7744
rect 5448 7692 5500 7744
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 11060 7828 11112 7880
rect 11336 7828 11388 7880
rect 11612 7828 11664 7880
rect 8484 7760 8536 7812
rect 9128 7760 9180 7812
rect 10692 7692 10744 7744
rect 11612 7692 11664 7744
rect 12348 7828 12400 7880
rect 12900 7803 12952 7812
rect 12900 7769 12909 7803
rect 12909 7769 12943 7803
rect 12943 7769 12952 7803
rect 12900 7760 12952 7769
rect 14004 7896 14056 7948
rect 15016 7896 15068 7948
rect 17868 7964 17920 8016
rect 13084 7692 13136 7744
rect 15292 7692 15344 7744
rect 15660 7760 15712 7812
rect 17224 7760 17276 7812
rect 17868 7692 17920 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 4252 7488 4304 7540
rect 4712 7488 4764 7540
rect 5540 7531 5592 7540
rect 5540 7497 5549 7531
rect 5549 7497 5583 7531
rect 5583 7497 5592 7531
rect 5540 7488 5592 7497
rect 7196 7531 7248 7540
rect 7196 7497 7205 7531
rect 7205 7497 7239 7531
rect 7239 7497 7248 7531
rect 7196 7488 7248 7497
rect 8024 7488 8076 7540
rect 9588 7488 9640 7540
rect 2136 7352 2188 7404
rect 4896 7352 4948 7404
rect 5080 7352 5132 7404
rect 6644 7420 6696 7472
rect 6368 7352 6420 7404
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 3056 7284 3108 7336
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 5816 7284 5868 7336
rect 8208 7420 8260 7472
rect 8024 7352 8076 7404
rect 12348 7488 12400 7540
rect 8300 7284 8352 7336
rect 9220 7284 9272 7336
rect 9680 7284 9732 7336
rect 4160 7216 4212 7268
rect 3424 7148 3476 7200
rect 3608 7191 3660 7200
rect 3608 7157 3617 7191
rect 3617 7157 3651 7191
rect 3651 7157 3660 7191
rect 3608 7148 3660 7157
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 8484 7216 8536 7268
rect 8576 7216 8628 7268
rect 4712 7148 4764 7157
rect 8208 7148 8260 7200
rect 12072 7352 12124 7404
rect 12900 7352 12952 7404
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 11060 7284 11112 7336
rect 13176 7284 13228 7336
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12992 7216 13044 7268
rect 12440 7148 12492 7157
rect 13176 7148 13228 7200
rect 13912 7488 13964 7540
rect 15108 7531 15160 7540
rect 15108 7497 15117 7531
rect 15117 7497 15151 7531
rect 15151 7497 15160 7531
rect 15108 7488 15160 7497
rect 15016 7148 15068 7200
rect 16120 7216 16172 7268
rect 16488 7148 16540 7200
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 4160 6944 4212 6996
rect 4712 6944 4764 6996
rect 4988 6944 5040 6996
rect 5080 6944 5132 6996
rect 6000 6944 6052 6996
rect 8116 6944 8168 6996
rect 3148 6919 3200 6928
rect 3148 6885 3157 6919
rect 3157 6885 3191 6919
rect 3191 6885 3200 6919
rect 3148 6876 3200 6885
rect 3792 6808 3844 6860
rect 5908 6876 5960 6928
rect 9496 6876 9548 6928
rect 13636 6944 13688 6996
rect 14096 6944 14148 6996
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 16580 6944 16632 6996
rect 16856 6876 16908 6928
rect 5816 6808 5868 6860
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 8024 6808 8076 6860
rect 3056 6740 3108 6792
rect 3884 6740 3936 6792
rect 2412 6672 2464 6724
rect 2964 6604 3016 6656
rect 4252 6604 4304 6656
rect 5448 6604 5500 6656
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 6000 6604 6052 6656
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 8852 6783 8904 6792
rect 7656 6740 7708 6749
rect 8852 6749 8861 6783
rect 8861 6749 8895 6783
rect 8895 6749 8904 6783
rect 8852 6740 8904 6749
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 10508 6808 10560 6860
rect 11520 6808 11572 6860
rect 8944 6740 8996 6749
rect 10692 6740 10744 6792
rect 10968 6783 11020 6792
rect 10968 6749 10977 6783
rect 10977 6749 11011 6783
rect 11011 6749 11020 6783
rect 12440 6808 12492 6860
rect 13176 6808 13228 6860
rect 12256 6783 12308 6792
rect 10968 6740 11020 6749
rect 8116 6672 8168 6724
rect 10416 6715 10468 6724
rect 8484 6604 8536 6656
rect 9680 6604 9732 6656
rect 10416 6681 10425 6715
rect 10425 6681 10459 6715
rect 10459 6681 10468 6715
rect 10416 6672 10468 6681
rect 12256 6749 12265 6783
rect 12265 6749 12299 6783
rect 12299 6749 12308 6783
rect 12256 6740 12308 6749
rect 13084 6740 13136 6792
rect 17408 6808 17460 6860
rect 13820 6740 13872 6792
rect 14648 6783 14700 6792
rect 14648 6749 14657 6783
rect 14657 6749 14691 6783
rect 14691 6749 14700 6783
rect 14648 6740 14700 6749
rect 15476 6740 15528 6792
rect 11520 6604 11572 6656
rect 14004 6647 14056 6656
rect 14004 6613 14013 6647
rect 14013 6613 14047 6647
rect 14047 6613 14056 6647
rect 14004 6604 14056 6613
rect 15108 6672 15160 6724
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 16672 6715 16724 6724
rect 16672 6681 16681 6715
rect 16681 6681 16715 6715
rect 16715 6681 16724 6715
rect 16672 6672 16724 6681
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 3792 6443 3844 6452
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 3792 6409 3801 6443
rect 3801 6409 3835 6443
rect 3835 6409 3844 6443
rect 3792 6400 3844 6409
rect 5264 6400 5316 6452
rect 6276 6400 6328 6452
rect 7748 6400 7800 6452
rect 8300 6400 8352 6452
rect 12164 6400 12216 6452
rect 12716 6400 12768 6452
rect 4436 6264 4488 6316
rect 4252 6196 4304 6248
rect 4712 6196 4764 6248
rect 6276 6196 6328 6248
rect 10968 6332 11020 6384
rect 13636 6332 13688 6384
rect 2596 6128 2648 6180
rect 1860 6103 1912 6112
rect 1860 6069 1869 6103
rect 1869 6069 1903 6103
rect 1903 6069 1912 6103
rect 1860 6060 1912 6069
rect 6000 6103 6052 6112
rect 6000 6069 6009 6103
rect 6009 6069 6043 6103
rect 6043 6069 6052 6103
rect 6000 6060 6052 6069
rect 6184 6060 6236 6112
rect 6736 6060 6788 6112
rect 7656 6264 7708 6316
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 9220 6307 9272 6316
rect 8576 6264 8628 6273
rect 9220 6273 9229 6307
rect 9229 6273 9263 6307
rect 9263 6273 9272 6307
rect 9220 6264 9272 6273
rect 11612 6307 11664 6316
rect 11612 6273 11621 6307
rect 11621 6273 11655 6307
rect 11655 6273 11664 6307
rect 11612 6264 11664 6273
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 11888 6264 11940 6316
rect 14740 6400 14792 6452
rect 15660 6400 15712 6452
rect 16120 6332 16172 6384
rect 17132 6332 17184 6384
rect 14004 6264 14056 6316
rect 16488 6307 16540 6316
rect 8760 6196 8812 6248
rect 10324 6196 10376 6248
rect 11520 6239 11572 6248
rect 11520 6205 11529 6239
rect 11529 6205 11563 6239
rect 11563 6205 11572 6239
rect 11520 6196 11572 6205
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 16488 6273 16497 6307
rect 16497 6273 16531 6307
rect 16531 6273 16540 6307
rect 16488 6264 16540 6273
rect 16856 6264 16908 6316
rect 17040 6264 17092 6316
rect 17132 6196 17184 6248
rect 7380 6128 7432 6180
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 8392 6103 8444 6112
rect 8392 6069 8401 6103
rect 8401 6069 8435 6103
rect 8435 6069 8444 6103
rect 8392 6060 8444 6069
rect 9128 6128 9180 6180
rect 13176 6128 13228 6180
rect 14648 6128 14700 6180
rect 15200 6128 15252 6180
rect 16672 6128 16724 6180
rect 17316 6060 17368 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 4436 5856 4488 5908
rect 5632 5856 5684 5908
rect 6276 5856 6328 5908
rect 6736 5856 6788 5908
rect 7288 5856 7340 5908
rect 1768 5652 1820 5704
rect 3792 5652 3844 5704
rect 5908 5788 5960 5840
rect 7380 5788 7432 5840
rect 9128 5831 9180 5840
rect 4436 5763 4488 5772
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 9128 5797 9137 5831
rect 9137 5797 9171 5831
rect 9171 5797 9180 5831
rect 9128 5788 9180 5797
rect 9312 5856 9364 5908
rect 10968 5856 11020 5908
rect 11796 5856 11848 5908
rect 12164 5788 12216 5840
rect 16764 5856 16816 5908
rect 17316 5899 17368 5908
rect 17316 5865 17325 5899
rect 17325 5865 17359 5899
rect 17359 5865 17368 5899
rect 17316 5856 17368 5865
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 16120 5788 16172 5840
rect 9496 5720 9548 5772
rect 12256 5720 12308 5772
rect 3792 5516 3844 5568
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 6184 5652 6236 5704
rect 9036 5652 9088 5704
rect 9220 5652 9272 5704
rect 9588 5652 9640 5704
rect 10968 5652 11020 5704
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 8484 5584 8536 5636
rect 9312 5584 9364 5636
rect 9128 5516 9180 5568
rect 10416 5516 10468 5568
rect 14096 5720 14148 5772
rect 15660 5720 15712 5772
rect 17500 5788 17552 5840
rect 18328 5788 18380 5840
rect 16580 5695 16632 5704
rect 16580 5661 16589 5695
rect 16589 5661 16623 5695
rect 16623 5661 16632 5695
rect 16580 5652 16632 5661
rect 17040 5652 17092 5704
rect 18972 5695 19024 5704
rect 18972 5661 18981 5695
rect 18981 5661 19015 5695
rect 19015 5661 19024 5695
rect 18972 5652 19024 5661
rect 15200 5516 15252 5568
rect 15660 5516 15712 5568
rect 16120 5559 16172 5568
rect 16120 5525 16129 5559
rect 16129 5525 16163 5559
rect 16163 5525 16172 5559
rect 16120 5516 16172 5525
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 1860 5355 1912 5364
rect 1860 5321 1869 5355
rect 1869 5321 1903 5355
rect 1903 5321 1912 5355
rect 1860 5312 1912 5321
rect 4436 5312 4488 5364
rect 8300 5312 8352 5364
rect 9496 5355 9548 5364
rect 9496 5321 9505 5355
rect 9505 5321 9539 5355
rect 9539 5321 9548 5355
rect 9496 5312 9548 5321
rect 9588 5312 9640 5364
rect 6276 5287 6328 5296
rect 1676 5151 1728 5160
rect 1676 5117 1685 5151
rect 1685 5117 1719 5151
rect 1719 5117 1728 5151
rect 1676 5108 1728 5117
rect 6276 5253 6285 5287
rect 6285 5253 6319 5287
rect 6319 5253 6328 5287
rect 6276 5244 6328 5253
rect 6368 5244 6420 5296
rect 2872 5176 2924 5228
rect 3240 5176 3292 5228
rect 4712 5176 4764 5228
rect 3332 5108 3384 5160
rect 4252 5108 4304 5160
rect 6184 5108 6236 5160
rect 6736 5108 6788 5160
rect 7380 5108 7432 5160
rect 7748 5108 7800 5160
rect 9864 5108 9916 5160
rect 2872 5083 2924 5092
rect 2872 5049 2881 5083
rect 2881 5049 2915 5083
rect 2915 5049 2924 5083
rect 2872 5040 2924 5049
rect 5080 5040 5132 5092
rect 9036 5040 9088 5092
rect 11704 5312 11756 5364
rect 13544 5312 13596 5364
rect 13820 5312 13872 5364
rect 15476 5355 15528 5364
rect 15476 5321 15485 5355
rect 15485 5321 15519 5355
rect 15519 5321 15528 5355
rect 15476 5312 15528 5321
rect 16672 5355 16724 5364
rect 16672 5321 16681 5355
rect 16681 5321 16715 5355
rect 16715 5321 16724 5355
rect 16672 5312 16724 5321
rect 16304 5244 16356 5296
rect 13636 5176 13688 5228
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 16488 5176 16540 5228
rect 17040 5176 17092 5228
rect 10968 5108 11020 5160
rect 12716 5108 12768 5160
rect 16120 5108 16172 5160
rect 17316 5108 17368 5160
rect 10416 5040 10468 5092
rect 11152 5040 11204 5092
rect 11704 5040 11756 5092
rect 13360 5040 13412 5092
rect 5632 4972 5684 5024
rect 6000 4972 6052 5024
rect 9404 4972 9456 5024
rect 10784 4972 10836 5024
rect 15936 5015 15988 5024
rect 15936 4981 15945 5015
rect 15945 4981 15979 5015
rect 15979 4981 15988 5015
rect 15936 4972 15988 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 1860 4811 1912 4820
rect 1860 4777 1869 4811
rect 1869 4777 1903 4811
rect 1903 4777 1912 4811
rect 1860 4768 1912 4777
rect 2780 4768 2832 4820
rect 4804 4768 4856 4820
rect 5356 4768 5408 4820
rect 5632 4811 5684 4820
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 3240 4700 3292 4752
rect 2412 4675 2464 4684
rect 2412 4641 2421 4675
rect 2421 4641 2455 4675
rect 2455 4641 2464 4675
rect 2412 4632 2464 4641
rect 5172 4632 5224 4684
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 8852 4768 8904 4820
rect 9036 4811 9088 4820
rect 9036 4777 9045 4811
rect 9045 4777 9079 4811
rect 9079 4777 9088 4811
rect 9036 4768 9088 4777
rect 11060 4768 11112 4820
rect 6000 4743 6052 4752
rect 6000 4709 6009 4743
rect 6009 4709 6043 4743
rect 6043 4709 6052 4743
rect 11152 4743 11204 4752
rect 6000 4700 6052 4709
rect 11152 4709 11161 4743
rect 11161 4709 11195 4743
rect 11195 4709 11204 4743
rect 11152 4700 11204 4709
rect 11980 4743 12032 4752
rect 11980 4709 11989 4743
rect 11989 4709 12023 4743
rect 12023 4709 12032 4743
rect 11980 4700 12032 4709
rect 12072 4743 12124 4752
rect 12072 4709 12081 4743
rect 12081 4709 12115 4743
rect 12115 4709 12124 4743
rect 12072 4700 12124 4709
rect 12440 4700 12492 4752
rect 13820 4743 13872 4752
rect 13820 4709 13829 4743
rect 13829 4709 13863 4743
rect 13863 4709 13872 4743
rect 13820 4700 13872 4709
rect 15108 4700 15160 4752
rect 15936 4768 15988 4820
rect 17132 4768 17184 4820
rect 16396 4743 16448 4752
rect 5448 4496 5500 4548
rect 6276 4564 6328 4616
rect 7748 4632 7800 4684
rect 8484 4632 8536 4684
rect 8852 4632 8904 4684
rect 10784 4675 10836 4684
rect 10784 4641 10793 4675
rect 10793 4641 10827 4675
rect 10827 4641 10836 4675
rect 10784 4632 10836 4641
rect 16396 4709 16405 4743
rect 16405 4709 16439 4743
rect 16439 4709 16448 4743
rect 16396 4700 16448 4709
rect 16764 4632 16816 4684
rect 17040 4632 17092 4684
rect 9864 4564 9916 4616
rect 10508 4564 10560 4616
rect 14372 4607 14424 4616
rect 8944 4496 8996 4548
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 15384 4607 15436 4616
rect 15384 4573 15393 4607
rect 15393 4573 15427 4607
rect 15427 4573 15436 4607
rect 15384 4564 15436 4573
rect 17316 4607 17368 4616
rect 17316 4573 17325 4607
rect 17325 4573 17359 4607
rect 17359 4573 17368 4607
rect 17316 4564 17368 4573
rect 14280 4496 14332 4548
rect 3240 4428 3292 4480
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 9588 4428 9640 4480
rect 11796 4428 11848 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 1860 4267 1912 4276
rect 1860 4233 1869 4267
rect 1869 4233 1903 4267
rect 1903 4233 1912 4267
rect 1860 4224 1912 4233
rect 3332 4224 3384 4276
rect 4436 4131 4488 4140
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 4712 4156 4764 4208
rect 4988 4224 5040 4276
rect 6000 4224 6052 4276
rect 5448 4156 5500 4208
rect 11060 4224 11112 4276
rect 2136 3995 2188 4004
rect 2136 3961 2145 3995
rect 2145 3961 2179 3995
rect 2179 3961 2188 3995
rect 2136 3952 2188 3961
rect 4712 4020 4764 4072
rect 4804 4020 4856 4072
rect 5356 4020 5408 4072
rect 8392 4156 8444 4208
rect 8944 4156 8996 4208
rect 6276 4088 6328 4140
rect 10324 4156 10376 4208
rect 3056 3952 3108 4004
rect 3884 3952 3936 4004
rect 7840 4020 7892 4072
rect 13176 4088 13228 4140
rect 13360 4131 13412 4140
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 15936 4088 15988 4140
rect 16948 4131 17000 4140
rect 16948 4097 16957 4131
rect 16957 4097 16991 4131
rect 16991 4097 17000 4131
rect 16948 4088 17000 4097
rect 7288 3952 7340 4004
rect 10048 4020 10100 4072
rect 10968 4020 11020 4072
rect 10416 3952 10468 4004
rect 10784 3952 10836 4004
rect 12532 3952 12584 4004
rect 14096 3952 14148 4004
rect 14556 3995 14608 4004
rect 14556 3961 14565 3995
rect 14565 3961 14599 3995
rect 14599 3961 14608 3995
rect 14556 3952 14608 3961
rect 15936 3952 15988 4004
rect 2780 3884 2832 3936
rect 3332 3927 3384 3936
rect 3332 3893 3341 3927
rect 3341 3893 3375 3927
rect 3375 3893 3384 3927
rect 3332 3884 3384 3893
rect 3792 3884 3844 3936
rect 5264 3884 5316 3936
rect 6460 3884 6512 3936
rect 8484 3884 8536 3936
rect 10968 3884 11020 3936
rect 15200 3884 15252 3936
rect 15752 3884 15804 3936
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 4896 3680 4948 3732
rect 5448 3723 5500 3732
rect 5448 3689 5457 3723
rect 5457 3689 5491 3723
rect 5491 3689 5500 3723
rect 5448 3680 5500 3689
rect 3884 3544 3936 3596
rect 4252 3612 4304 3664
rect 4436 3612 4488 3664
rect 5080 3612 5132 3664
rect 4620 3544 4672 3596
rect 6276 3680 6328 3732
rect 7288 3723 7340 3732
rect 7288 3689 7297 3723
rect 7297 3689 7331 3723
rect 7331 3689 7340 3723
rect 7288 3680 7340 3689
rect 8668 3680 8720 3732
rect 7380 3612 7432 3664
rect 7656 3612 7708 3664
rect 6460 3544 6512 3596
rect 8944 3612 8996 3664
rect 9220 3612 9272 3664
rect 10600 3612 10652 3664
rect 10784 3612 10836 3664
rect 11428 3655 11480 3664
rect 11428 3621 11437 3655
rect 11437 3621 11471 3655
rect 11471 3621 11480 3655
rect 11428 3612 11480 3621
rect 12348 3655 12400 3664
rect 12348 3621 12357 3655
rect 12357 3621 12391 3655
rect 12391 3621 12400 3655
rect 12348 3612 12400 3621
rect 8392 3587 8444 3596
rect 8392 3553 8401 3587
rect 8401 3553 8435 3587
rect 8435 3553 8444 3587
rect 8392 3544 8444 3553
rect 9036 3544 9088 3596
rect 9588 3544 9640 3596
rect 10324 3544 10376 3596
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 10968 3544 11020 3596
rect 12256 3544 12308 3596
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 7196 3476 7248 3528
rect 11060 3476 11112 3528
rect 11612 3476 11664 3528
rect 13544 3612 13596 3664
rect 14648 3680 14700 3732
rect 15384 3680 15436 3732
rect 15844 3723 15896 3732
rect 15844 3689 15853 3723
rect 15853 3689 15887 3723
rect 15887 3689 15896 3723
rect 15844 3680 15896 3689
rect 16580 3680 16632 3732
rect 16764 3680 16816 3732
rect 17316 3612 17368 3664
rect 13820 3544 13872 3596
rect 15384 3544 15436 3596
rect 15476 3544 15528 3596
rect 17040 3587 17092 3596
rect 17040 3553 17049 3587
rect 17049 3553 17083 3587
rect 17083 3553 17092 3587
rect 17040 3544 17092 3553
rect 17868 3680 17920 3732
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 15752 3476 15804 3528
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 7748 3408 7800 3460
rect 9956 3408 10008 3460
rect 10048 3451 10100 3460
rect 10048 3417 10057 3451
rect 10057 3417 10091 3451
rect 10091 3417 10100 3451
rect 10048 3408 10100 3417
rect 12624 3408 12676 3460
rect 14372 3408 14424 3460
rect 5172 3340 5224 3392
rect 10416 3340 10468 3392
rect 11704 3340 11756 3392
rect 15200 3340 15252 3392
rect 15384 3340 15436 3392
rect 16396 3340 16448 3392
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 7656 3136 7708 3188
rect 204 3000 256 3052
rect 1768 3000 1820 3052
rect 1584 2932 1636 2984
rect 3792 2932 3844 2984
rect 4528 3000 4580 3052
rect 664 2864 716 2916
rect 2136 2864 2188 2916
rect 3148 2864 3200 2916
rect 6460 3068 6512 3120
rect 12256 3136 12308 3188
rect 12348 3136 12400 3188
rect 17040 3136 17092 3188
rect 7564 3000 7616 3052
rect 11152 3068 11204 3120
rect 11428 3068 11480 3120
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 10876 3000 10928 3052
rect 11244 3043 11296 3052
rect 11244 3009 11253 3043
rect 11253 3009 11287 3043
rect 11287 3009 11296 3043
rect 11244 3000 11296 3009
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 13084 3000 13136 3052
rect 14556 3000 14608 3052
rect 14740 3000 14792 3052
rect 5356 2932 5408 2984
rect 6736 2932 6788 2984
rect 7288 2932 7340 2984
rect 8668 2932 8720 2984
rect 15568 3000 15620 3052
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 1676 2796 1728 2848
rect 7564 2864 7616 2916
rect 4712 2796 4764 2848
rect 7748 2796 7800 2848
rect 8668 2796 8720 2848
rect 9772 2864 9824 2916
rect 10508 2907 10560 2916
rect 10508 2873 10517 2907
rect 10517 2873 10551 2907
rect 10551 2873 10560 2907
rect 10508 2864 10560 2873
rect 10784 2864 10836 2916
rect 13084 2864 13136 2916
rect 10600 2796 10652 2848
rect 10692 2796 10744 2848
rect 14372 2907 14424 2916
rect 14372 2873 14381 2907
rect 14381 2873 14415 2907
rect 14415 2873 14424 2907
rect 14372 2864 14424 2873
rect 14832 2864 14884 2916
rect 15660 2864 15712 2916
rect 15936 2907 15988 2916
rect 15936 2873 15945 2907
rect 15945 2873 15979 2907
rect 15979 2873 15988 2907
rect 15936 2864 15988 2873
rect 14556 2796 14608 2848
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 2780 2592 2832 2644
rect 8116 2592 8168 2644
rect 15200 2592 15252 2644
rect 17684 2635 17736 2644
rect 17684 2601 17693 2635
rect 17693 2601 17727 2635
rect 17727 2601 17736 2635
rect 17684 2592 17736 2601
rect 3516 2524 3568 2576
rect 10232 2567 10284 2576
rect 1124 2388 1176 2440
rect 4804 2456 4856 2508
rect 7196 2456 7248 2508
rect 7380 2456 7432 2508
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 4988 2388 5040 2440
rect 4436 2320 4488 2372
rect 7564 2388 7616 2440
rect 7932 2388 7984 2440
rect 6736 2320 6788 2372
rect 8392 2388 8444 2440
rect 10232 2533 10241 2567
rect 10241 2533 10275 2567
rect 10275 2533 10284 2567
rect 10232 2524 10284 2533
rect 10416 2524 10468 2576
rect 11336 2524 11388 2576
rect 13452 2524 13504 2576
rect 14280 2567 14332 2576
rect 14280 2533 14289 2567
rect 14289 2533 14323 2567
rect 14323 2533 14332 2567
rect 14280 2524 14332 2533
rect 15016 2524 15068 2576
rect 11704 2456 11756 2508
rect 12532 2388 12584 2440
rect 12624 2388 12676 2440
rect 9772 2320 9824 2372
rect 3424 2295 3476 2304
rect 3424 2261 3433 2295
rect 3433 2261 3467 2295
rect 3467 2261 3476 2295
rect 3424 2252 3476 2261
rect 3516 2252 3568 2304
rect 10508 2252 10560 2304
rect 17776 2456 17828 2508
rect 15108 2388 15160 2440
rect 16488 2431 16540 2440
rect 16488 2397 16497 2431
rect 16497 2397 16531 2431
rect 16531 2397 16540 2431
rect 16488 2388 16540 2397
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 7932 1980 7984 2032
rect 10416 1980 10468 2032
rect 14556 1980 14608 2032
rect 13912 1368 13964 1420
rect 16672 1368 16724 1420
<< metal2 >>
rect 294 16520 350 17000
rect 938 16520 994 17000
rect 1582 16520 1638 17000
rect 2226 16520 2282 17000
rect 2870 16520 2926 17000
rect 3514 16520 3570 17000
rect 3698 16688 3754 16697
rect 3698 16623 3754 16632
rect 308 13530 336 16520
rect 952 14618 980 16520
rect 940 14612 992 14618
rect 940 14554 992 14560
rect 1596 14074 1624 16520
rect 2240 14618 2268 16520
rect 2594 16280 2650 16289
rect 2594 16215 2650 16224
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 296 13524 348 13530
rect 296 13466 348 13472
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10266 1624 11086
rect 1688 11014 1716 12174
rect 1872 11694 1900 13398
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1964 12782 1992 13126
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 2056 12442 2084 12582
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 9042 1624 9454
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 8090 1532 8298
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 204 3052 256 3058
rect 204 2994 256 3000
rect 216 480 244 2994
rect 1596 2990 1624 8502
rect 1688 5166 1716 10950
rect 1780 7993 1808 11494
rect 1872 11354 1900 11494
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 2148 11150 2176 12786
rect 2608 12442 2636 16215
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 2792 13870 2820 14486
rect 2884 14074 2912 16520
rect 3330 15872 3386 15881
rect 3330 15807 3386 15816
rect 3146 14648 3202 14657
rect 3146 14583 3202 14592
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 3068 13870 3096 14214
rect 2780 13864 2832 13870
rect 2686 13832 2742 13841
rect 2780 13806 2832 13812
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 2686 13767 2742 13776
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2516 11762 2544 12106
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2516 10606 2544 11698
rect 2700 11694 2728 13767
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2976 12714 3004 13262
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2792 11830 2820 12582
rect 2976 12238 3004 12650
rect 3160 12345 3188 14583
rect 3146 12336 3202 12345
rect 3146 12271 3202 12280
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2792 11354 2820 11494
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2424 9518 2452 10542
rect 2516 10062 2544 10542
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2056 8022 2084 8570
rect 2044 8016 2096 8022
rect 1766 7984 1822 7993
rect 2044 7958 2096 7964
rect 1766 7919 1822 7928
rect 2148 7886 2176 9046
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2148 7410 2176 7822
rect 2240 7546 2268 8230
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2608 7342 2636 7686
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2792 6769 2820 10406
rect 2884 8401 2912 12038
rect 2962 11384 3018 11393
rect 2962 11319 2964 11328
rect 3016 11319 3018 11328
rect 2964 11290 3016 11296
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 3068 10266 3096 10406
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2964 10056 3016 10062
rect 2962 10024 2964 10033
rect 3016 10024 3018 10033
rect 2962 9959 3018 9968
rect 2976 9761 3004 9959
rect 2962 9752 3018 9761
rect 3068 9722 3096 10066
rect 2962 9687 3018 9696
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2976 9178 3004 9386
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2976 8498 3004 9114
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2870 8392 2926 8401
rect 2870 8327 2926 8336
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2976 6848 3004 8298
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 3068 7342 3096 8230
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3160 6934 3188 12271
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 2884 6820 3004 6848
rect 2778 6760 2834 6769
rect 2412 6724 2464 6730
rect 2778 6695 2834 6704
rect 2412 6666 2464 6672
rect 2424 6322 2452 6666
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1872 5953 1900 6054
rect 1858 5944 1914 5953
rect 1858 5879 1914 5888
rect 2608 5817 2636 6122
rect 2594 5808 2650 5817
rect 2594 5743 2650 5752
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 2410 5672 2466 5681
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1780 3058 1808 5646
rect 2410 5607 2466 5616
rect 1858 5536 1914 5545
rect 1858 5471 1914 5480
rect 1872 5370 1900 5471
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1858 5128 1914 5137
rect 1858 5063 1914 5072
rect 1872 4826 1900 5063
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 2424 4690 2452 5607
rect 2884 5234 2912 6820
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2792 4729 2820 4762
rect 2778 4720 2834 4729
rect 2412 4684 2464 4690
rect 2778 4655 2834 4664
rect 2412 4626 2464 4632
rect 1858 4312 1914 4321
rect 1858 4247 1860 4256
rect 1912 4247 1914 4256
rect 1860 4218 1912 4224
rect 2134 4040 2190 4049
rect 2134 3975 2136 3984
rect 2188 3975 2190 3984
rect 2136 3946 2188 3952
rect 2780 3936 2832 3942
rect 2778 3904 2780 3913
rect 2832 3904 2834 3913
rect 2778 3839 2834 3848
rect 1858 3496 1914 3505
rect 1858 3431 1860 3440
rect 1912 3431 1914 3440
rect 1860 3402 1912 3408
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1584 2984 1636 2990
rect 2884 2938 2912 5034
rect 1584 2926 1636 2932
rect 664 2916 716 2922
rect 664 2858 716 2864
rect 2136 2916 2188 2922
rect 2136 2858 2188 2864
rect 2700 2910 2912 2938
rect 676 480 704 2858
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1124 2440 1176 2446
rect 1124 2382 1176 2388
rect 1136 480 1164 2382
rect 1688 480 1716 2790
rect 2148 480 2176 2858
rect 2700 480 2728 2910
rect 2778 2680 2834 2689
rect 2778 2615 2780 2624
rect 2832 2615 2834 2624
rect 2780 2586 2832 2592
rect 2976 1873 3004 6598
rect 3068 6225 3096 6734
rect 3252 6338 3280 11290
rect 3344 11234 3372 15807
rect 3528 13734 3556 16520
rect 3712 15298 3740 16623
rect 4158 16520 4214 17000
rect 4802 16520 4858 17000
rect 5446 16520 5502 17000
rect 6090 16520 6146 17000
rect 6734 16520 6790 17000
rect 7378 16520 7434 17000
rect 8022 16520 8078 17000
rect 8666 16520 8722 17000
rect 9310 16520 9366 17000
rect 9954 16520 10010 17000
rect 10598 16520 10654 17000
rect 11242 16520 11298 17000
rect 11886 16520 11942 17000
rect 12346 16688 12402 16697
rect 12346 16623 12402 16632
rect 4066 15464 4122 15473
rect 4066 15399 4122 15408
rect 3700 15292 3752 15298
rect 3700 15234 3752 15240
rect 4080 15230 4108 15399
rect 4068 15224 4120 15230
rect 4068 15166 4120 15172
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 4080 14346 4108 14991
rect 4068 14340 4120 14346
rect 4172 14328 4200 16520
rect 4172 14300 4292 14328
rect 4068 14282 4120 14288
rect 3698 14240 3754 14249
rect 3698 14175 3754 14184
rect 3712 14074 3740 14175
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 4264 13530 4292 14300
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 3698 13424 3754 13433
rect 4816 13394 4844 16520
rect 5460 13462 5488 16520
rect 6000 15292 6052 15298
rect 6000 15234 6052 15240
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 3698 13359 3754 13368
rect 4804 13388 4856 13394
rect 3712 13190 3740 13359
rect 4804 13330 4856 13336
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3422 13016 3478 13025
rect 3921 13008 4217 13028
rect 3422 12951 3478 12960
rect 4436 12980 4488 12986
rect 3436 11354 3464 12951
rect 4436 12922 4488 12928
rect 3792 12640 3844 12646
rect 3606 12608 3662 12617
rect 3792 12582 3844 12588
rect 3606 12543 3662 12552
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3344 11206 3464 11234
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3344 10538 3372 11086
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3344 10062 3372 10474
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3344 9586 3372 9998
rect 3436 9625 3464 11206
rect 3422 9616 3478 9625
rect 3332 9580 3384 9586
rect 3422 9551 3478 9560
rect 3332 9522 3384 9528
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3344 7886 3372 8434
rect 3436 8430 3464 9551
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3422 7848 3478 7857
rect 3422 7783 3478 7792
rect 3436 7342 3464 7783
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3252 6310 3372 6338
rect 3054 6216 3110 6225
rect 3054 6151 3110 6160
rect 3068 4010 3096 6151
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3252 4758 3280 5170
rect 3344 5166 3372 6310
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2962 1864 3018 1873
rect 2962 1799 3018 1808
rect 202 0 258 480
rect 662 0 718 480
rect 1122 0 1178 480
rect 1674 0 1730 480
rect 2134 0 2190 480
rect 2686 0 2742 480
rect 3068 241 3096 3470
rect 3148 2916 3200 2922
rect 3148 2858 3200 2864
rect 3160 480 3188 2858
rect 3252 649 3280 4422
rect 3344 4282 3372 5102
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3344 3097 3372 3878
rect 3330 3088 3386 3097
rect 3330 3023 3386 3032
rect 3436 2394 3464 7142
rect 3528 2582 3556 11290
rect 3620 9081 3648 12543
rect 3804 11626 3832 12582
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 3792 11620 3844 11626
rect 3792 11562 3844 11568
rect 4448 11354 4476 12922
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4540 11898 4568 12174
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 3698 10976 3754 10985
rect 3698 10911 3754 10920
rect 3712 10266 3740 10911
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4540 10742 4568 11834
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4528 10736 4580 10742
rect 4528 10678 4580 10684
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 4066 10160 4122 10169
rect 3606 9072 3662 9081
rect 3606 9007 3662 9016
rect 3606 8528 3662 8537
rect 3606 8463 3662 8472
rect 3620 8430 3648 8463
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3608 8016 3660 8022
rect 3606 7984 3608 7993
rect 3660 7984 3662 7993
rect 3606 7919 3662 7928
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3620 6361 3648 7142
rect 3804 6984 3832 10134
rect 4122 10130 4200 10146
rect 4122 10124 4212 10130
rect 4122 10118 4160 10124
rect 4066 10095 4122 10104
rect 4160 10066 4212 10072
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 4264 9704 4292 10678
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4080 9676 4292 9704
rect 4080 9518 4108 9676
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4080 8974 4108 9454
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4068 8968 4120 8974
rect 4172 8945 4200 9386
rect 4344 9036 4396 9042
rect 4264 8996 4344 9024
rect 4068 8910 4120 8916
rect 4158 8936 4214 8945
rect 4158 8871 4214 8880
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 4264 8498 4292 8996
rect 4344 8978 4396 8984
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4264 7546 4292 8298
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4356 7426 4384 8502
rect 4080 7398 4384 7426
rect 4080 7177 4108 7398
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 4172 7002 4200 7210
rect 3712 6956 3832 6984
rect 4160 6996 4212 7002
rect 3606 6352 3662 6361
rect 3606 6287 3662 6296
rect 3712 4978 3740 6956
rect 4160 6938 4212 6944
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3804 6458 3832 6802
rect 3884 6792 3936 6798
rect 3882 6760 3884 6769
rect 3936 6760 3938 6769
rect 3882 6695 3938 6704
rect 4252 6656 4304 6662
rect 4448 6610 4476 9930
rect 4252 6598 4304 6604
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3804 5710 3832 6394
rect 4264 6254 4292 6598
rect 4356 6582 4476 6610
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3620 4950 3740 4978
rect 3516 2576 3568 2582
rect 3516 2518 3568 2524
rect 3344 2366 3464 2394
rect 3344 1057 3372 2366
rect 3424 2304 3476 2310
rect 3422 2272 3424 2281
rect 3516 2304 3568 2310
rect 3476 2272 3478 2281
rect 3516 2246 3568 2252
rect 3422 2207 3478 2216
rect 3528 1465 3556 2246
rect 3514 1456 3570 1465
rect 3514 1391 3570 1400
rect 3330 1048 3386 1057
rect 3330 983 3386 992
rect 3238 640 3294 649
rect 3238 575 3294 584
rect 3620 480 3648 4950
rect 3804 3942 3832 5510
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4264 5166 4292 6190
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3790 3632 3846 3641
rect 3896 3602 3924 3946
rect 4264 3670 4292 5102
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 3790 3567 3846 3576
rect 3884 3596 3936 3602
rect 3804 2990 3832 3567
rect 3884 3538 3936 3544
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 4356 1306 4384 6582
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4448 5914 4476 6258
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4448 5370 4476 5714
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4146 4476 4422
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4448 2378 4476 3606
rect 4540 3058 4568 10406
rect 4632 7818 4660 12582
rect 4724 9489 4752 13126
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4908 11898 4936 12242
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4908 11150 4936 11834
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4802 10568 4858 10577
rect 4802 10503 4858 10512
rect 4710 9480 4766 9489
rect 4710 9415 4766 9424
rect 4724 8430 4752 9415
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4724 7546 4752 8230
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4724 7002 4752 7142
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4618 5808 4674 5817
rect 4618 5743 4674 5752
rect 4632 5710 4660 5743
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4724 5234 4752 6190
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4724 4214 4752 5170
rect 4816 4826 4844 10503
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4908 9722 4936 10202
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 4908 7410 4936 9658
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 5000 7188 5028 12718
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 11762 5580 12582
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5644 11937 5672 12378
rect 5630 11928 5686 11937
rect 5630 11863 5686 11872
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5354 11656 5410 11665
rect 5354 11591 5410 11600
rect 5368 11286 5396 11591
rect 5736 11558 5764 14010
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5368 10606 5396 10950
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5092 10266 5120 10406
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5170 10024 5226 10033
rect 5170 9959 5226 9968
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5092 7732 5120 9318
rect 5184 8838 5212 9959
rect 5276 9382 5304 10474
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 9994 5396 10406
rect 5460 10266 5488 11494
rect 5828 11234 5856 13806
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5736 11206 5856 11234
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5460 9722 5488 9998
rect 5552 9994 5580 10678
rect 5644 10577 5672 11154
rect 5630 10568 5686 10577
rect 5630 10503 5686 10512
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5184 7886 5212 8434
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5092 7704 5212 7732
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 4908 7160 5028 7188
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 4172 1278 4384 1306
rect 4172 480 4200 1278
rect 4632 480 4660 3538
rect 4724 2854 4752 4014
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4816 2514 4844 4014
rect 4908 3738 4936 7160
rect 5092 7002 5120 7346
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5000 4434 5028 6938
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5092 4622 5120 5034
rect 5184 4690 5212 7704
rect 5276 6458 5304 9318
rect 5368 8634 5396 9454
rect 5446 8936 5502 8945
rect 5446 8871 5502 8880
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5460 8242 5488 8871
rect 5552 8401 5580 9930
rect 5538 8392 5594 8401
rect 5538 8327 5594 8336
rect 5368 8214 5488 8242
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5368 4826 5396 8214
rect 5552 8090 5580 8230
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5460 7834 5488 7890
rect 5460 7806 5580 7834
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 6662 5488 7686
rect 5552 7546 5580 7806
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5644 5914 5672 10134
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4826 5672 4966
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5000 4406 5120 4434
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 5000 2446 5028 4218
rect 5092 3670 5120 4406
rect 5460 4214 5488 4490
rect 5448 4208 5500 4214
rect 5354 4176 5410 4185
rect 5448 4150 5500 4156
rect 5354 4111 5410 4120
rect 5368 4078 5396 4111
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 5276 3482 5304 3878
rect 5460 3738 5488 4150
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5276 3454 5396 3482
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5184 480 5212 3334
rect 5368 2990 5396 3454
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5736 2530 5764 11206
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5828 10266 5856 11086
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5828 9110 5856 10066
rect 5920 9466 5948 13942
rect 6012 13682 6040 15234
rect 6104 13870 6132 16520
rect 6748 14074 6776 16520
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 7392 13802 7420 16520
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 6012 13654 6132 13682
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6012 11801 6040 12582
rect 5998 11792 6054 11801
rect 5998 11727 6054 11736
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 6012 11234 6040 11494
rect 6104 11354 6132 13654
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6656 12374 6684 12786
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 6184 12368 6236 12374
rect 6644 12368 6696 12374
rect 6184 12310 6236 12316
rect 6472 12316 6644 12322
rect 6472 12310 6696 12316
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6012 11206 6132 11234
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6012 10062 6040 11086
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6104 10010 6132 11206
rect 6196 10470 6224 12310
rect 6472 12294 6684 12310
rect 6472 12102 6500 12294
rect 6656 12245 6684 12294
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6380 11558 6408 11630
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6104 9982 6224 10010
rect 5920 9438 6132 9466
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 9178 5948 9318
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5920 8362 5948 8978
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5828 6866 5856 7278
rect 5920 6934 5948 8298
rect 6012 7954 6040 8434
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6012 7002 6040 7890
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5920 5846 5948 6598
rect 6012 6118 6040 6598
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5908 5840 5960 5846
rect 6012 5817 6040 6054
rect 5908 5782 5960 5788
rect 5998 5808 6054 5817
rect 5998 5743 6054 5752
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4758 6040 4966
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 6012 4282 6040 4694
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6104 4060 6132 9438
rect 6196 9382 6224 9982
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6196 7585 6224 7958
rect 6182 7576 6238 7585
rect 6182 7511 6238 7520
rect 6288 7018 6316 11222
rect 6380 10266 6408 11290
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 9586 6408 9998
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6366 9344 6422 9353
rect 6366 9279 6422 9288
rect 6380 9178 6408 9279
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6380 8362 6408 9114
rect 6472 8974 6500 12038
rect 6748 11762 6776 12038
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6748 11626 6776 11698
rect 6932 11694 6960 12310
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6380 7410 6408 7890
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6288 6990 6408 7018
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6288 6458 6316 6802
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5710 6224 6054
rect 6288 5914 6316 6190
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6196 5166 6224 5646
rect 6288 5302 6316 5850
rect 6380 5302 6408 6990
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6196 4604 6224 5102
rect 6276 4616 6328 4622
rect 6196 4576 6276 4604
rect 6196 4128 6224 4576
rect 6276 4558 6328 4564
rect 6276 4140 6328 4146
rect 6196 4100 6276 4128
rect 6276 4082 6328 4088
rect 6104 4032 6215 4060
rect 6187 4026 6215 4032
rect 6187 3998 6224 4026
rect 5644 2502 5764 2530
rect 5644 480 5672 2502
rect 6196 480 6224 3998
rect 6288 3738 6316 4082
rect 6472 3942 6500 8774
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6472 3126 6500 3538
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 6564 626 6592 11018
rect 6656 10742 6684 11154
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 7300 10606 7328 12582
rect 7484 12374 7512 13194
rect 8036 12782 8064 16520
rect 8116 15224 8168 15230
rect 8116 15166 8168 15172
rect 8128 13433 8156 15166
rect 8114 13424 8170 13433
rect 8114 13359 8170 13368
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 7472 12368 7524 12374
rect 7852 12322 7880 12718
rect 7472 12310 7524 12316
rect 7760 12294 7880 12322
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7472 11688 7524 11694
rect 7564 11688 7616 11694
rect 7472 11630 7524 11636
rect 7562 11656 7564 11665
rect 7616 11656 7618 11665
rect 7484 11150 7512 11630
rect 7562 11591 7618 11600
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7484 10554 7512 11086
rect 7668 10674 7696 12038
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 6748 10266 6776 10542
rect 7484 10526 7604 10554
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 9058 6684 9318
rect 6748 9178 6776 9386
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 7300 9178 7328 9930
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 6656 9030 6776 9058
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6656 7478 6684 8910
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6748 6769 6776 9030
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7208 7546 7236 7890
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 6734 6760 6790 6769
rect 6734 6695 6790 6704
rect 7300 6118 7328 8366
rect 7392 8090 7420 8366
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 6748 5914 6776 6054
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 7300 5914 7328 6054
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7392 5846 7420 6122
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7392 5166 7420 5782
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 6748 2990 6776 5102
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 7300 3738 7328 3946
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6748 2378 6776 2926
rect 7208 2836 7236 3470
rect 7300 2990 7328 3674
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7208 2808 7328 2836
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 7196 2508 7248 2514
rect 7300 2496 7328 2808
rect 7392 2514 7420 3606
rect 7248 2468 7328 2496
rect 7380 2508 7432 2514
rect 7196 2450 7248 2456
rect 7380 2450 7432 2456
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 7484 1442 7512 10406
rect 7576 10130 7604 10526
rect 7668 10130 7696 10610
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7576 9450 7604 10066
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7562 9072 7618 9081
rect 7562 9007 7618 9016
rect 7576 8294 7604 9007
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 3058 7604 7686
rect 7668 6882 7696 8298
rect 7760 7256 7788 12294
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7852 8498 7880 11766
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7760 7228 7880 7256
rect 7668 6854 7788 6882
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6322 7696 6734
rect 7760 6458 7788 6854
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7668 3670 7696 5510
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7760 4690 7788 5102
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7852 4078 7880 7228
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7576 2446 7604 2858
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7116 1414 7512 1442
rect 6564 598 6684 626
rect 6656 480 6684 598
rect 7116 480 7144 1414
rect 7668 480 7696 3130
rect 7760 2854 7788 3402
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7944 2446 7972 10542
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8036 7546 8064 8434
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8036 7410 8064 7482
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8128 7002 8156 13359
rect 8680 12782 8708 16520
rect 9324 13802 9352 16520
rect 9968 14498 9996 16520
rect 10612 14498 10640 16520
rect 9968 14470 10548 14498
rect 10612 14470 11008 14498
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8576 12708 8628 12714
rect 8576 12650 8628 12656
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11286 8248 11494
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8300 10192 8352 10198
rect 8298 10160 8300 10169
rect 8352 10160 8354 10169
rect 8298 10095 8354 10104
rect 8404 10044 8432 12038
rect 8312 10016 8432 10044
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8220 7478 8248 8978
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8220 7206 8248 7414
rect 8312 7342 8340 10016
rect 8390 9888 8446 9897
rect 8390 9823 8446 9832
rect 8404 7857 8432 9823
rect 8482 9752 8538 9761
rect 8482 9687 8538 9696
rect 8496 9382 8524 9687
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8496 8276 8524 9318
rect 8588 8430 8616 12650
rect 8772 12306 8800 12650
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8496 8248 8616 8276
rect 8482 7984 8538 7993
rect 8482 7919 8484 7928
rect 8536 7919 8538 7928
rect 8484 7890 8536 7896
rect 8390 7848 8446 7857
rect 8390 7783 8446 7792
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8496 7274 8524 7754
rect 8588 7274 8616 8248
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8390 6896 8446 6905
rect 8024 6860 8076 6866
rect 8390 6831 8446 6840
rect 8024 6802 8076 6808
rect 8036 5681 8064 6802
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8022 5672 8078 5681
rect 8022 5607 8078 5616
rect 8128 3641 8156 6666
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8312 5370 8340 6394
rect 8404 6118 8432 6831
rect 8484 6656 8536 6662
rect 8588 6633 8616 7210
rect 8484 6598 8536 6604
rect 8574 6624 8630 6633
rect 8496 6322 8524 6598
rect 8574 6559 8630 6568
rect 8588 6322 8616 6559
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8404 5658 8432 6054
rect 8404 5642 8524 5658
rect 8404 5636 8536 5642
rect 8404 5630 8484 5636
rect 8484 5578 8536 5584
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 8114 3632 8170 3641
rect 8404 3602 8432 4150
rect 8496 3942 8524 4626
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8114 3567 8170 3576
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7944 2038 7972 2382
rect 7932 2032 7984 2038
rect 7932 1974 7984 1980
rect 8128 480 8156 2586
rect 8404 2446 8432 3538
rect 8496 2514 8524 3878
rect 8680 3738 8708 12242
rect 8772 11257 8800 12242
rect 9128 12232 9180 12238
rect 8942 12200 8998 12209
rect 9128 12174 9180 12180
rect 8942 12135 8998 12144
rect 8758 11248 8814 11257
rect 8758 11183 8814 11192
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8772 6254 8800 11086
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8864 10742 8892 10950
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8864 10441 8892 10678
rect 8850 10432 8906 10441
rect 8850 10367 8906 10376
rect 8956 10198 8984 12135
rect 9140 11762 9168 12174
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9140 11665 9168 11698
rect 9126 11656 9182 11665
rect 9126 11591 9182 11600
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8944 10192 8996 10198
rect 8864 10140 8944 10146
rect 8864 10134 8996 10140
rect 8864 10118 8984 10134
rect 8864 6905 8892 10118
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8956 9586 8984 9862
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8956 8974 8984 9522
rect 9048 9178 9076 11494
rect 9140 9654 9168 11494
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8850 6896 8906 6905
rect 8850 6831 8906 6840
rect 8956 6798 8984 8910
rect 9048 8265 9076 8978
rect 9034 8256 9090 8265
rect 9034 8191 9090 8200
rect 9140 7818 9168 8978
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9232 7426 9260 13738
rect 9416 10062 9444 13874
rect 10232 13796 10284 13802
rect 10232 13738 10284 13744
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9600 12238 9628 12378
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9586 11928 9642 11937
rect 9586 11863 9588 11872
rect 9640 11863 9642 11872
rect 9588 11834 9640 11840
rect 9586 11792 9642 11801
rect 9586 11727 9642 11736
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9324 8945 9352 9318
rect 9310 8936 9366 8945
rect 9310 8871 9366 8880
rect 9324 8566 9352 8871
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9416 8430 9444 9386
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9048 7398 9260 7426
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8864 4826 8892 6734
rect 9048 5710 9076 7398
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9232 6322 9260 7278
rect 9508 6934 9536 10406
rect 9600 8401 9628 11727
rect 9678 11112 9734 11121
rect 9678 11047 9734 11056
rect 9692 9994 9720 11047
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9692 8974 9720 9590
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9678 8800 9734 8809
rect 9678 8735 9734 8744
rect 9692 8498 9720 8735
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9586 8392 9642 8401
rect 9586 8327 9642 8336
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9600 7546 9628 7890
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9692 7342 9720 7822
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9140 5846 9168 6122
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 9232 5710 9260 6258
rect 9310 6216 9366 6225
rect 9310 6151 9366 6160
rect 9324 5914 9352 6151
rect 9508 5930 9536 6870
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9416 5902 9536 5930
rect 9036 5704 9088 5710
rect 8956 5664 9036 5692
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8864 4690 8892 4762
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8956 4554 8984 5664
rect 9036 5646 9088 5652
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9048 4826 9076 5034
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8944 4548 8996 4554
rect 8944 4490 8996 4496
rect 8956 4214 8984 4490
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8668 2984 8720 2990
rect 8956 2972 8984 3606
rect 9048 3602 9076 4762
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8720 2944 8984 2972
rect 8668 2926 8720 2932
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8680 480 8708 2790
rect 9140 480 9168 5510
rect 9218 4856 9274 4865
rect 9218 4791 9274 4800
rect 9232 3670 9260 4791
rect 9324 4185 9352 5578
rect 9416 5030 9444 5902
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9508 5370 9536 5714
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 5370 9628 5646
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9310 4176 9366 4185
rect 9310 4111 9366 4120
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9600 3602 9628 4422
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9692 480 9720 6598
rect 9784 3058 9812 13262
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 10138 10704 10194 10713
rect 10138 10639 10194 10648
rect 10152 10470 10180 10639
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 10140 9376 10192 9382
rect 10138 9344 10140 9353
rect 10192 9344 10194 9353
rect 10138 9279 10194 9288
rect 10046 9072 10102 9081
rect 10046 9007 10102 9016
rect 10060 8906 10088 9007
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 10060 7857 10088 8502
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10152 8090 10180 8298
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10046 7848 10102 7857
rect 10046 7783 10102 7792
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9876 4622 9904 5102
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9954 3496 10010 3505
rect 10060 3466 10088 4014
rect 9954 3431 9956 3440
rect 10008 3431 10010 3440
rect 10048 3460 10100 3466
rect 9956 3402 10008 3408
rect 10048 3402 10100 3408
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9784 2378 9812 2858
rect 10244 2582 10272 13738
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10336 10606 10364 11086
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10428 10674 10456 10950
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10062 10364 10406
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 6254 10364 9998
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10428 6730 10456 9318
rect 10520 7426 10548 14470
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10704 10198 10732 10406
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10612 7562 10640 9658
rect 10704 9042 10732 9862
rect 10796 9042 10824 10542
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10796 8945 10824 8978
rect 10782 8936 10838 8945
rect 10782 8871 10838 8880
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10704 7750 10732 8366
rect 10796 7857 10824 8774
rect 10782 7848 10838 7857
rect 10782 7783 10838 7792
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10612 7534 10824 7562
rect 10520 7398 10640 7426
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10520 6497 10548 6802
rect 10506 6488 10562 6497
rect 10506 6423 10562 6432
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10520 5658 10548 6423
rect 10336 5630 10548 5658
rect 10336 4214 10364 5630
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10428 5098 10456 5510
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10428 4010 10456 5034
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 9772 2372 9824 2378
rect 9772 2314 9824 2320
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 10336 1442 10364 3538
rect 10428 3398 10456 3538
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10520 2922 10548 4558
rect 10612 3670 10640 7398
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 6361 10732 6734
rect 10690 6352 10746 6361
rect 10690 6287 10746 6296
rect 10796 5930 10824 7534
rect 10704 5902 10824 5930
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 10508 2916 10560 2922
rect 10508 2858 10560 2864
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 10428 2038 10456 2518
rect 10520 2310 10548 2858
rect 10704 2854 10732 5902
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10796 4690 10824 4966
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10796 4010 10824 4626
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 10796 2922 10824 3606
rect 10888 3058 10916 12718
rect 10980 9722 11008 14470
rect 11150 13832 11206 13841
rect 11256 13802 11284 16520
rect 11150 13767 11206 13776
rect 11244 13796 11296 13802
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11072 11898 11100 12378
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 11072 10606 11100 11834
rect 11164 10674 11192 13767
rect 11244 13738 11296 13744
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11058 10432 11114 10441
rect 11058 10367 11114 10376
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 11072 9466 11100 10367
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10980 9438 11100 9466
rect 10980 9058 11008 9438
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11072 9178 11100 9318
rect 11164 9178 11192 9522
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 10980 9030 11192 9058
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10980 6798 11008 8842
rect 11058 8800 11114 8809
rect 11058 8735 11114 8744
rect 11072 8022 11100 8735
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11072 7342 11100 7822
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10980 5914 11008 6326
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10980 5166 11008 5646
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10980 4078 11008 5102
rect 11164 5098 11192 9030
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11072 4282 11100 4762
rect 11152 4752 11204 4758
rect 11150 4720 11152 4729
rect 11204 4720 11206 4729
rect 11150 4655 11206 4664
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10980 3602 11008 3878
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11072 3097 11100 3470
rect 11152 3120 11204 3126
rect 11058 3088 11114 3097
rect 10876 3052 10928 3058
rect 11152 3062 11204 3068
rect 11058 3023 11114 3032
rect 10876 2994 10928 3000
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10416 2032 10468 2038
rect 10416 1974 10468 1980
rect 10152 1414 10364 1442
rect 10152 480 10180 1414
rect 10612 480 10640 2790
rect 11164 480 11192 3062
rect 11256 3058 11284 12310
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11348 10674 11376 11154
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11348 9654 11376 10066
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11348 7886 11376 9114
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11440 6066 11468 12786
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11532 9382 11560 9590
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11532 8498 11560 9046
rect 11624 9042 11652 11834
rect 11716 9654 11744 12242
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11808 10470 11836 10950
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11808 10062 11836 10406
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11704 9648 11756 9654
rect 11900 9602 11928 16520
rect 12164 15224 12216 15230
rect 12164 15166 12216 15172
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11704 9590 11756 9596
rect 11808 9574 11928 9602
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11716 9110 11744 9318
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11624 8566 11652 8978
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11532 6866 11560 8026
rect 11624 7886 11652 8230
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11532 6254 11560 6598
rect 11624 6322 11652 7686
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11348 6038 11468 6066
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11348 2582 11376 6038
rect 11716 5370 11744 9046
rect 11808 7834 11836 9574
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11900 8090 11928 9454
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11808 7806 11928 7834
rect 11900 6322 11928 7806
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11808 5914 11836 6258
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11704 5092 11756 5098
rect 11704 5034 11756 5040
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11440 3126 11468 3606
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11624 480 11652 3470
rect 11716 3398 11744 5034
rect 11992 4758 12020 13738
rect 12176 12306 12204 15166
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12084 9602 12112 12174
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 11529 12204 11630
rect 12162 11520 12218 11529
rect 12162 11455 12218 11464
rect 12268 11336 12296 14350
rect 12360 12170 12388 16623
rect 12530 16520 12586 17000
rect 13174 16520 13230 17000
rect 13818 16520 13874 17000
rect 14462 16520 14518 17000
rect 15106 16520 15162 17000
rect 15750 16520 15806 17000
rect 16394 16520 16450 17000
rect 17038 16520 17094 17000
rect 17682 16520 17738 17000
rect 18326 16520 18382 17000
rect 18970 16520 19026 17000
rect 19614 16520 19670 17000
rect 12544 13682 12572 16520
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12452 13654 12572 13682
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12176 11308 12296 11336
rect 12176 10044 12204 11308
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12268 10713 12296 10746
rect 12254 10704 12310 10713
rect 12254 10639 12310 10648
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12268 10169 12296 10542
rect 12360 10538 12388 11698
rect 12452 11665 12480 13654
rect 12728 13190 12756 14282
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 13188 13410 13216 16520
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13464 13705 13492 14214
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13450 13696 13506 13705
rect 13450 13631 13506 13640
rect 13556 13530 13584 14010
rect 13648 13530 13676 14486
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13188 13382 13584 13410
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12438 11656 12494 11665
rect 12438 11591 12494 11600
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12254 10160 12310 10169
rect 12254 10095 12310 10104
rect 12256 10056 12308 10062
rect 12176 10016 12256 10044
rect 12256 9998 12308 10004
rect 12084 9574 12296 9602
rect 12360 9586 12388 10474
rect 12452 10266 12480 11494
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 12084 8634 12112 9454
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12176 9353 12204 9386
rect 12162 9344 12218 9353
rect 12162 9279 12218 9288
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12072 8288 12124 8294
rect 12070 8256 12072 8265
rect 12124 8256 12126 8265
rect 12070 8191 12126 8200
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12084 7410 12112 7890
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12176 6458 12204 8774
rect 12268 8294 12296 9574
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12360 8430 12388 9386
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12360 7546 12388 7822
rect 12348 7540 12400 7546
rect 12268 7500 12348 7528
rect 12268 6798 12296 7500
rect 12348 7482 12400 7488
rect 12452 7290 12480 9998
rect 12360 7262 12480 7290
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12164 5840 12216 5846
rect 12162 5808 12164 5817
rect 12216 5808 12218 5817
rect 12268 5778 12296 6734
rect 12162 5743 12218 5752
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12070 4856 12126 4865
rect 12070 4791 12126 4800
rect 12084 4758 12112 4791
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11716 2514 11744 3334
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11808 1873 11836 4422
rect 12360 3670 12388 7262
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6866 12480 7142
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12438 6760 12494 6769
rect 12438 6695 12494 6704
rect 12452 4758 12480 6695
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12544 4010 12572 12038
rect 12636 10305 12664 12718
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12728 10996 12756 12242
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 12728 10968 12848 10996
rect 12820 10452 12848 10968
rect 12990 10840 13046 10849
rect 12990 10775 12992 10784
rect 13044 10775 13046 10784
rect 12992 10746 13044 10752
rect 13096 10674 13124 11222
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12728 10424 12848 10452
rect 12622 10296 12678 10305
rect 12622 10231 12678 10240
rect 12728 10248 12756 10424
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 12728 10220 12848 10248
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12714 10024 12770 10033
rect 12636 9722 12664 9998
rect 12714 9959 12770 9968
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12728 9568 12756 9959
rect 12636 9540 12756 9568
rect 12636 8265 12664 9540
rect 12820 9518 12848 10220
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 8634 12756 9318
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13082 9072 13138 9081
rect 13082 9007 13138 9016
rect 13096 8974 13124 9007
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12622 8256 12678 8265
rect 12622 8191 12678 8200
rect 12728 8106 12756 8366
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12636 8078 12756 8106
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12268 3482 12296 3538
rect 12176 3454 12296 3482
rect 12346 3496 12402 3505
rect 11794 1864 11850 1873
rect 11794 1799 11850 1808
rect 12176 480 12204 3454
rect 12636 3466 12664 8078
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 13096 7857 13124 7958
rect 13082 7848 13138 7857
rect 12900 7812 12952 7818
rect 13082 7783 13138 7792
rect 12900 7754 12952 7760
rect 12912 7410 12940 7754
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 7410 13124 7686
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13188 7342 13216 13126
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13280 8956 13308 12582
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 10266 13400 11494
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13372 9178 13400 9318
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13280 8928 13400 8956
rect 13266 8664 13322 8673
rect 13266 8599 13322 8608
rect 13176 7336 13228 7342
rect 12990 7304 13046 7313
rect 13176 7278 13228 7284
rect 12990 7239 12992 7248
rect 13044 7239 13046 7248
rect 12992 7210 13044 7216
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 13082 6896 13138 6905
rect 13188 6866 13216 7142
rect 13082 6831 13138 6840
rect 13176 6860 13228 6866
rect 13096 6798 13124 6831
rect 13176 6802 13228 6808
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12728 5166 12756 6394
rect 13176 6180 13228 6186
rect 13280 6168 13308 8599
rect 13228 6140 13308 6168
rect 13176 6122 13228 6128
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 13372 5098 13400 8928
rect 13360 5092 13412 5098
rect 13360 5034 13412 5040
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 12346 3431 12402 3440
rect 12624 3460 12676 3466
rect 12360 3194 12388 3431
rect 12624 3402 12676 3408
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12268 2961 12296 3130
rect 12254 2952 12310 2961
rect 12254 2887 12310 2896
rect 12636 2530 12664 3402
rect 12990 3224 13046 3233
rect 12990 3159 13046 3168
rect 13004 3058 13032 3159
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13096 2961 13124 2994
rect 13082 2952 13138 2961
rect 13082 2887 13084 2896
rect 13136 2887 13138 2896
rect 13084 2858 13136 2864
rect 13096 2827 13124 2858
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 12544 2502 12664 2530
rect 12544 2446 12572 2502
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12636 480 12664 2382
rect 13188 480 13216 4082
rect 13372 4049 13400 4082
rect 13358 4040 13414 4049
rect 13358 3975 13414 3984
rect 13464 2582 13492 12038
rect 13556 11801 13584 13382
rect 13648 13297 13676 13466
rect 13634 13288 13690 13297
rect 13634 13223 13690 13232
rect 13542 11792 13598 11801
rect 13542 11727 13598 11736
rect 13636 11756 13688 11762
rect 13740 11744 13768 14282
rect 13832 13705 13860 16520
rect 13910 14648 13966 14657
rect 13910 14583 13966 14592
rect 13818 13696 13874 13705
rect 13818 13631 13874 13640
rect 13924 12714 13952 14583
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14016 13734 14044 14214
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14372 13864 14424 13870
rect 14476 13852 14504 16520
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 14424 13824 14504 13852
rect 14924 13864 14976 13870
rect 14372 13806 14424 13812
rect 14924 13806 14976 13812
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13818 12336 13874 12345
rect 13818 12271 13874 12280
rect 13832 12238 13860 12271
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13740 11716 13860 11744
rect 13636 11698 13688 11704
rect 13648 11642 13676 11698
rect 13544 11620 13596 11626
rect 13648 11614 13768 11642
rect 13544 11562 13596 11568
rect 13556 11286 13584 11562
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13556 10470 13584 11086
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10062 13584 10406
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 8974 13584 9998
rect 13648 9654 13676 11494
rect 13740 11150 13768 11614
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13740 10010 13768 10746
rect 13832 10713 13860 11716
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13818 10704 13874 10713
rect 13818 10639 13874 10648
rect 13924 10266 13952 11086
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13740 9982 13860 10010
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 8498 13584 8910
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13556 7721 13584 8230
rect 13542 7712 13598 7721
rect 13542 7647 13598 7656
rect 13542 7440 13598 7449
rect 13542 7375 13598 7384
rect 13556 5522 13584 7375
rect 13648 7002 13676 9318
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13634 6896 13690 6905
rect 13634 6831 13690 6840
rect 13648 6390 13676 6831
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13740 5522 13768 9862
rect 13832 9586 13860 9982
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13832 9178 13860 9522
rect 13924 9353 13952 10202
rect 13910 9344 13966 9353
rect 13910 9279 13966 9288
rect 14016 9217 14044 12718
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14002 9208 14058 9217
rect 13820 9172 13872 9178
rect 13872 9132 13952 9160
rect 14002 9143 14058 9152
rect 13820 9114 13872 9120
rect 13818 9072 13874 9081
rect 13818 9007 13820 9016
rect 13872 9007 13874 9016
rect 13820 8978 13872 8984
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13832 6798 13860 8774
rect 13924 8498 13952 9132
rect 14108 9024 14136 11494
rect 14016 8996 14136 9024
rect 14016 8566 14044 8996
rect 14094 8936 14150 8945
rect 14094 8871 14150 8880
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13924 7546 13952 8434
rect 14016 7954 14044 8502
rect 14108 7993 14136 8871
rect 14094 7984 14150 7993
rect 14004 7948 14056 7954
rect 14094 7919 14150 7928
rect 14004 7890 14056 7896
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13910 7440 13966 7449
rect 13910 7375 13966 7384
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13556 5494 13676 5522
rect 13740 5494 13860 5522
rect 13544 5364 13596 5370
rect 13648 5352 13676 5494
rect 13832 5370 13860 5494
rect 13820 5364 13872 5370
rect 13648 5324 13768 5352
rect 13544 5306 13596 5312
rect 13556 3670 13584 5306
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13648 480 13676 5170
rect 13740 4185 13768 5324
rect 13820 5306 13872 5312
rect 13818 4856 13874 4865
rect 13818 4791 13874 4800
rect 13832 4758 13860 4791
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13818 4312 13874 4321
rect 13818 4247 13874 4256
rect 13726 4176 13782 4185
rect 13726 4111 13782 4120
rect 13726 4040 13782 4049
rect 13726 3975 13782 3984
rect 13740 3534 13768 3975
rect 13832 3602 13860 4247
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13924 1426 13952 7375
rect 14108 7002 14136 7919
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14016 6322 14044 6598
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14108 5778 14136 6190
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14200 5234 14228 13806
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14292 4554 14320 11494
rect 14384 11393 14412 12718
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14370 11384 14426 11393
rect 14370 11319 14426 11328
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14384 4622 14412 11154
rect 14476 10198 14504 11562
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14280 4548 14332 4554
rect 14280 4490 14332 4496
rect 14096 4004 14148 4010
rect 14096 3946 14148 3952
rect 13912 1420 13964 1426
rect 13912 1362 13964 1368
rect 14108 480 14136 3946
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14384 2922 14412 3402
rect 14372 2916 14424 2922
rect 14372 2858 14424 2864
rect 14278 2680 14334 2689
rect 14278 2615 14334 2624
rect 14292 2582 14320 2615
rect 14280 2576 14332 2582
rect 14280 2518 14332 2524
rect 3054 232 3110 241
rect 3054 167 3110 176
rect 3146 0 3202 480
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4618 0 4674 480
rect 5170 0 5226 480
rect 5630 0 5686 480
rect 6182 0 6238 480
rect 6642 0 6698 480
rect 7102 0 7158 480
rect 7654 0 7710 480
rect 8114 0 8170 480
rect 8666 0 8722 480
rect 9126 0 9182 480
rect 9678 0 9734 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 11150 0 11206 480
rect 11610 0 11666 480
rect 12162 0 12218 480
rect 12622 0 12678 480
rect 13174 0 13230 480
rect 13634 0 13690 480
rect 14094 0 14150 480
rect 14476 241 14504 8774
rect 14568 8401 14596 12582
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14660 11354 14688 11562
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14660 10713 14688 10950
rect 14646 10704 14702 10713
rect 14646 10639 14702 10648
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14554 8392 14610 8401
rect 14554 8327 14610 8336
rect 14660 6882 14688 10066
rect 14568 6854 14688 6882
rect 14568 4162 14596 6854
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14660 6186 14688 6734
rect 14752 6458 14780 12650
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14738 5672 14794 5681
rect 14738 5607 14794 5616
rect 14568 4134 14688 4162
rect 14554 4040 14610 4049
rect 14554 3975 14556 3984
rect 14608 3975 14610 3984
rect 14556 3946 14608 3952
rect 14660 3890 14688 4134
rect 14568 3862 14688 3890
rect 14568 3058 14596 3862
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14568 2038 14596 2790
rect 14556 2032 14608 2038
rect 14556 1974 14608 1980
rect 14660 480 14688 3674
rect 14752 3058 14780 5607
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14844 2922 14872 12038
rect 14936 4146 14964 13806
rect 15028 13258 15056 14418
rect 15120 13870 15148 16520
rect 15382 15056 15438 15065
rect 15382 14991 15438 15000
rect 15396 14346 15424 14991
rect 15764 14482 15792 16520
rect 15934 16280 15990 16289
rect 15934 16215 15990 16224
rect 15948 15230 15976 16215
rect 15936 15224 15988 15230
rect 15936 15166 15988 15172
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 16210 14240 16266 14249
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15212 13394 15240 14214
rect 15782 14172 16078 14192
rect 16210 14175 16266 14184
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15580 13462 15608 14010
rect 16224 13938 16252 14175
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15672 13705 15700 13806
rect 15658 13696 15714 13705
rect 15658 13631 15714 13640
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15028 13161 15056 13194
rect 15384 13184 15436 13190
rect 15014 13152 15070 13161
rect 15384 13126 15436 13132
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15014 13087 15070 13096
rect 15396 12918 15424 13126
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15028 8673 15056 12582
rect 15108 11688 15160 11694
rect 15212 11665 15240 12854
rect 15488 12730 15516 13126
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15304 12702 15516 12730
rect 15108 11630 15160 11636
rect 15198 11656 15254 11665
rect 15120 11558 15148 11630
rect 15198 11591 15254 11600
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15212 11218 15240 11290
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15106 11112 15162 11121
rect 15304 11098 15332 12702
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15106 11047 15162 11056
rect 15212 11070 15332 11098
rect 15120 11014 15148 11047
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 15120 10033 15148 10134
rect 15106 10024 15162 10033
rect 15106 9959 15162 9968
rect 15014 8664 15070 8673
rect 15014 8599 15070 8608
rect 15120 8514 15148 9959
rect 15028 8486 15148 8514
rect 15028 7954 15056 8486
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15028 7206 15056 7890
rect 15120 7546 15148 8298
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15120 6730 15148 7482
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 15212 6440 15240 11070
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15304 8809 15332 10134
rect 15396 9330 15424 12242
rect 15566 12200 15622 12209
rect 15566 12135 15622 12144
rect 15580 11354 15608 12135
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15948 11257 15976 11698
rect 15934 11248 15990 11257
rect 15934 11183 15990 11192
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15476 10532 15528 10538
rect 15580 10520 15608 11018
rect 15528 10492 15608 10520
rect 15476 10474 15528 10480
rect 15580 9738 15608 10492
rect 15672 10266 15700 11086
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 16040 10180 16068 10542
rect 16132 10305 16160 12038
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16224 11558 16252 11766
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16118 10296 16174 10305
rect 16118 10231 16174 10240
rect 16040 10152 16160 10180
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 15571 9722 15608 9738
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 16132 9625 16160 10152
rect 16118 9616 16174 9625
rect 16118 9551 16174 9560
rect 16132 9450 16160 9551
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 15396 9302 15608 9330
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15290 8800 15346 8809
rect 15290 8735 15346 8744
rect 15396 8294 15424 8978
rect 15384 8288 15436 8294
rect 15290 8256 15346 8265
rect 15384 8230 15436 8236
rect 15290 8191 15346 8200
rect 15304 8022 15332 8191
rect 15292 8016 15344 8022
rect 15292 7958 15344 7964
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15028 6412 15240 6440
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 15028 2582 15056 6412
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15212 5574 15240 6122
rect 15200 5568 15252 5574
rect 15106 5536 15162 5545
rect 15200 5510 15252 5516
rect 15106 5471 15162 5480
rect 15120 4758 15148 5471
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15212 3942 15240 5510
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15198 3632 15254 3641
rect 15198 3567 15254 3576
rect 15212 3398 15240 3567
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 15198 2680 15254 2689
rect 15198 2615 15200 2624
rect 15252 2615 15254 2624
rect 15200 2586 15252 2592
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15120 480 15148 2382
rect 15304 1465 15332 7686
rect 15396 5250 15424 8230
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15488 6905 15516 7958
rect 15474 6896 15530 6905
rect 15474 6831 15530 6840
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15488 5370 15516 6734
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15396 5222 15516 5250
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15396 3738 15424 4558
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15488 3602 15516 5222
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15396 3398 15424 3538
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15580 3058 15608 9302
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15672 8634 15700 9046
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 16224 8634 16252 11086
rect 16316 10962 16344 14418
rect 16408 13705 16436 16520
rect 16394 13696 16450 13705
rect 16394 13631 16450 13640
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16408 11150 16436 12582
rect 16500 12345 16528 13330
rect 17052 13326 17080 16520
rect 17696 14414 17724 16520
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 18340 13530 18368 16520
rect 18418 15872 18474 15881
rect 18418 15807 18474 15816
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 17866 13424 17922 13433
rect 17866 13359 17868 13368
rect 17920 13359 17922 13368
rect 17868 13330 17920 13336
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17960 12912 18012 12918
rect 17866 12880 17922 12889
rect 17960 12854 18012 12860
rect 17866 12815 17922 12824
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 16486 12336 16542 12345
rect 16486 12271 16542 12280
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16316 10934 16436 10962
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16316 8634 16344 9998
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 15672 7818 15700 8570
rect 15750 8528 15806 8537
rect 15750 8463 15806 8472
rect 15764 8430 15792 8463
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16302 8392 16358 8401
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15672 6458 15700 6938
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 16132 6390 16160 7210
rect 16120 6384 16172 6390
rect 15658 6352 15714 6361
rect 16120 6326 16172 6332
rect 15658 6287 15714 6296
rect 15672 5778 15700 6287
rect 16132 5846 16160 6326
rect 16120 5840 16172 5846
rect 16120 5782 16172 5788
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 15672 3097 15700 5510
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 16132 5166 16160 5510
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 15936 5024 15988 5030
rect 16224 5012 16252 8366
rect 16302 8327 16358 8336
rect 16316 5409 16344 8327
rect 16302 5400 16358 5409
rect 16302 5335 16358 5344
rect 16304 5296 16356 5302
rect 16304 5238 16356 5244
rect 15936 4966 15988 4972
rect 16132 4984 16252 5012
rect 15948 4826 15976 4966
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 15934 4176 15990 4185
rect 15934 4111 15936 4120
rect 15988 4111 15990 4120
rect 15936 4082 15988 4088
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15752 3936 15804 3942
rect 15948 3913 15976 3946
rect 15752 3878 15804 3884
rect 15934 3904 15990 3913
rect 15764 3534 15792 3878
rect 15934 3839 15990 3848
rect 15842 3768 15898 3777
rect 15842 3703 15844 3712
rect 15896 3703 15898 3712
rect 15844 3674 15896 3680
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 15658 3088 15714 3097
rect 15568 3052 15620 3058
rect 15658 3023 15714 3032
rect 15568 2994 15620 3000
rect 15934 2952 15990 2961
rect 15660 2916 15712 2922
rect 15934 2887 15936 2896
rect 15660 2858 15712 2864
rect 15988 2887 15990 2896
rect 15936 2858 15988 2864
rect 15290 1456 15346 1465
rect 15290 1391 15346 1400
rect 15672 480 15700 2858
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16132 480 16160 4984
rect 16316 2281 16344 5238
rect 16408 4758 16436 10934
rect 16500 10606 16528 11630
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16500 10062 16528 10406
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16500 9518 16528 9998
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16486 9072 16542 9081
rect 16486 9007 16542 9016
rect 16500 7290 16528 9007
rect 16592 7449 16620 11494
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16684 9518 16712 10474
rect 16776 9654 16804 11086
rect 16868 10266 16896 11154
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16854 10160 16910 10169
rect 16854 10095 16910 10104
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16684 9178 16712 9454
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16684 8498 16712 9114
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16578 7440 16634 7449
rect 16578 7375 16634 7384
rect 16500 7262 16620 7290
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16500 6322 16528 7142
rect 16592 7002 16620 7262
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16684 6730 16712 8298
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 8090 16804 8230
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16868 6934 16896 10095
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16500 5234 16528 6258
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16486 5128 16542 5137
rect 16486 5063 16542 5072
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16302 2272 16358 2281
rect 16302 2207 16358 2216
rect 16408 1057 16436 3334
rect 16500 2446 16528 5063
rect 16592 3738 16620 5646
rect 16684 5370 16712 6122
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16776 4690 16804 5850
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16776 3738 16804 4626
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16868 3058 16896 6258
rect 16960 4146 16988 12242
rect 17420 12186 17448 12582
rect 17420 12158 17724 12186
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 17052 10470 17080 11086
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 17144 10282 17172 11698
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17236 10305 17264 10542
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17052 10254 17172 10282
rect 17222 10296 17278 10305
rect 17052 6322 17080 10254
rect 17222 10231 17278 10240
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17144 9178 17172 10066
rect 17236 9586 17264 10066
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17222 9480 17278 9489
rect 17222 9415 17224 9424
rect 17276 9415 17278 9424
rect 17224 9386 17276 9392
rect 17222 9344 17278 9353
rect 17222 9279 17278 9288
rect 17236 9178 17264 9279
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17236 8004 17264 9114
rect 17144 7976 17264 8004
rect 17144 6390 17172 7976
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 17236 6798 17264 7754
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17328 6610 17356 10406
rect 17420 8265 17448 11494
rect 17406 8256 17462 8265
rect 17406 8191 17462 8200
rect 17512 7857 17540 12038
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17604 9110 17632 11834
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17604 8090 17632 8910
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17498 7848 17554 7857
rect 17498 7783 17554 7792
rect 17406 7032 17462 7041
rect 17406 6967 17462 6976
rect 17420 6866 17448 6967
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17236 6582 17356 6610
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 17052 5234 17080 5646
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17052 4690 17080 5170
rect 17144 4826 17172 6190
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17130 4720 17186 4729
rect 17040 4684 17092 4690
rect 17130 4655 17186 4664
rect 17040 4626 17092 4632
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17052 3194 17080 3538
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16672 1420 16724 1426
rect 16672 1362 16724 1368
rect 16394 1048 16450 1057
rect 16394 983 16450 992
rect 16684 480 16712 1362
rect 17144 480 17172 4655
rect 17236 649 17264 6582
rect 17696 6497 17724 12158
rect 17880 11762 17908 12815
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17866 11656 17922 11665
rect 17866 11591 17922 11600
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17788 9586 17816 9998
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17788 8974 17816 9522
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17682 6488 17738 6497
rect 17682 6423 17738 6432
rect 17788 6338 17816 8774
rect 17880 8022 17908 11591
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17604 6310 17816 6338
rect 17498 6216 17554 6225
rect 17498 6151 17554 6160
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17328 5914 17356 6054
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17314 5672 17370 5681
rect 17314 5607 17370 5616
rect 17328 5166 17356 5607
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17420 4865 17448 6054
rect 17512 5846 17540 6151
rect 17500 5840 17552 5846
rect 17500 5782 17552 5788
rect 17406 4856 17462 4865
rect 17406 4791 17462 4800
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17328 3670 17356 4558
rect 17316 3664 17368 3670
rect 17316 3606 17368 3612
rect 17222 640 17278 649
rect 17222 575 17278 584
rect 17604 480 17632 6310
rect 17880 6236 17908 7686
rect 17788 6208 17908 6236
rect 17682 5944 17738 5953
rect 17682 5879 17684 5888
rect 17736 5879 17738 5888
rect 17684 5850 17736 5856
rect 17682 4040 17738 4049
rect 17682 3975 17738 3984
rect 17696 2650 17724 3975
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17788 2514 17816 6208
rect 17972 4842 18000 12854
rect 18064 7041 18092 13126
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18050 7032 18106 7041
rect 18050 6967 18106 6976
rect 18156 5273 18184 11018
rect 18248 6089 18276 12038
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18234 6080 18290 6089
rect 18234 6015 18290 6024
rect 18340 5846 18368 11698
rect 18432 10266 18460 15807
rect 18694 13288 18750 13297
rect 18984 13258 19012 16520
rect 19628 13734 19656 16520
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 18694 13223 18750 13232
rect 18972 13252 19024 13258
rect 18510 10840 18566 10849
rect 18510 10775 18566 10784
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18524 9926 18552 10775
rect 18602 10568 18658 10577
rect 18602 10503 18658 10512
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 18142 5264 18198 5273
rect 18142 5199 18198 5208
rect 17972 4814 18184 4842
rect 17866 4448 17922 4457
rect 17866 4383 17922 4392
rect 17880 3738 17908 4383
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 18156 480 18184 4814
rect 18616 480 18644 10503
rect 18708 9761 18736 13223
rect 18972 13194 19024 13200
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 18694 9752 18750 9761
rect 18694 9687 18750 9696
rect 18972 5704 19024 5710
rect 18970 5672 18972 5681
rect 19024 5672 19026 5681
rect 18970 5607 19026 5616
rect 19168 480 19196 12106
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 19628 480 19656 11766
rect 14462 232 14518 241
rect 14462 167 14518 176
rect 14646 0 14702 480
rect 15106 0 15162 480
rect 15658 0 15714 480
rect 16118 0 16174 480
rect 16670 0 16726 480
rect 17130 0 17186 480
rect 17590 0 17646 480
rect 18142 0 18198 480
rect 18602 0 18658 480
rect 19154 0 19210 480
rect 19614 0 19670 480
<< via2 >>
rect 3698 16632 3754 16688
rect 2594 16224 2650 16280
rect 3330 15816 3386 15872
rect 3146 14592 3202 14648
rect 2686 13776 2742 13832
rect 3146 12280 3202 12336
rect 1766 7928 1822 7984
rect 2962 11348 3018 11384
rect 2962 11328 2964 11348
rect 2964 11328 3016 11348
rect 3016 11328 3018 11348
rect 2962 10004 2964 10024
rect 2964 10004 3016 10024
rect 3016 10004 3018 10024
rect 2962 9968 3018 10004
rect 2962 9696 3018 9752
rect 2870 8336 2926 8392
rect 2778 6704 2834 6760
rect 1858 5888 1914 5944
rect 2594 5752 2650 5808
rect 2410 5616 2466 5672
rect 1858 5480 1914 5536
rect 1858 5072 1914 5128
rect 2778 4664 2834 4720
rect 1858 4276 1914 4312
rect 1858 4256 1860 4276
rect 1860 4256 1912 4276
rect 1912 4256 1914 4276
rect 2134 4004 2190 4040
rect 2134 3984 2136 4004
rect 2136 3984 2188 4004
rect 2188 3984 2190 4004
rect 2778 3884 2780 3904
rect 2780 3884 2832 3904
rect 2832 3884 2834 3904
rect 2778 3848 2834 3884
rect 1858 3460 1914 3496
rect 1858 3440 1860 3460
rect 1860 3440 1912 3460
rect 1912 3440 1914 3460
rect 2778 2644 2834 2680
rect 2778 2624 2780 2644
rect 2780 2624 2832 2644
rect 2832 2624 2834 2644
rect 12346 16632 12402 16688
rect 4066 15408 4122 15464
rect 4066 15000 4122 15056
rect 3698 14184 3754 14240
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 3698 13368 3754 13424
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3422 12960 3478 13016
rect 3606 12552 3662 12608
rect 3422 9560 3478 9616
rect 3422 7792 3478 7848
rect 3054 6160 3110 6216
rect 2962 1808 3018 1864
rect 3330 3032 3386 3088
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3698 10920 3754 10976
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 3606 9016 3662 9072
rect 3606 8472 3662 8528
rect 3606 7964 3608 7984
rect 3608 7964 3660 7984
rect 3660 7964 3662 7984
rect 3606 7928 3662 7964
rect 4066 10104 4122 10160
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 4158 8880 4214 8936
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 4066 7112 4122 7168
rect 3606 6296 3662 6352
rect 3882 6740 3884 6760
rect 3884 6740 3936 6760
rect 3936 6740 3938 6760
rect 3882 6704 3938 6740
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 3422 2252 3424 2272
rect 3424 2252 3476 2272
rect 3476 2252 3478 2272
rect 3422 2216 3478 2252
rect 3514 1400 3570 1456
rect 3330 992 3386 1048
rect 3238 584 3294 640
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 3790 3576 3846 3632
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 4802 10512 4858 10568
rect 4710 9424 4766 9480
rect 4618 5752 4674 5808
rect 5630 11872 5686 11928
rect 5354 11600 5410 11656
rect 5170 9968 5226 10024
rect 5630 10512 5686 10568
rect 5446 8880 5502 8936
rect 5538 8336 5594 8392
rect 5354 4120 5410 4176
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 5998 11736 6054 11792
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 5998 5752 6054 5808
rect 6182 7520 6238 7576
rect 6366 9288 6422 9344
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 8114 13368 8170 13424
rect 7562 11636 7564 11656
rect 7564 11636 7616 11656
rect 7616 11636 7618 11656
rect 7562 11600 7618 11636
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6734 6704 6790 6760
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 7562 9016 7618 9072
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 8298 10140 8300 10160
rect 8300 10140 8352 10160
rect 8352 10140 8354 10160
rect 8298 10104 8354 10140
rect 8390 9832 8446 9888
rect 8482 9696 8538 9752
rect 8482 7948 8538 7984
rect 8482 7928 8484 7948
rect 8484 7928 8536 7948
rect 8536 7928 8538 7948
rect 8390 7792 8446 7848
rect 8390 6840 8446 6896
rect 8022 5616 8078 5672
rect 8574 6568 8630 6624
rect 8114 3576 8170 3632
rect 8942 12144 8998 12200
rect 8758 11192 8814 11248
rect 8850 10376 8906 10432
rect 9126 11600 9182 11656
rect 8850 6840 8906 6896
rect 9034 8200 9090 8256
rect 9586 11892 9642 11928
rect 9586 11872 9588 11892
rect 9588 11872 9640 11892
rect 9640 11872 9642 11892
rect 9586 11736 9642 11792
rect 9310 8880 9366 8936
rect 9678 11056 9734 11112
rect 9678 8744 9734 8800
rect 9586 8336 9642 8392
rect 9310 6160 9366 6216
rect 9218 4800 9274 4856
rect 9310 4120 9366 4176
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 10138 10648 10194 10704
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 10138 9324 10140 9344
rect 10140 9324 10192 9344
rect 10192 9324 10194 9344
rect 10138 9288 10194 9324
rect 10046 9016 10102 9072
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10046 7792 10102 7848
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9954 3460 10010 3496
rect 9954 3440 9956 3460
rect 9956 3440 10008 3460
rect 10008 3440 10010 3460
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 10782 8880 10838 8936
rect 10782 7792 10838 7848
rect 10506 6432 10562 6488
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 10690 6296 10746 6352
rect 11150 13776 11206 13832
rect 11058 10376 11114 10432
rect 11058 8744 11114 8800
rect 11150 4700 11152 4720
rect 11152 4700 11204 4720
rect 11204 4700 11206 4720
rect 11150 4664 11206 4700
rect 11058 3032 11114 3088
rect 12162 11464 12218 11520
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 12254 10648 12310 10704
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 13450 13640 13506 13696
rect 12438 11600 12494 11656
rect 12254 10104 12310 10160
rect 12162 9288 12218 9344
rect 12070 8236 12072 8256
rect 12072 8236 12124 8256
rect 12124 8236 12126 8256
rect 12070 8200 12126 8236
rect 12162 5788 12164 5808
rect 12164 5788 12216 5808
rect 12216 5788 12218 5808
rect 12162 5752 12218 5788
rect 12070 4800 12126 4856
rect 12438 6704 12494 6760
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12990 10804 13046 10840
rect 12990 10784 12992 10804
rect 12992 10784 13044 10804
rect 13044 10784 13046 10804
rect 12622 10240 12678 10296
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12714 9968 12770 10024
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 13082 9016 13138 9072
rect 12622 8200 12678 8256
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 11794 1808 11850 1864
rect 12346 3440 12402 3496
rect 13082 7792 13138 7848
rect 13266 8608 13322 8664
rect 12990 7268 13046 7304
rect 12990 7248 12992 7268
rect 12992 7248 13044 7268
rect 13044 7248 13046 7268
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 13082 6840 13138 6896
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 12254 2896 12310 2952
rect 12990 3168 13046 3224
rect 13082 2916 13138 2952
rect 13082 2896 13084 2916
rect 13084 2896 13136 2916
rect 13136 2896 13138 2916
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 13358 3984 13414 4040
rect 13634 13232 13690 13288
rect 13542 11736 13598 11792
rect 13910 14592 13966 14648
rect 13818 13640 13874 13696
rect 13818 12280 13874 12336
rect 13818 10648 13874 10704
rect 13542 7656 13598 7712
rect 13542 7384 13598 7440
rect 13634 6840 13690 6896
rect 13910 9288 13966 9344
rect 14002 9152 14058 9208
rect 13818 9036 13874 9072
rect 13818 9016 13820 9036
rect 13820 9016 13872 9036
rect 13872 9016 13874 9036
rect 14094 8880 14150 8936
rect 14094 7928 14150 7984
rect 13910 7384 13966 7440
rect 13818 4800 13874 4856
rect 13818 4256 13874 4312
rect 13726 4120 13782 4176
rect 13726 3984 13782 4040
rect 14370 11328 14426 11384
rect 14278 2624 14334 2680
rect 3054 176 3110 232
rect 14646 10648 14702 10704
rect 14554 8336 14610 8392
rect 14738 5616 14794 5672
rect 14554 4004 14610 4040
rect 14554 3984 14556 4004
rect 14556 3984 14608 4004
rect 14608 3984 14610 4004
rect 15382 15000 15438 15056
rect 15934 16224 15990 16280
rect 16210 14184 16266 14240
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 15658 13640 15714 13696
rect 15014 13096 15070 13152
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15198 11600 15254 11656
rect 15106 11056 15162 11112
rect 15106 9968 15162 10024
rect 15014 8608 15070 8664
rect 15566 12144 15622 12200
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 15934 11192 15990 11248
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 16118 10240 16174 10296
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 16118 9560 16174 9616
rect 15290 8744 15346 8800
rect 15290 8200 15346 8256
rect 15106 5480 15162 5536
rect 15198 3576 15254 3632
rect 15198 2644 15254 2680
rect 15198 2624 15200 2644
rect 15200 2624 15252 2644
rect 15252 2624 15254 2644
rect 15474 6840 15530 6896
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 16394 13640 16450 13696
rect 18418 15816 18474 15872
rect 17866 13388 17922 13424
rect 17866 13368 17868 13388
rect 17868 13368 17920 13388
rect 17920 13368 17922 13388
rect 17866 12824 17922 12880
rect 16486 12280 16542 12336
rect 15750 8472 15806 8528
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15658 6296 15714 6352
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 16302 8336 16358 8392
rect 16302 5344 16358 5400
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 15934 4140 15990 4176
rect 15934 4120 15936 4140
rect 15936 4120 15988 4140
rect 15988 4120 15990 4140
rect 15934 3848 15990 3904
rect 15842 3732 15898 3768
rect 15842 3712 15844 3732
rect 15844 3712 15896 3732
rect 15896 3712 15898 3732
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 15658 3032 15714 3088
rect 15934 2916 15990 2952
rect 15934 2896 15936 2916
rect 15936 2896 15988 2916
rect 15988 2896 15990 2916
rect 15290 1400 15346 1456
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 16486 9016 16542 9072
rect 16854 10104 16910 10160
rect 16578 7384 16634 7440
rect 16486 5072 16542 5128
rect 16302 2216 16358 2272
rect 17222 10240 17278 10296
rect 17222 9444 17278 9480
rect 17222 9424 17224 9444
rect 17224 9424 17276 9444
rect 17276 9424 17278 9444
rect 17222 9288 17278 9344
rect 17406 8200 17462 8256
rect 17498 7792 17554 7848
rect 17406 6976 17462 7032
rect 17130 4664 17186 4720
rect 16394 992 16450 1048
rect 17866 11600 17922 11656
rect 17682 6432 17738 6488
rect 17498 6160 17554 6216
rect 17314 5616 17370 5672
rect 17406 4800 17462 4856
rect 17222 584 17278 640
rect 17682 5908 17738 5944
rect 17682 5888 17684 5908
rect 17684 5888 17736 5908
rect 17736 5888 17738 5908
rect 17682 3984 17738 4040
rect 18050 6976 18106 7032
rect 18234 6024 18290 6080
rect 18694 13232 18750 13288
rect 18510 10784 18566 10840
rect 18602 10512 18658 10568
rect 18142 5208 18198 5264
rect 17866 4392 17922 4448
rect 18694 9696 18750 9752
rect 18970 5652 18972 5672
rect 18972 5652 19024 5672
rect 19024 5652 19026 5672
rect 18970 5616 19026 5652
rect 14462 176 14518 232
<< metal3 >>
rect 0 16690 480 16720
rect 3693 16690 3759 16693
rect 0 16688 3759 16690
rect 0 16632 3698 16688
rect 3754 16632 3759 16688
rect 0 16630 3759 16632
rect 0 16600 480 16630
rect 3693 16627 3759 16630
rect 12341 16690 12407 16693
rect 19520 16690 20000 16720
rect 12341 16688 20000 16690
rect 12341 16632 12346 16688
rect 12402 16632 20000 16688
rect 12341 16630 20000 16632
rect 12341 16627 12407 16630
rect 19520 16600 20000 16630
rect 0 16282 480 16312
rect 2589 16282 2655 16285
rect 0 16280 2655 16282
rect 0 16224 2594 16280
rect 2650 16224 2655 16280
rect 0 16222 2655 16224
rect 0 16192 480 16222
rect 2589 16219 2655 16222
rect 15929 16282 15995 16285
rect 19520 16282 20000 16312
rect 15929 16280 20000 16282
rect 15929 16224 15934 16280
rect 15990 16224 20000 16280
rect 15929 16222 20000 16224
rect 15929 16219 15995 16222
rect 19520 16192 20000 16222
rect 0 15874 480 15904
rect 3325 15874 3391 15877
rect 0 15872 3391 15874
rect 0 15816 3330 15872
rect 3386 15816 3391 15872
rect 0 15814 3391 15816
rect 0 15784 480 15814
rect 3325 15811 3391 15814
rect 18413 15874 18479 15877
rect 19520 15874 20000 15904
rect 18413 15872 20000 15874
rect 18413 15816 18418 15872
rect 18474 15816 20000 15872
rect 18413 15814 20000 15816
rect 18413 15811 18479 15814
rect 19520 15784 20000 15814
rect 0 15466 480 15496
rect 4061 15466 4127 15469
rect 0 15464 4127 15466
rect 0 15408 4066 15464
rect 4122 15408 4127 15464
rect 0 15406 4127 15408
rect 0 15376 480 15406
rect 4061 15403 4127 15406
rect 16430 15404 16436 15468
rect 16500 15466 16506 15468
rect 19520 15466 20000 15496
rect 16500 15406 20000 15466
rect 16500 15404 16506 15406
rect 19520 15376 20000 15406
rect 0 15058 480 15088
rect 4061 15058 4127 15061
rect 0 15056 4127 15058
rect 0 15000 4066 15056
rect 4122 15000 4127 15056
rect 0 14998 4127 15000
rect 0 14968 480 14998
rect 4061 14995 4127 14998
rect 15377 15058 15443 15061
rect 19520 15058 20000 15088
rect 15377 15056 20000 15058
rect 15377 15000 15382 15056
rect 15438 15000 20000 15056
rect 15377 14998 20000 15000
rect 15377 14995 15443 14998
rect 19520 14968 20000 14998
rect 6874 14720 7194 14721
rect 0 14650 480 14680
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 14655 13125 14656
rect 3141 14650 3207 14653
rect 0 14648 3207 14650
rect 0 14592 3146 14648
rect 3202 14592 3207 14648
rect 0 14590 3207 14592
rect 0 14560 480 14590
rect 3141 14587 3207 14590
rect 13905 14650 13971 14653
rect 19520 14650 20000 14680
rect 13905 14648 20000 14650
rect 13905 14592 13910 14648
rect 13966 14592 20000 14648
rect 13905 14590 20000 14592
rect 13905 14587 13971 14590
rect 19520 14560 20000 14590
rect 0 14242 480 14272
rect 3693 14242 3759 14245
rect 0 14240 3759 14242
rect 0 14184 3698 14240
rect 3754 14184 3759 14240
rect 0 14182 3759 14184
rect 0 14152 480 14182
rect 3693 14179 3759 14182
rect 16205 14242 16271 14245
rect 19520 14242 20000 14272
rect 16205 14240 20000 14242
rect 16205 14184 16210 14240
rect 16266 14184 20000 14240
rect 16205 14182 20000 14184
rect 16205 14179 16271 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19520 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13834 480 13864
rect 2681 13834 2747 13837
rect 0 13832 2747 13834
rect 0 13776 2686 13832
rect 2742 13776 2747 13832
rect 0 13774 2747 13776
rect 0 13744 480 13774
rect 2681 13771 2747 13774
rect 11145 13834 11211 13837
rect 19520 13834 20000 13864
rect 11145 13832 20000 13834
rect 11145 13776 11150 13832
rect 11206 13776 20000 13832
rect 11145 13774 20000 13776
rect 11145 13771 11211 13774
rect 19520 13744 20000 13774
rect 13445 13700 13511 13701
rect 13445 13696 13492 13700
rect 13556 13698 13562 13700
rect 13813 13698 13879 13701
rect 14774 13698 14780 13700
rect 13445 13640 13450 13696
rect 13445 13636 13492 13640
rect 13556 13638 13602 13698
rect 13813 13696 14780 13698
rect 13813 13640 13818 13696
rect 13874 13640 14780 13696
rect 13813 13638 14780 13640
rect 13556 13636 13562 13638
rect 13445 13635 13511 13636
rect 13813 13635 13879 13638
rect 14774 13636 14780 13638
rect 14844 13636 14850 13700
rect 15653 13698 15719 13701
rect 16389 13698 16455 13701
rect 16614 13698 16620 13700
rect 15653 13696 16620 13698
rect 15653 13640 15658 13696
rect 15714 13640 16394 13696
rect 16450 13640 16620 13696
rect 15653 13638 16620 13640
rect 15653 13635 15719 13638
rect 16389 13635 16455 13638
rect 16614 13636 16620 13638
rect 16684 13636 16690 13700
rect 6874 13632 7194 13633
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 0 13426 480 13456
rect 3693 13426 3759 13429
rect 0 13424 3759 13426
rect 0 13368 3698 13424
rect 3754 13368 3759 13424
rect 0 13366 3759 13368
rect 0 13336 480 13366
rect 3693 13363 3759 13366
rect 8109 13426 8175 13429
rect 17718 13426 17724 13428
rect 8109 13424 17724 13426
rect 8109 13368 8114 13424
rect 8170 13368 17724 13424
rect 8109 13366 17724 13368
rect 8109 13363 8175 13366
rect 17718 13364 17724 13366
rect 17788 13426 17794 13428
rect 17861 13426 17927 13429
rect 17788 13424 17927 13426
rect 17788 13368 17866 13424
rect 17922 13368 17927 13424
rect 17788 13366 17927 13368
rect 17788 13364 17794 13366
rect 17861 13363 17927 13366
rect 13629 13292 13695 13293
rect 13629 13288 13676 13292
rect 13740 13290 13746 13292
rect 18689 13290 18755 13293
rect 19520 13290 20000 13320
rect 13629 13232 13634 13288
rect 13629 13228 13676 13232
rect 13740 13230 13786 13290
rect 18689 13288 20000 13290
rect 18689 13232 18694 13288
rect 18750 13232 20000 13288
rect 18689 13230 20000 13232
rect 13740 13228 13746 13230
rect 13629 13227 13695 13228
rect 18689 13227 18755 13230
rect 19520 13200 20000 13230
rect 14406 13092 14412 13156
rect 14476 13154 14482 13156
rect 15009 13154 15075 13157
rect 14476 13152 15075 13154
rect 14476 13096 15014 13152
rect 15070 13096 15075 13152
rect 14476 13094 15075 13096
rect 14476 13092 14482 13094
rect 15009 13091 15075 13094
rect 3909 13088 4229 13089
rect 0 13018 480 13048
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 3417 13018 3483 13021
rect 0 13016 3483 13018
rect 0 12960 3422 13016
rect 3478 12960 3483 13016
rect 0 12958 3483 12960
rect 0 12928 480 12958
rect 3417 12955 3483 12958
rect 17861 12882 17927 12885
rect 19520 12882 20000 12912
rect 17861 12880 20000 12882
rect 17861 12824 17866 12880
rect 17922 12824 20000 12880
rect 17861 12822 20000 12824
rect 17861 12819 17927 12822
rect 19520 12792 20000 12822
rect 0 12610 480 12640
rect 3601 12610 3667 12613
rect 0 12608 3667 12610
rect 0 12552 3606 12608
rect 3662 12552 3667 12608
rect 0 12550 3667 12552
rect 0 12520 480 12550
rect 3601 12547 3667 12550
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 12479 13125 12480
rect 15142 12412 15148 12476
rect 15212 12474 15218 12476
rect 19520 12474 20000 12504
rect 15212 12414 20000 12474
rect 15212 12412 15218 12414
rect 19520 12384 20000 12414
rect 3141 12338 3207 12341
rect 13813 12338 13879 12341
rect 3141 12336 13879 12338
rect 3141 12280 3146 12336
rect 3202 12280 13818 12336
rect 13874 12280 13879 12336
rect 3141 12278 13879 12280
rect 3141 12275 3207 12278
rect 13813 12275 13879 12278
rect 16246 12276 16252 12340
rect 16316 12338 16322 12340
rect 16481 12338 16547 12341
rect 16316 12336 16547 12338
rect 16316 12280 16486 12336
rect 16542 12280 16547 12336
rect 16316 12278 16547 12280
rect 16316 12276 16322 12278
rect 16481 12275 16547 12278
rect 0 12202 480 12232
rect 8937 12202 9003 12205
rect 0 12200 9003 12202
rect 0 12144 8942 12200
rect 8998 12144 9003 12200
rect 0 12142 9003 12144
rect 0 12112 480 12142
rect 8937 12139 9003 12142
rect 15561 12202 15627 12205
rect 15561 12200 16314 12202
rect 15561 12144 15566 12200
rect 15622 12144 16314 12200
rect 15561 12142 16314 12144
rect 15561 12139 15627 12142
rect 16254 12066 16314 12142
rect 19520 12066 20000 12096
rect 16254 12006 20000 12066
rect 3909 12000 4229 12001
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 19520 11976 20000 12006
rect 15770 11935 16090 11936
rect 5625 11930 5691 11933
rect 9581 11930 9647 11933
rect 5625 11928 9647 11930
rect 5625 11872 5630 11928
rect 5686 11872 9586 11928
rect 9642 11872 9647 11928
rect 5625 11870 9647 11872
rect 5625 11867 5691 11870
rect 9581 11867 9647 11870
rect 0 11794 480 11824
rect 5993 11794 6059 11797
rect 9581 11794 9647 11797
rect 0 11792 9647 11794
rect 0 11736 5998 11792
rect 6054 11736 9586 11792
rect 9642 11736 9647 11792
rect 0 11734 9647 11736
rect 0 11704 480 11734
rect 5993 11731 6059 11734
rect 9581 11731 9647 11734
rect 13302 11732 13308 11796
rect 13372 11794 13378 11796
rect 13537 11794 13603 11797
rect 13372 11792 13603 11794
rect 13372 11736 13542 11792
rect 13598 11736 13603 11792
rect 13372 11734 13603 11736
rect 13372 11732 13378 11734
rect 13537 11731 13603 11734
rect 5349 11658 5415 11661
rect 7557 11658 7623 11661
rect 9121 11660 9187 11661
rect 12433 11660 12499 11661
rect 5349 11656 7623 11658
rect 5349 11600 5354 11656
rect 5410 11600 7562 11656
rect 7618 11600 7623 11656
rect 5349 11598 7623 11600
rect 5349 11595 5415 11598
rect 7557 11595 7623 11598
rect 9070 11596 9076 11660
rect 9140 11658 9187 11660
rect 9140 11656 9232 11658
rect 9182 11600 9232 11656
rect 9140 11598 9232 11600
rect 9140 11596 9187 11598
rect 12382 11596 12388 11660
rect 12452 11658 12499 11660
rect 15193 11658 15259 11661
rect 17861 11658 17927 11661
rect 19520 11658 20000 11688
rect 12452 11656 12544 11658
rect 12494 11600 12544 11656
rect 12452 11598 12544 11600
rect 15193 11656 20000 11658
rect 15193 11600 15198 11656
rect 15254 11600 17866 11656
rect 17922 11600 20000 11656
rect 15193 11598 20000 11600
rect 12452 11596 12499 11598
rect 9121 11595 9187 11596
rect 12433 11595 12499 11596
rect 15193 11595 15259 11598
rect 17861 11595 17927 11598
rect 19520 11568 20000 11598
rect 12157 11524 12223 11525
rect 12157 11522 12204 11524
rect 12112 11520 12204 11522
rect 12112 11464 12162 11520
rect 12112 11462 12204 11464
rect 12157 11460 12204 11462
rect 12268 11460 12274 11524
rect 12157 11459 12223 11460
rect 6874 11456 7194 11457
rect 0 11386 480 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 2957 11386 3023 11389
rect 0 11384 3023 11386
rect 0 11328 2962 11384
rect 3018 11328 3023 11384
rect 0 11326 3023 11328
rect 0 11296 480 11326
rect 2957 11323 3023 11326
rect 14222 11324 14228 11388
rect 14292 11386 14298 11388
rect 14365 11386 14431 11389
rect 14292 11384 14431 11386
rect 14292 11328 14370 11384
rect 14426 11328 14431 11384
rect 14292 11326 14431 11328
rect 14292 11324 14298 11326
rect 14365 11323 14431 11326
rect 8518 11188 8524 11252
rect 8588 11250 8594 11252
rect 8753 11250 8819 11253
rect 8588 11248 8819 11250
rect 8588 11192 8758 11248
rect 8814 11192 8819 11248
rect 8588 11190 8819 11192
rect 8588 11188 8594 11190
rect 8753 11187 8819 11190
rect 15929 11250 15995 11253
rect 19520 11250 20000 11280
rect 15929 11248 20000 11250
rect 15929 11192 15934 11248
rect 15990 11192 20000 11248
rect 15929 11190 20000 11192
rect 15929 11187 15995 11190
rect 19520 11160 20000 11190
rect 9673 11114 9739 11117
rect 15101 11114 15167 11117
rect 9673 11112 15167 11114
rect 9673 11056 9678 11112
rect 9734 11056 15106 11112
rect 15162 11056 15167 11112
rect 9673 11054 15167 11056
rect 9673 11051 9739 11054
rect 15101 11051 15167 11054
rect 0 10978 480 11008
rect 3693 10978 3759 10981
rect 0 10976 3759 10978
rect 0 10920 3698 10976
rect 3754 10920 3759 10976
rect 0 10918 3759 10920
rect 0 10888 480 10918
rect 3693 10915 3759 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 11646 10780 11652 10844
rect 11716 10842 11722 10844
rect 12985 10842 13051 10845
rect 11716 10840 13051 10842
rect 11716 10784 12990 10840
rect 13046 10784 13051 10840
rect 11716 10782 13051 10784
rect 11716 10780 11722 10782
rect 12985 10779 13051 10782
rect 18505 10842 18571 10845
rect 19520 10842 20000 10872
rect 18505 10840 20000 10842
rect 18505 10784 18510 10840
rect 18566 10784 20000 10840
rect 18505 10782 20000 10784
rect 18505 10779 18571 10782
rect 19520 10752 20000 10782
rect 10133 10706 10199 10709
rect 12249 10706 12315 10709
rect 12566 10706 12572 10708
rect 10133 10704 10978 10706
rect 10133 10648 10138 10704
rect 10194 10648 10978 10704
rect 10133 10646 10978 10648
rect 10133 10643 10199 10646
rect 0 10570 480 10600
rect 4797 10570 4863 10573
rect 0 10568 4863 10570
rect 0 10512 4802 10568
rect 4858 10512 4863 10568
rect 0 10510 4863 10512
rect 0 10480 480 10510
rect 4797 10507 4863 10510
rect 5625 10570 5691 10573
rect 10918 10570 10978 10646
rect 12249 10704 12572 10706
rect 12249 10648 12254 10704
rect 12310 10648 12572 10704
rect 12249 10646 12572 10648
rect 12249 10643 12315 10646
rect 12566 10644 12572 10646
rect 12636 10706 12642 10708
rect 13813 10706 13879 10709
rect 12636 10704 13879 10706
rect 12636 10648 13818 10704
rect 13874 10648 13879 10704
rect 12636 10646 13879 10648
rect 12636 10644 12642 10646
rect 13813 10643 13879 10646
rect 14641 10706 14707 10709
rect 14641 10704 15762 10706
rect 14641 10648 14646 10704
rect 14702 10648 15762 10704
rect 14641 10646 15762 10648
rect 14641 10643 14707 10646
rect 15702 10570 15762 10646
rect 18597 10570 18663 10573
rect 5625 10568 10794 10570
rect 5625 10512 5630 10568
rect 5686 10512 10794 10568
rect 5625 10510 10794 10512
rect 10918 10510 13370 10570
rect 15702 10568 18663 10570
rect 15702 10512 18602 10568
rect 18658 10512 18663 10568
rect 15702 10510 18663 10512
rect 5625 10507 5691 10510
rect 8845 10434 8911 10437
rect 8526 10432 8911 10434
rect 8526 10376 8850 10432
rect 8906 10376 8911 10432
rect 8526 10374 8911 10376
rect 10734 10434 10794 10510
rect 11053 10434 11119 10437
rect 10734 10432 11119 10434
rect 10734 10376 11058 10432
rect 11114 10376 11119 10432
rect 10734 10374 11119 10376
rect 13310 10434 13370 10510
rect 18597 10507 18663 10510
rect 19520 10434 20000 10464
rect 13310 10374 20000 10434
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 8526 10196 8586 10374
rect 8845 10371 8911 10374
rect 11053 10371 11119 10374
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19520 10344 20000 10374
rect 12805 10303 13125 10304
rect 12014 10236 12020 10300
rect 12084 10298 12090 10300
rect 12617 10298 12683 10301
rect 12084 10296 12683 10298
rect 12084 10240 12622 10296
rect 12678 10240 12683 10296
rect 12084 10238 12683 10240
rect 12084 10236 12090 10238
rect 12617 10235 12683 10238
rect 16113 10298 16179 10301
rect 16798 10298 16804 10300
rect 16113 10296 16804 10298
rect 16113 10240 16118 10296
rect 16174 10240 16804 10296
rect 16113 10238 16804 10240
rect 16113 10235 16179 10238
rect 16798 10236 16804 10238
rect 16868 10236 16874 10300
rect 17217 10298 17283 10301
rect 17174 10296 17283 10298
rect 17174 10240 17222 10296
rect 17278 10240 17283 10296
rect 17174 10235 17283 10240
rect 0 10162 480 10192
rect 8342 10165 8586 10196
rect 4061 10162 4127 10165
rect 0 10160 4127 10162
rect 0 10104 4066 10160
rect 4122 10104 4127 10160
rect 0 10102 4127 10104
rect 0 10072 480 10102
rect 4061 10099 4127 10102
rect 8293 10160 8586 10165
rect 8293 10104 8298 10160
rect 8354 10136 8586 10160
rect 12249 10160 12315 10165
rect 8354 10104 8402 10136
rect 8293 10102 8402 10104
rect 12249 10104 12254 10160
rect 12310 10104 12315 10160
rect 8293 10099 8359 10102
rect 12249 10099 12315 10104
rect 16849 10162 16915 10165
rect 17174 10162 17234 10235
rect 16849 10160 17234 10162
rect 16849 10104 16854 10160
rect 16910 10104 17234 10160
rect 16849 10102 17234 10104
rect 16849 10099 16915 10102
rect 2957 10026 3023 10029
rect 5165 10026 5231 10029
rect 2957 10024 5231 10026
rect 2957 9968 2962 10024
rect 3018 9968 5170 10024
rect 5226 9968 5231 10024
rect 2957 9966 5231 9968
rect 12252 10026 12312 10099
rect 12709 10026 12775 10029
rect 12252 10024 12775 10026
rect 12252 9968 12714 10024
rect 12770 9968 12775 10024
rect 12252 9966 12775 9968
rect 2957 9963 3023 9966
rect 5165 9963 5231 9966
rect 12709 9963 12775 9966
rect 15101 10026 15167 10029
rect 15101 10024 16314 10026
rect 15101 9968 15106 10024
rect 15162 9968 16314 10024
rect 15101 9966 16314 9968
rect 15101 9963 15167 9966
rect 8385 9890 8451 9893
rect 8518 9890 8524 9892
rect 8385 9888 8524 9890
rect 8385 9832 8390 9888
rect 8446 9832 8524 9888
rect 8385 9830 8524 9832
rect 8385 9827 8451 9830
rect 8518 9828 8524 9830
rect 8588 9828 8594 9892
rect 16254 9890 16314 9966
rect 19520 9890 20000 9920
rect 16254 9830 20000 9890
rect 3909 9824 4229 9825
rect 0 9754 480 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 19520 9800 20000 9830
rect 15770 9759 16090 9760
rect 2957 9754 3023 9757
rect 0 9752 3023 9754
rect 0 9696 2962 9752
rect 3018 9696 3023 9752
rect 0 9694 3023 9696
rect 0 9664 480 9694
rect 2957 9691 3023 9694
rect 8477 9754 8543 9757
rect 9070 9754 9076 9756
rect 8477 9752 9076 9754
rect 8477 9696 8482 9752
rect 8538 9696 9076 9752
rect 8477 9694 9076 9696
rect 8477 9691 8543 9694
rect 9070 9692 9076 9694
rect 9140 9692 9146 9756
rect 18689 9754 18755 9757
rect 16254 9752 18755 9754
rect 16254 9696 18694 9752
rect 18750 9696 18755 9752
rect 16254 9694 18755 9696
rect 3417 9618 3483 9621
rect 16113 9618 16179 9621
rect 3417 9616 16179 9618
rect 3417 9560 3422 9616
rect 3478 9560 16118 9616
rect 16174 9560 16179 9616
rect 3417 9558 16179 9560
rect 3417 9555 3483 9558
rect 16113 9555 16179 9558
rect 4705 9482 4771 9485
rect 4705 9480 15210 9482
rect 4705 9424 4710 9480
rect 4766 9424 15210 9480
rect 4705 9422 15210 9424
rect 4705 9419 4771 9422
rect 0 9346 480 9376
rect 6361 9346 6427 9349
rect 0 9344 6427 9346
rect 0 9288 6366 9344
rect 6422 9288 6427 9344
rect 0 9286 6427 9288
rect 0 9256 480 9286
rect 6361 9283 6427 9286
rect 10133 9346 10199 9349
rect 12157 9346 12223 9349
rect 13905 9348 13971 9349
rect 13854 9346 13860 9348
rect 10133 9344 12223 9346
rect 10133 9288 10138 9344
rect 10194 9288 12162 9344
rect 12218 9288 12223 9344
rect 10133 9286 12223 9288
rect 13814 9286 13860 9346
rect 13924 9344 13971 9348
rect 13966 9288 13971 9344
rect 10133 9283 10199 9286
rect 12157 9283 12223 9286
rect 13854 9284 13860 9286
rect 13924 9284 13971 9288
rect 15150 9346 15210 9422
rect 15326 9420 15332 9484
rect 15396 9482 15402 9484
rect 16254 9482 16314 9694
rect 17220 9485 17280 9694
rect 18689 9691 18755 9694
rect 15396 9422 16314 9482
rect 17217 9480 17283 9485
rect 19520 9482 20000 9512
rect 17217 9424 17222 9480
rect 17278 9424 17283 9480
rect 15396 9420 15402 9422
rect 17217 9419 17283 9424
rect 17358 9422 20000 9482
rect 17217 9346 17283 9349
rect 15150 9344 17283 9346
rect 15150 9288 17222 9344
rect 17278 9288 17283 9344
rect 15150 9286 17283 9288
rect 13905 9283 13971 9284
rect 17217 9283 17283 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 13997 9212 14063 9213
rect 13997 9208 14044 9212
rect 14108 9210 14114 9212
rect 17358 9210 17418 9422
rect 19520 9392 20000 9422
rect 13997 9152 14002 9208
rect 13997 9148 14044 9152
rect 14108 9150 14154 9210
rect 14230 9150 17418 9210
rect 14108 9148 14114 9150
rect 13997 9147 14063 9148
rect 3601 9074 3667 9077
rect 7557 9074 7623 9077
rect 3601 9072 7623 9074
rect 3601 9016 3606 9072
rect 3662 9016 7562 9072
rect 7618 9016 7623 9072
rect 3601 9014 7623 9016
rect 3601 9011 3667 9014
rect 7557 9011 7623 9014
rect 10041 9074 10107 9077
rect 13077 9074 13143 9077
rect 10041 9072 13143 9074
rect 10041 9016 10046 9072
rect 10102 9016 13082 9072
rect 13138 9016 13143 9072
rect 10041 9014 13143 9016
rect 10041 9011 10107 9014
rect 13077 9011 13143 9014
rect 13813 9074 13879 9077
rect 14230 9074 14290 9150
rect 13813 9072 14290 9074
rect 13813 9016 13818 9072
rect 13874 9016 14290 9072
rect 13813 9014 14290 9016
rect 16481 9074 16547 9077
rect 19520 9074 20000 9104
rect 16481 9072 20000 9074
rect 16481 9016 16486 9072
rect 16542 9016 20000 9072
rect 16481 9014 20000 9016
rect 13813 9011 13879 9014
rect 0 8938 480 8968
rect 14046 8941 14106 9014
rect 16481 9011 16547 9014
rect 19520 8984 20000 9014
rect 4153 8938 4219 8941
rect 5441 8938 5507 8941
rect 9305 8938 9371 8941
rect 10777 8938 10843 8941
rect 0 8936 9371 8938
rect 0 8880 4158 8936
rect 4214 8880 5446 8936
rect 5502 8880 9310 8936
rect 9366 8880 9371 8936
rect 0 8878 9371 8880
rect 0 8848 480 8878
rect 4153 8875 4219 8878
rect 5441 8875 5507 8878
rect 9305 8875 9371 8878
rect 9676 8936 10843 8938
rect 9676 8880 10782 8936
rect 10838 8880 10843 8936
rect 9676 8878 10843 8880
rect 14046 8936 14155 8941
rect 14046 8880 14094 8936
rect 14150 8880 14155 8936
rect 14046 8878 14155 8880
rect 9676 8805 9736 8878
rect 10777 8875 10843 8878
rect 14089 8875 14155 8878
rect 9673 8800 9739 8805
rect 9673 8744 9678 8800
rect 9734 8744 9739 8800
rect 9673 8739 9739 8744
rect 11053 8802 11119 8805
rect 15285 8802 15351 8805
rect 11053 8800 15351 8802
rect 11053 8744 11058 8800
rect 11114 8744 15290 8800
rect 15346 8744 15351 8800
rect 11053 8742 15351 8744
rect 11053 8739 11119 8742
rect 15285 8739 15351 8742
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 8671 16090 8672
rect 12014 8604 12020 8668
rect 12084 8666 12090 8668
rect 13261 8666 13327 8669
rect 15009 8668 15075 8669
rect 12084 8664 13327 8666
rect 12084 8608 13266 8664
rect 13322 8608 13327 8664
rect 12084 8606 13327 8608
rect 12084 8604 12090 8606
rect 13261 8603 13327 8606
rect 14958 8604 14964 8668
rect 15028 8666 15075 8668
rect 19520 8666 20000 8696
rect 15028 8664 15120 8666
rect 15070 8608 15120 8664
rect 15028 8606 15120 8608
rect 16208 8606 20000 8666
rect 15028 8604 15075 8606
rect 15009 8603 15075 8604
rect 3601 8530 3667 8533
rect 15326 8530 15332 8532
rect 3601 8528 15332 8530
rect 3601 8472 3606 8528
rect 3662 8472 15332 8528
rect 3601 8470 15332 8472
rect 3601 8467 3667 8470
rect 15326 8468 15332 8470
rect 15396 8468 15402 8532
rect 15745 8530 15811 8533
rect 16208 8530 16268 8606
rect 19520 8576 20000 8606
rect 15702 8528 16268 8530
rect 15702 8472 15750 8528
rect 15806 8472 16268 8528
rect 15702 8470 16268 8472
rect 15702 8467 15811 8470
rect 0 8394 480 8424
rect 2865 8394 2931 8397
rect 0 8392 2931 8394
rect 0 8336 2870 8392
rect 2926 8336 2931 8392
rect 0 8334 2931 8336
rect 0 8304 480 8334
rect 2865 8331 2931 8334
rect 5390 8332 5396 8396
rect 5460 8394 5466 8396
rect 5533 8394 5599 8397
rect 5460 8392 5599 8394
rect 5460 8336 5538 8392
rect 5594 8336 5599 8392
rect 5460 8334 5599 8336
rect 5460 8332 5466 8334
rect 5533 8331 5599 8334
rect 9581 8394 9647 8397
rect 14549 8396 14615 8397
rect 14549 8394 14596 8396
rect 9581 8392 14336 8394
rect 9581 8336 9586 8392
rect 9642 8336 14336 8392
rect 9581 8334 14336 8336
rect 14504 8392 14596 8394
rect 14504 8336 14554 8392
rect 14504 8334 14596 8336
rect 9581 8331 9647 8334
rect 9029 8258 9095 8261
rect 9029 8256 9874 8258
rect 9029 8200 9034 8256
rect 9090 8200 9874 8256
rect 9029 8198 9874 8200
rect 9029 8195 9095 8198
rect 6874 8192 7194 8193
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 0 7986 480 8016
rect 1761 7986 1827 7989
rect 0 7984 1827 7986
rect 0 7928 1766 7984
rect 1822 7928 1827 7984
rect 0 7926 1827 7928
rect 0 7896 480 7926
rect 1761 7923 1827 7926
rect 3601 7986 3667 7989
rect 8477 7986 8543 7989
rect 3601 7984 8543 7986
rect 3601 7928 3606 7984
rect 3662 7928 8482 7984
rect 8538 7928 8543 7984
rect 3601 7926 8543 7928
rect 9814 7986 9874 8198
rect 11830 8196 11836 8260
rect 11900 8258 11906 8260
rect 12065 8258 12131 8261
rect 12617 8258 12683 8261
rect 11900 8256 12131 8258
rect 11900 8200 12070 8256
rect 12126 8200 12131 8256
rect 11900 8198 12131 8200
rect 11900 8196 11906 8198
rect 12065 8195 12131 8198
rect 12206 8256 12683 8258
rect 12206 8200 12622 8256
rect 12678 8200 12683 8256
rect 12206 8198 12683 8200
rect 14276 8258 14336 8334
rect 14549 8332 14596 8334
rect 14660 8332 14666 8396
rect 15510 8332 15516 8396
rect 15580 8394 15586 8396
rect 15702 8394 15762 8467
rect 15580 8334 15762 8394
rect 16297 8394 16363 8397
rect 16614 8394 16620 8396
rect 16297 8392 16620 8394
rect 16297 8336 16302 8392
rect 16358 8336 16620 8392
rect 16297 8334 16620 8336
rect 15580 8332 15586 8334
rect 14549 8331 14615 8332
rect 16297 8331 16363 8334
rect 16614 8332 16620 8334
rect 16684 8332 16690 8396
rect 15285 8258 15351 8261
rect 14276 8256 15351 8258
rect 14276 8200 15290 8256
rect 15346 8200 15351 8256
rect 14276 8198 15351 8200
rect 12014 8060 12020 8124
rect 12084 8122 12090 8124
rect 12206 8122 12266 8198
rect 12617 8195 12683 8198
rect 15285 8195 15351 8198
rect 17401 8258 17467 8261
rect 19520 8258 20000 8288
rect 17401 8256 20000 8258
rect 17401 8200 17406 8256
rect 17462 8200 20000 8256
rect 17401 8198 20000 8200
rect 17401 8195 17467 8198
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 19520 8168 20000 8198
rect 12805 8127 13125 8128
rect 12084 8062 12266 8122
rect 12084 8060 12090 8062
rect 14089 7986 14155 7989
rect 9814 7984 14155 7986
rect 9814 7928 14094 7984
rect 14150 7928 14155 7984
rect 9814 7926 14155 7928
rect 3601 7923 3667 7926
rect 8477 7923 8543 7926
rect 14089 7923 14155 7926
rect 3417 7850 3483 7853
rect 8385 7850 8451 7853
rect 3417 7848 8451 7850
rect 3417 7792 3422 7848
rect 3478 7792 8390 7848
rect 8446 7792 8451 7848
rect 3417 7790 8451 7792
rect 3417 7787 3483 7790
rect 8385 7787 8451 7790
rect 10041 7850 10107 7853
rect 10777 7850 10843 7853
rect 13077 7850 13143 7853
rect 10041 7848 10426 7850
rect 10041 7792 10046 7848
rect 10102 7792 10426 7848
rect 10041 7790 10426 7792
rect 10041 7787 10107 7790
rect 10366 7714 10426 7790
rect 10777 7848 13143 7850
rect 10777 7792 10782 7848
rect 10838 7792 13082 7848
rect 13138 7792 13143 7848
rect 10777 7790 13143 7792
rect 10777 7787 10843 7790
rect 13077 7787 13143 7790
rect 17493 7850 17559 7853
rect 19520 7850 20000 7880
rect 17493 7848 20000 7850
rect 17493 7792 17498 7848
rect 17554 7792 20000 7848
rect 17493 7790 20000 7792
rect 17493 7787 17559 7790
rect 19520 7760 20000 7790
rect 13537 7714 13603 7717
rect 10366 7712 13603 7714
rect 10366 7656 13542 7712
rect 13598 7656 13603 7712
rect 10366 7654 13603 7656
rect 13537 7651 13603 7654
rect 3909 7648 4229 7649
rect 0 7578 480 7608
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 6177 7578 6243 7581
rect 0 7518 3802 7578
rect 0 7488 480 7518
rect 3742 7442 3802 7518
rect 4294 7576 6243 7578
rect 4294 7520 6182 7576
rect 6238 7520 6243 7576
rect 4294 7518 6243 7520
rect 4294 7442 4354 7518
rect 6177 7515 6243 7518
rect 11646 7516 11652 7580
rect 11716 7578 11722 7580
rect 11716 7518 13968 7578
rect 11716 7516 11722 7518
rect 13908 7445 13968 7518
rect 3742 7382 4354 7442
rect 13302 7380 13308 7444
rect 13372 7442 13378 7444
rect 13537 7442 13603 7445
rect 13372 7440 13603 7442
rect 13372 7384 13542 7440
rect 13598 7384 13603 7440
rect 13372 7382 13603 7384
rect 13372 7380 13378 7382
rect 13537 7379 13603 7382
rect 13905 7440 13971 7445
rect 13905 7384 13910 7440
rect 13966 7384 13971 7440
rect 13905 7379 13971 7384
rect 16573 7442 16639 7445
rect 19520 7442 20000 7472
rect 16573 7440 20000 7442
rect 16573 7384 16578 7440
rect 16634 7384 20000 7440
rect 16573 7382 20000 7384
rect 16573 7379 16639 7382
rect 19520 7352 20000 7382
rect 12985 7306 13051 7309
rect 13302 7306 13308 7308
rect 12985 7304 13308 7306
rect 12985 7248 12990 7304
rect 13046 7248 13308 7304
rect 12985 7246 13308 7248
rect 12985 7243 13051 7246
rect 13302 7244 13308 7246
rect 13372 7306 13378 7308
rect 15142 7306 15148 7308
rect 13372 7246 15148 7306
rect 13372 7244 13378 7246
rect 15142 7244 15148 7246
rect 15212 7244 15218 7308
rect 0 7170 480 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 480 7110
rect 4061 7107 4127 7110
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 17401 7034 17467 7037
rect 13494 7032 17467 7034
rect 13494 6976 17406 7032
rect 17462 6976 17467 7032
rect 13494 6974 17467 6976
rect 8385 6898 8451 6901
rect 8845 6898 8911 6901
rect 8385 6896 8911 6898
rect 8385 6840 8390 6896
rect 8446 6840 8850 6896
rect 8906 6840 8911 6896
rect 8385 6838 8911 6840
rect 8385 6835 8451 6838
rect 8845 6835 8911 6838
rect 12566 6836 12572 6900
rect 12636 6898 12642 6900
rect 13077 6898 13143 6901
rect 12636 6896 13143 6898
rect 12636 6840 13082 6896
rect 13138 6840 13143 6896
rect 12636 6838 13143 6840
rect 12636 6836 12642 6838
rect 13077 6835 13143 6838
rect 0 6762 480 6792
rect 2773 6762 2839 6765
rect 0 6760 2839 6762
rect 0 6704 2778 6760
rect 2834 6704 2839 6760
rect 0 6702 2839 6704
rect 0 6672 480 6702
rect 2773 6699 2839 6702
rect 3877 6762 3943 6765
rect 6729 6762 6795 6765
rect 12433 6764 12499 6765
rect 3877 6760 6562 6762
rect 3877 6704 3882 6760
rect 3938 6704 6562 6760
rect 3877 6702 6562 6704
rect 3877 6699 3943 6702
rect 6502 6626 6562 6702
rect 6729 6760 12312 6762
rect 6729 6704 6734 6760
rect 6790 6704 12312 6760
rect 6729 6702 12312 6704
rect 6729 6699 6795 6702
rect 8569 6626 8635 6629
rect 6502 6624 8635 6626
rect 6502 6568 8574 6624
rect 8630 6568 8635 6624
rect 6502 6566 8635 6568
rect 12252 6626 12312 6702
rect 12382 6700 12388 6764
rect 12452 6762 12499 6764
rect 12452 6760 12544 6762
rect 12494 6704 12544 6760
rect 12452 6702 12544 6704
rect 12452 6700 12499 6702
rect 12433 6699 12499 6700
rect 13494 6626 13554 6974
rect 17401 6971 17467 6974
rect 18045 7034 18111 7037
rect 19520 7034 20000 7064
rect 18045 7032 20000 7034
rect 18045 6976 18050 7032
rect 18106 6976 20000 7032
rect 18045 6974 20000 6976
rect 18045 6971 18111 6974
rect 19520 6944 20000 6974
rect 13629 6898 13695 6901
rect 13854 6898 13860 6900
rect 13629 6896 13860 6898
rect 13629 6840 13634 6896
rect 13690 6840 13860 6896
rect 13629 6838 13860 6840
rect 13629 6835 13695 6838
rect 13854 6836 13860 6838
rect 13924 6836 13930 6900
rect 15469 6898 15535 6901
rect 15469 6896 15578 6898
rect 15469 6840 15474 6896
rect 15530 6840 15578 6896
rect 15469 6835 15578 6840
rect 12252 6566 13554 6626
rect 8569 6563 8635 6566
rect 3909 6560 4229 6561
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 10501 6490 10567 6493
rect 14038 6490 14044 6492
rect 10501 6488 14044 6490
rect 10501 6432 10506 6488
rect 10562 6432 14044 6488
rect 10501 6430 14044 6432
rect 10501 6427 10567 6430
rect 14038 6428 14044 6430
rect 14108 6428 14114 6492
rect 0 6354 480 6384
rect 3601 6354 3667 6357
rect 0 6352 3667 6354
rect 0 6296 3606 6352
rect 3662 6296 3667 6352
rect 0 6294 3667 6296
rect 0 6264 480 6294
rect 3601 6291 3667 6294
rect 10685 6354 10751 6357
rect 15518 6354 15578 6835
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 6495 16090 6496
rect 17677 6490 17743 6493
rect 19520 6490 20000 6520
rect 17677 6488 20000 6490
rect 17677 6432 17682 6488
rect 17738 6432 20000 6488
rect 17677 6430 20000 6432
rect 17677 6427 17743 6430
rect 19520 6400 20000 6430
rect 15653 6354 15719 6357
rect 10685 6352 15394 6354
rect 10685 6296 10690 6352
rect 10746 6296 15394 6352
rect 10685 6294 15394 6296
rect 15518 6352 15719 6354
rect 15518 6296 15658 6352
rect 15714 6296 15719 6352
rect 15518 6294 15719 6296
rect 10685 6291 10751 6294
rect 3049 6218 3115 6221
rect 9305 6218 9371 6221
rect 3049 6216 9371 6218
rect 3049 6160 3054 6216
rect 3110 6160 9310 6216
rect 9366 6160 9371 6216
rect 3049 6158 9371 6160
rect 15334 6218 15394 6294
rect 15653 6291 15719 6294
rect 17493 6218 17559 6221
rect 15334 6216 17559 6218
rect 15334 6160 17498 6216
rect 17554 6160 17559 6216
rect 15334 6158 17559 6160
rect 3049 6155 3115 6158
rect 9305 6155 9371 6158
rect 17493 6155 17559 6158
rect 18229 6082 18295 6085
rect 19520 6082 20000 6112
rect 18229 6080 20000 6082
rect 18229 6024 18234 6080
rect 18290 6024 20000 6080
rect 18229 6022 20000 6024
rect 18229 6019 18295 6022
rect 6874 6016 7194 6017
rect 0 5946 480 5976
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 19520 5992 20000 6022
rect 12805 5951 13125 5952
rect 1853 5946 1919 5949
rect 17677 5948 17743 5949
rect 17677 5946 17724 5948
rect 0 5944 1919 5946
rect 0 5888 1858 5944
rect 1914 5888 1919 5944
rect 0 5886 1919 5888
rect 17632 5944 17724 5946
rect 17632 5888 17682 5944
rect 17632 5886 17724 5888
rect 0 5856 480 5886
rect 1853 5883 1919 5886
rect 17677 5884 17724 5886
rect 17788 5884 17794 5948
rect 17677 5883 17743 5884
rect 2589 5810 2655 5813
rect 4613 5810 4679 5813
rect 5993 5810 6059 5813
rect 2589 5808 6059 5810
rect 2589 5752 2594 5808
rect 2650 5752 4618 5808
rect 4674 5752 5998 5808
rect 6054 5752 6059 5808
rect 2589 5750 6059 5752
rect 2589 5747 2655 5750
rect 4613 5747 4679 5750
rect 5993 5747 6059 5750
rect 12157 5810 12223 5813
rect 12157 5808 16498 5810
rect 12157 5752 12162 5808
rect 12218 5752 16498 5808
rect 12157 5750 16498 5752
rect 12157 5747 12223 5750
rect 2405 5674 2471 5677
rect 8017 5674 8083 5677
rect 14733 5676 14799 5677
rect 16438 5676 16498 5750
rect 14733 5674 14780 5676
rect 2405 5672 8083 5674
rect 2405 5616 2410 5672
rect 2466 5616 8022 5672
rect 8078 5616 8083 5672
rect 2405 5614 8083 5616
rect 14688 5672 14780 5674
rect 14688 5616 14738 5672
rect 14688 5614 14780 5616
rect 2405 5611 2471 5614
rect 8017 5611 8083 5614
rect 14733 5612 14780 5614
rect 14844 5612 14850 5676
rect 16430 5612 16436 5676
rect 16500 5674 16506 5676
rect 17309 5674 17375 5677
rect 16500 5672 17375 5674
rect 16500 5616 17314 5672
rect 17370 5616 17375 5672
rect 16500 5614 17375 5616
rect 16500 5612 16506 5614
rect 14733 5611 14799 5612
rect 17309 5611 17375 5614
rect 18965 5674 19031 5677
rect 19520 5674 20000 5704
rect 18965 5672 20000 5674
rect 18965 5616 18970 5672
rect 19026 5616 20000 5672
rect 18965 5614 20000 5616
rect 18965 5611 19031 5614
rect 19520 5584 20000 5614
rect 0 5538 480 5568
rect 1853 5538 1919 5541
rect 0 5536 1919 5538
rect 0 5480 1858 5536
rect 1914 5480 1919 5536
rect 0 5478 1919 5480
rect 0 5448 480 5478
rect 1853 5475 1919 5478
rect 14958 5476 14964 5540
rect 15028 5538 15034 5540
rect 15101 5538 15167 5541
rect 15028 5536 15167 5538
rect 15028 5480 15106 5536
rect 15162 5480 15167 5536
rect 15028 5478 15167 5480
rect 15028 5476 15034 5478
rect 15101 5475 15167 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 16297 5402 16363 5405
rect 16297 5400 16498 5402
rect 16297 5344 16302 5400
rect 16358 5344 16498 5400
rect 16297 5342 16498 5344
rect 16297 5339 16363 5342
rect 0 5130 480 5160
rect 16438 5133 16498 5342
rect 18137 5266 18203 5269
rect 19520 5266 20000 5296
rect 18137 5264 20000 5266
rect 18137 5208 18142 5264
rect 18198 5208 20000 5264
rect 18137 5206 20000 5208
rect 18137 5203 18203 5206
rect 19520 5176 20000 5206
rect 1853 5130 1919 5133
rect 0 5128 1919 5130
rect 0 5072 1858 5128
rect 1914 5072 1919 5128
rect 0 5070 1919 5072
rect 16438 5128 16547 5133
rect 16438 5072 16486 5128
rect 16542 5072 16547 5128
rect 16438 5070 16547 5072
rect 0 5040 480 5070
rect 1853 5067 1919 5070
rect 16481 5067 16547 5070
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 9213 4858 9279 4861
rect 11830 4858 11836 4860
rect 9213 4856 11836 4858
rect 9213 4800 9218 4856
rect 9274 4800 11836 4856
rect 9213 4798 11836 4800
rect 9213 4795 9279 4798
rect 11830 4796 11836 4798
rect 11900 4858 11906 4860
rect 12065 4858 12131 4861
rect 11900 4856 12131 4858
rect 11900 4800 12070 4856
rect 12126 4800 12131 4856
rect 11900 4798 12131 4800
rect 11900 4796 11906 4798
rect 12065 4795 12131 4798
rect 13813 4858 13879 4861
rect 14038 4858 14044 4860
rect 13813 4856 14044 4858
rect 13813 4800 13818 4856
rect 13874 4800 14044 4856
rect 13813 4798 14044 4800
rect 13813 4795 13879 4798
rect 14038 4796 14044 4798
rect 14108 4796 14114 4860
rect 17401 4858 17467 4861
rect 19520 4858 20000 4888
rect 17401 4856 20000 4858
rect 17401 4800 17406 4856
rect 17462 4800 20000 4856
rect 17401 4798 20000 4800
rect 17401 4795 17467 4798
rect 19520 4768 20000 4798
rect 0 4722 480 4752
rect 2773 4722 2839 4725
rect 0 4720 2839 4722
rect 0 4664 2778 4720
rect 2834 4664 2839 4720
rect 0 4662 2839 4664
rect 0 4632 480 4662
rect 2773 4659 2839 4662
rect 11145 4722 11211 4725
rect 14222 4722 14228 4724
rect 11145 4720 14228 4722
rect 11145 4664 11150 4720
rect 11206 4664 14228 4720
rect 11145 4662 14228 4664
rect 11145 4659 11211 4662
rect 14222 4660 14228 4662
rect 14292 4660 14298 4724
rect 16798 4660 16804 4724
rect 16868 4722 16874 4724
rect 17125 4722 17191 4725
rect 16868 4720 17191 4722
rect 16868 4664 17130 4720
rect 17186 4664 17191 4720
rect 16868 4662 17191 4664
rect 16868 4660 16874 4662
rect 17125 4659 17191 4662
rect 17861 4450 17927 4453
rect 19520 4450 20000 4480
rect 17861 4448 20000 4450
rect 17861 4392 17866 4448
rect 17922 4392 20000 4448
rect 17861 4390 20000 4392
rect 17861 4387 17927 4390
rect 3909 4384 4229 4385
rect 0 4314 480 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19520 4360 20000 4390
rect 15770 4319 16090 4320
rect 1853 4314 1919 4317
rect 13813 4314 13879 4317
rect 0 4312 1919 4314
rect 0 4256 1858 4312
rect 1914 4256 1919 4312
rect 0 4254 1919 4256
rect 0 4224 480 4254
rect 1853 4251 1919 4254
rect 12022 4312 13879 4314
rect 12022 4256 13818 4312
rect 13874 4256 13879 4312
rect 12022 4254 13879 4256
rect 5349 4180 5415 4181
rect 5349 4178 5396 4180
rect 5304 4176 5396 4178
rect 5304 4120 5354 4176
rect 5304 4118 5396 4120
rect 5349 4116 5396 4118
rect 5460 4116 5466 4180
rect 9305 4178 9371 4181
rect 12022 4178 12082 4254
rect 13813 4251 13879 4254
rect 13302 4178 13308 4180
rect 9305 4176 12082 4178
rect 9305 4120 9310 4176
rect 9366 4120 12082 4176
rect 9305 4118 12082 4120
rect 13126 4118 13308 4178
rect 5349 4115 5415 4116
rect 9305 4115 9371 4118
rect 2129 4042 2195 4045
rect 13126 4042 13186 4118
rect 13302 4116 13308 4118
rect 13372 4116 13378 4180
rect 13721 4178 13787 4181
rect 15929 4178 15995 4181
rect 13721 4176 15995 4178
rect 13721 4120 13726 4176
rect 13782 4120 15934 4176
rect 15990 4120 15995 4176
rect 13721 4118 15995 4120
rect 13721 4115 13787 4118
rect 15929 4115 15995 4118
rect 2129 4040 13186 4042
rect 2129 3984 2134 4040
rect 2190 3984 13186 4040
rect 2129 3982 13186 3984
rect 13353 4042 13419 4045
rect 13721 4044 13787 4045
rect 13486 4042 13492 4044
rect 13353 4040 13492 4042
rect 13353 3984 13358 4040
rect 13414 3984 13492 4040
rect 13353 3982 13492 3984
rect 2129 3979 2195 3982
rect 13353 3979 13419 3982
rect 13486 3980 13492 3982
rect 13556 3980 13562 4044
rect 13670 4042 13676 4044
rect 13630 3982 13676 4042
rect 13740 4040 13787 4044
rect 13782 3984 13787 4040
rect 13670 3980 13676 3982
rect 13740 3980 13787 3984
rect 13721 3979 13787 3980
rect 14549 4044 14615 4045
rect 14549 4040 14596 4044
rect 14660 4042 14666 4044
rect 17677 4042 17743 4045
rect 19520 4042 20000 4072
rect 14549 3984 14554 4040
rect 14549 3980 14596 3984
rect 14660 3982 14706 4042
rect 17677 4040 20000 4042
rect 17677 3984 17682 4040
rect 17738 3984 20000 4040
rect 17677 3982 20000 3984
rect 14660 3980 14666 3982
rect 14549 3979 14615 3980
rect 17677 3979 17743 3982
rect 19520 3952 20000 3982
rect 0 3906 480 3936
rect 2773 3906 2839 3909
rect 0 3904 2839 3906
rect 0 3848 2778 3904
rect 2834 3848 2839 3904
rect 0 3846 2839 3848
rect 0 3816 480 3846
rect 2773 3843 2839 3846
rect 14222 3844 14228 3908
rect 14292 3906 14298 3908
rect 15929 3906 15995 3909
rect 14292 3904 15995 3906
rect 14292 3848 15934 3904
rect 15990 3848 15995 3904
rect 14292 3846 15995 3848
rect 14292 3844 14298 3846
rect 15929 3843 15995 3846
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 15510 3708 15516 3772
rect 15580 3770 15586 3772
rect 15837 3770 15903 3773
rect 15580 3768 15903 3770
rect 15580 3712 15842 3768
rect 15898 3712 15903 3768
rect 15580 3710 15903 3712
rect 15580 3708 15586 3710
rect 15837 3707 15903 3710
rect 3785 3634 3851 3637
rect 8109 3634 8175 3637
rect 3785 3632 8175 3634
rect 3785 3576 3790 3632
rect 3846 3576 8114 3632
rect 8170 3576 8175 3632
rect 3785 3574 8175 3576
rect 3785 3571 3851 3574
rect 8109 3571 8175 3574
rect 15193 3634 15259 3637
rect 19520 3634 20000 3664
rect 15193 3632 20000 3634
rect 15193 3576 15198 3632
rect 15254 3576 20000 3632
rect 15193 3574 20000 3576
rect 15193 3571 15259 3574
rect 19520 3544 20000 3574
rect 0 3498 480 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 480 3438
rect 1853 3435 1919 3438
rect 9949 3498 10015 3501
rect 12198 3498 12204 3500
rect 9949 3496 12204 3498
rect 9949 3440 9954 3496
rect 10010 3440 12204 3496
rect 9949 3438 12204 3440
rect 9949 3435 10015 3438
rect 12198 3436 12204 3438
rect 12268 3498 12274 3500
rect 12341 3498 12407 3501
rect 12268 3496 12407 3498
rect 12268 3440 12346 3496
rect 12402 3440 12407 3496
rect 12268 3438 12407 3440
rect 12268 3436 12274 3438
rect 12341 3435 12407 3438
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 12014 3164 12020 3228
rect 12084 3226 12090 3228
rect 12985 3226 13051 3229
rect 12084 3224 13051 3226
rect 12084 3168 12990 3224
rect 13046 3168 13051 3224
rect 12084 3166 13051 3168
rect 12084 3164 12090 3166
rect 12985 3163 13051 3166
rect 0 3090 480 3120
rect 3325 3090 3391 3093
rect 0 3088 3391 3090
rect 0 3032 3330 3088
rect 3386 3032 3391 3088
rect 0 3030 3391 3032
rect 0 3000 480 3030
rect 3325 3027 3391 3030
rect 11053 3090 11119 3093
rect 15653 3090 15719 3093
rect 19520 3090 20000 3120
rect 11053 3088 13370 3090
rect 11053 3032 11058 3088
rect 11114 3032 13370 3088
rect 11053 3030 13370 3032
rect 11053 3027 11119 3030
rect 12249 2954 12315 2957
rect 13077 2954 13143 2957
rect 12249 2952 13143 2954
rect 12249 2896 12254 2952
rect 12310 2896 13082 2952
rect 13138 2896 13143 2952
rect 12249 2894 13143 2896
rect 13310 2954 13370 3030
rect 15653 3088 20000 3090
rect 15653 3032 15658 3088
rect 15714 3032 20000 3088
rect 15653 3030 20000 3032
rect 15653 3027 15719 3030
rect 19520 3000 20000 3030
rect 15929 2954 15995 2957
rect 16246 2954 16252 2956
rect 13310 2952 16252 2954
rect 13310 2896 15934 2952
rect 15990 2896 16252 2952
rect 13310 2894 16252 2896
rect 12249 2891 12315 2894
rect 13077 2891 13143 2894
rect 15929 2891 15995 2894
rect 16246 2892 16252 2894
rect 16316 2892 16322 2956
rect 6874 2752 7194 2753
rect 0 2682 480 2712
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2687 13125 2688
rect 2773 2682 2839 2685
rect 0 2680 2839 2682
rect 0 2624 2778 2680
rect 2834 2624 2839 2680
rect 0 2622 2839 2624
rect 0 2592 480 2622
rect 2773 2619 2839 2622
rect 14273 2682 14339 2685
rect 14406 2682 14412 2684
rect 14273 2680 14412 2682
rect 14273 2624 14278 2680
rect 14334 2624 14412 2680
rect 14273 2622 14412 2624
rect 14273 2619 14339 2622
rect 14406 2620 14412 2622
rect 14476 2620 14482 2684
rect 15193 2682 15259 2685
rect 19520 2682 20000 2712
rect 15193 2680 20000 2682
rect 15193 2624 15198 2680
rect 15254 2624 20000 2680
rect 15193 2622 20000 2624
rect 15193 2619 15259 2622
rect 19520 2592 20000 2622
rect 0 2274 480 2304
rect 3417 2274 3483 2277
rect 0 2272 3483 2274
rect 0 2216 3422 2272
rect 3478 2216 3483 2272
rect 0 2214 3483 2216
rect 0 2184 480 2214
rect 3417 2211 3483 2214
rect 16297 2274 16363 2277
rect 19520 2274 20000 2304
rect 16297 2272 20000 2274
rect 16297 2216 16302 2272
rect 16358 2216 20000 2272
rect 16297 2214 20000 2216
rect 16297 2211 16363 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 19520 2184 20000 2214
rect 15770 2143 16090 2144
rect 0 1866 480 1896
rect 2957 1866 3023 1869
rect 0 1864 3023 1866
rect 0 1808 2962 1864
rect 3018 1808 3023 1864
rect 0 1806 3023 1808
rect 0 1776 480 1806
rect 2957 1803 3023 1806
rect 11789 1866 11855 1869
rect 19520 1866 20000 1896
rect 11789 1864 20000 1866
rect 11789 1808 11794 1864
rect 11850 1808 20000 1864
rect 11789 1806 20000 1808
rect 11789 1803 11855 1806
rect 19520 1776 20000 1806
rect 0 1458 480 1488
rect 3509 1458 3575 1461
rect 0 1456 3575 1458
rect 0 1400 3514 1456
rect 3570 1400 3575 1456
rect 0 1398 3575 1400
rect 0 1368 480 1398
rect 3509 1395 3575 1398
rect 15285 1458 15351 1461
rect 19520 1458 20000 1488
rect 15285 1456 20000 1458
rect 15285 1400 15290 1456
rect 15346 1400 20000 1456
rect 15285 1398 20000 1400
rect 15285 1395 15351 1398
rect 19520 1368 20000 1398
rect 0 1050 480 1080
rect 3325 1050 3391 1053
rect 0 1048 3391 1050
rect 0 992 3330 1048
rect 3386 992 3391 1048
rect 0 990 3391 992
rect 0 960 480 990
rect 3325 987 3391 990
rect 16389 1050 16455 1053
rect 19520 1050 20000 1080
rect 16389 1048 20000 1050
rect 16389 992 16394 1048
rect 16450 992 20000 1048
rect 16389 990 20000 992
rect 16389 987 16455 990
rect 19520 960 20000 990
rect 0 642 480 672
rect 3233 642 3299 645
rect 0 640 3299 642
rect 0 584 3238 640
rect 3294 584 3299 640
rect 0 582 3299 584
rect 0 552 480 582
rect 3233 579 3299 582
rect 17217 642 17283 645
rect 19520 642 20000 672
rect 17217 640 20000 642
rect 17217 584 17222 640
rect 17278 584 20000 640
rect 17217 582 20000 584
rect 17217 579 17283 582
rect 19520 552 20000 582
rect 0 234 480 264
rect 3049 234 3115 237
rect 0 232 3115 234
rect 0 176 3054 232
rect 3110 176 3115 232
rect 0 174 3115 176
rect 0 144 480 174
rect 3049 171 3115 174
rect 14457 234 14523 237
rect 19520 234 20000 264
rect 14457 232 20000 234
rect 14457 176 14462 232
rect 14518 176 20000 232
rect 14457 174 20000 176
rect 14457 171 14523 174
rect 19520 144 20000 174
<< via3 >>
rect 16436 15404 16500 15468
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 13492 13696 13556 13700
rect 13492 13640 13506 13696
rect 13506 13640 13556 13696
rect 13492 13636 13556 13640
rect 14780 13636 14844 13700
rect 16620 13636 16684 13700
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 17724 13364 17788 13428
rect 13676 13288 13740 13292
rect 13676 13232 13690 13288
rect 13690 13232 13740 13288
rect 13676 13228 13740 13232
rect 14412 13092 14476 13156
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 15148 12412 15212 12476
rect 16252 12276 16316 12340
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 13308 11732 13372 11796
rect 9076 11656 9140 11660
rect 9076 11600 9126 11656
rect 9126 11600 9140 11656
rect 9076 11596 9140 11600
rect 12388 11656 12452 11660
rect 12388 11600 12438 11656
rect 12438 11600 12452 11656
rect 12388 11596 12452 11600
rect 12204 11520 12268 11524
rect 12204 11464 12218 11520
rect 12218 11464 12268 11520
rect 12204 11460 12268 11464
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 14228 11324 14292 11388
rect 8524 11188 8588 11252
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 11652 10780 11716 10844
rect 12572 10644 12636 10708
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 12020 10236 12084 10300
rect 16804 10236 16868 10300
rect 8524 9828 8588 9892
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 9076 9692 9140 9756
rect 13860 9344 13924 9348
rect 13860 9288 13910 9344
rect 13910 9288 13924 9344
rect 13860 9284 13924 9288
rect 15332 9420 15396 9484
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 14044 9208 14108 9212
rect 14044 9152 14058 9208
rect 14058 9152 14108 9208
rect 14044 9148 14108 9152
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 12020 8604 12084 8668
rect 14964 8664 15028 8668
rect 14964 8608 15014 8664
rect 15014 8608 15028 8664
rect 14964 8604 15028 8608
rect 15332 8468 15396 8532
rect 5396 8332 5460 8396
rect 14596 8392 14660 8396
rect 14596 8336 14610 8392
rect 14610 8336 14660 8392
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 11836 8196 11900 8260
rect 14596 8332 14660 8336
rect 15516 8332 15580 8396
rect 16620 8332 16684 8396
rect 12020 8060 12084 8124
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 11652 7516 11716 7580
rect 13308 7380 13372 7444
rect 13308 7244 13372 7308
rect 15148 7244 15212 7308
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 12572 6836 12636 6900
rect 12388 6760 12452 6764
rect 12388 6704 12438 6760
rect 12438 6704 12452 6760
rect 12388 6700 12452 6704
rect 13860 6836 13924 6900
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 14044 6428 14108 6492
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 17724 5944 17788 5948
rect 17724 5888 17738 5944
rect 17738 5888 17788 5944
rect 17724 5884 17788 5888
rect 14780 5672 14844 5676
rect 14780 5616 14794 5672
rect 14794 5616 14844 5672
rect 14780 5612 14844 5616
rect 16436 5612 16500 5676
rect 14964 5476 15028 5540
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 11836 4796 11900 4860
rect 14044 4796 14108 4860
rect 14228 4660 14292 4724
rect 16804 4660 16868 4724
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 5396 4176 5460 4180
rect 5396 4120 5410 4176
rect 5410 4120 5460 4176
rect 5396 4116 5460 4120
rect 13308 4116 13372 4180
rect 13492 3980 13556 4044
rect 13676 4040 13740 4044
rect 13676 3984 13726 4040
rect 13726 3984 13740 4040
rect 13676 3980 13740 3984
rect 14596 4040 14660 4044
rect 14596 3984 14610 4040
rect 14610 3984 14660 4040
rect 14596 3980 14660 3984
rect 14228 3844 14292 3908
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 15516 3708 15580 3772
rect 12204 3436 12268 3500
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 12020 3164 12084 3228
rect 16252 2892 16316 2956
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 14412 2620 14476 2684
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 16435 15468 16501 15469
rect 16435 15404 16436 15468
rect 16500 15404 16501 15468
rect 16435 15403 16501 15404
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9075 11660 9141 11661
rect 9075 11596 9076 11660
rect 9140 11596 9141 11660
rect 9075 11595 9141 11596
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 8523 11252 8589 11253
rect 8523 11188 8524 11252
rect 8588 11188 8589 11252
rect 8523 11187 8589 11188
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 8526 9893 8586 11187
rect 8523 9892 8589 9893
rect 8523 9828 8524 9892
rect 8588 9828 8589 9892
rect 8523 9827 8589 9828
rect 9078 9757 9138 11595
rect 9840 10912 10160 11936
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 15770 14176 16090 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 13491 13700 13557 13701
rect 13491 13636 13492 13700
rect 13556 13636 13557 13700
rect 13491 13635 13557 13636
rect 14779 13700 14845 13701
rect 14779 13636 14780 13700
rect 14844 13636 14845 13700
rect 14779 13635 14845 13636
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12387 11660 12453 11661
rect 12387 11596 12388 11660
rect 12452 11596 12453 11660
rect 12387 11595 12453 11596
rect 12203 11524 12269 11525
rect 12203 11460 12204 11524
rect 12268 11460 12269 11524
rect 12203 11459 12269 11460
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 11651 10844 11717 10845
rect 11651 10780 11652 10844
rect 11716 10780 11717 10844
rect 11651 10779 11717 10780
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9075 9756 9141 9757
rect 9075 9692 9076 9756
rect 9140 9692 9141 9756
rect 9075 9691 9141 9692
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 5395 8396 5461 8397
rect 5395 8332 5396 8396
rect 5460 8332 5461 8396
rect 5395 8331 5461 8332
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 5398 4181 5458 8331
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 5395 4180 5461 4181
rect 5395 4116 5396 4180
rect 5460 4116 5461 4180
rect 5395 4115 5461 4116
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 11654 7581 11714 10779
rect 12019 10300 12085 10301
rect 12019 10236 12020 10300
rect 12084 10236 12085 10300
rect 12019 10235 12085 10236
rect 12022 8669 12082 10235
rect 12019 8668 12085 8669
rect 12019 8604 12020 8668
rect 12084 8604 12085 8668
rect 12019 8603 12085 8604
rect 11835 8260 11901 8261
rect 11835 8196 11836 8260
rect 11900 8196 11901 8260
rect 11835 8195 11901 8196
rect 11651 7580 11717 7581
rect 11651 7516 11652 7580
rect 11716 7516 11717 7580
rect 11651 7515 11717 7516
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 11838 4861 11898 8195
rect 12019 8124 12085 8125
rect 12019 8060 12020 8124
rect 12084 8060 12085 8124
rect 12019 8059 12085 8060
rect 11835 4860 11901 4861
rect 11835 4796 11836 4860
rect 11900 4796 11901 4860
rect 11835 4795 11901 4796
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 12022 3229 12082 8059
rect 12206 3501 12266 11459
rect 12390 6765 12450 11595
rect 12805 11456 13125 12480
rect 13307 11796 13373 11797
rect 13307 11732 13308 11796
rect 13372 11732 13373 11796
rect 13307 11731 13373 11732
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12571 10708 12637 10709
rect 12571 10644 12572 10708
rect 12636 10644 12637 10708
rect 12571 10643 12637 10644
rect 12574 6901 12634 10643
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 13310 7445 13370 11731
rect 13307 7444 13373 7445
rect 13307 7380 13308 7444
rect 13372 7380 13373 7444
rect 13307 7379 13373 7380
rect 13307 7308 13373 7309
rect 13307 7244 13308 7308
rect 13372 7244 13373 7308
rect 13307 7243 13373 7244
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12571 6900 12637 6901
rect 12571 6836 12572 6900
rect 12636 6836 12637 6900
rect 12571 6835 12637 6836
rect 12387 6764 12453 6765
rect 12387 6700 12388 6764
rect 12452 6700 12453 6764
rect 12387 6699 12453 6700
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 3840 13125 4864
rect 13310 4181 13370 7243
rect 13307 4180 13373 4181
rect 13307 4116 13308 4180
rect 13372 4116 13373 4180
rect 13307 4115 13373 4116
rect 13494 4045 13554 13635
rect 13675 13292 13741 13293
rect 13675 13228 13676 13292
rect 13740 13228 13741 13292
rect 13675 13227 13741 13228
rect 13678 4045 13738 13227
rect 14411 13156 14477 13157
rect 14411 13092 14412 13156
rect 14476 13092 14477 13156
rect 14411 13091 14477 13092
rect 14227 11388 14293 11389
rect 14227 11324 14228 11388
rect 14292 11324 14293 11388
rect 14227 11323 14293 11324
rect 13859 9348 13925 9349
rect 13859 9284 13860 9348
rect 13924 9284 13925 9348
rect 13859 9283 13925 9284
rect 13862 6901 13922 9283
rect 14043 9212 14109 9213
rect 14043 9148 14044 9212
rect 14108 9148 14109 9212
rect 14043 9147 14109 9148
rect 13859 6900 13925 6901
rect 13859 6836 13860 6900
rect 13924 6836 13925 6900
rect 13859 6835 13925 6836
rect 14046 6493 14106 9147
rect 14043 6492 14109 6493
rect 14043 6428 14044 6492
rect 14108 6428 14109 6492
rect 14043 6427 14109 6428
rect 14046 4861 14106 6427
rect 14043 4860 14109 4861
rect 14043 4796 14044 4860
rect 14108 4796 14109 4860
rect 14043 4795 14109 4796
rect 14230 4725 14290 11323
rect 14227 4724 14293 4725
rect 14227 4660 14228 4724
rect 14292 4660 14293 4724
rect 14227 4659 14293 4660
rect 13491 4044 13557 4045
rect 13491 3980 13492 4044
rect 13556 3980 13557 4044
rect 13491 3979 13557 3980
rect 13675 4044 13741 4045
rect 13675 3980 13676 4044
rect 13740 3980 13741 4044
rect 13675 3979 13741 3980
rect 14230 3909 14290 4659
rect 14227 3908 14293 3909
rect 14227 3844 14228 3908
rect 14292 3844 14293 3908
rect 14227 3843 14293 3844
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12203 3500 12269 3501
rect 12203 3436 12204 3500
rect 12268 3436 12269 3500
rect 12203 3435 12269 3436
rect 12019 3228 12085 3229
rect 12019 3164 12020 3228
rect 12084 3164 12085 3228
rect 12019 3163 12085 3164
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 14414 2685 14474 13091
rect 14595 8396 14661 8397
rect 14595 8332 14596 8396
rect 14660 8332 14661 8396
rect 14595 8331 14661 8332
rect 14598 4045 14658 8331
rect 14782 5677 14842 13635
rect 15770 13088 16090 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15147 12476 15213 12477
rect 15147 12412 15148 12476
rect 15212 12412 15213 12476
rect 15147 12411 15213 12412
rect 14963 8668 15029 8669
rect 14963 8604 14964 8668
rect 15028 8604 15029 8668
rect 14963 8603 15029 8604
rect 14779 5676 14845 5677
rect 14779 5612 14780 5676
rect 14844 5612 14845 5676
rect 14779 5611 14845 5612
rect 14966 5541 15026 8603
rect 15150 7309 15210 12411
rect 15770 12000 16090 13024
rect 16251 12340 16317 12341
rect 16251 12276 16252 12340
rect 16316 12276 16317 12340
rect 16251 12275 16317 12276
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 10912 16090 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 9824 16090 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15331 9484 15397 9485
rect 15331 9420 15332 9484
rect 15396 9420 15397 9484
rect 15331 9419 15397 9420
rect 15334 8533 15394 9419
rect 15770 8736 16090 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15331 8532 15397 8533
rect 15331 8468 15332 8532
rect 15396 8468 15397 8532
rect 15331 8467 15397 8468
rect 15515 8396 15581 8397
rect 15515 8332 15516 8396
rect 15580 8332 15581 8396
rect 15515 8331 15581 8332
rect 15147 7308 15213 7309
rect 15147 7244 15148 7308
rect 15212 7244 15213 7308
rect 15147 7243 15213 7244
rect 14963 5540 15029 5541
rect 14963 5476 14964 5540
rect 15028 5476 15029 5540
rect 14963 5475 15029 5476
rect 14595 4044 14661 4045
rect 14595 3980 14596 4044
rect 14660 3980 14661 4044
rect 14595 3979 14661 3980
rect 15518 3773 15578 8331
rect 15770 7648 16090 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 6560 16090 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 5472 16090 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 4384 16090 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15515 3772 15581 3773
rect 15515 3708 15516 3772
rect 15580 3708 15581 3772
rect 15515 3707 15581 3708
rect 15770 3296 16090 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 14411 2684 14477 2685
rect 14411 2620 14412 2684
rect 14476 2620 14477 2684
rect 14411 2619 14477 2620
rect 15770 2208 16090 3232
rect 16254 2957 16314 12275
rect 16438 5677 16498 15403
rect 16619 13700 16685 13701
rect 16619 13636 16620 13700
rect 16684 13636 16685 13700
rect 16619 13635 16685 13636
rect 16622 8397 16682 13635
rect 17723 13428 17789 13429
rect 17723 13364 17724 13428
rect 17788 13364 17789 13428
rect 17723 13363 17789 13364
rect 16803 10300 16869 10301
rect 16803 10236 16804 10300
rect 16868 10236 16869 10300
rect 16803 10235 16869 10236
rect 16619 8396 16685 8397
rect 16619 8332 16620 8396
rect 16684 8332 16685 8396
rect 16619 8331 16685 8332
rect 16435 5676 16501 5677
rect 16435 5612 16436 5676
rect 16500 5612 16501 5676
rect 16435 5611 16501 5612
rect 16806 4725 16866 10235
rect 17726 5949 17786 13363
rect 17723 5948 17789 5949
rect 17723 5884 17724 5948
rect 17788 5884 17789 5948
rect 17723 5883 17789 5884
rect 16803 4724 16869 4725
rect 16803 4660 16804 4724
rect 16868 4660 16869 4724
rect 16803 4659 16869 4660
rect 16251 2956 16317 2957
rect 16251 2892 16252 2956
rect 16316 2892 16317 2956
rect 16251 2891 16317 2892
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2128 16090 2144
use sky130_fd_sc_hd__fill_1  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1564 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1472 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11
timestamp 1606256979
transform 1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1606256979
transform 1 0 2944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19
timestamp 1606256979
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2392 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _26_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1606256979
transform 1 0 3220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 4232 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 3312 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1606256979
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4416 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1606256979
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1606256979
transform 1 0 4784 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_49
timestamp 1606256979
transform 1 0 5612 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_44
timestamp 1606256979
transform 1 0 5152 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50
timestamp 1606256979
transform 1 0 5704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44
timestamp 1606256979
transform 1 0 5152 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606256979
transform 1 0 5244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606256979
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1606256979
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58
timestamp 1606256979
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606256979
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606256979
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606256979
transform 1 0 8004 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 8740 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606256979
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1606256979
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1606256979
transform 1 0 7636 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_79
timestamp 1606256979
transform 1 0 8372 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 10304 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 10120 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1606256979
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1606256979
transform 1 0 9936 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1606256979
transform 1 0 11500 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111
timestamp 1606256979
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1606256979
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1606256979
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1606256979
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1606256979
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 12604 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606256979
transform 1 0 13156 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 14168 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144
timestamp 1606256979
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1606256979
transform 1 0 13800 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 14720 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 15732 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1606256979
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_155
timestamp 1606256979
transform 1 0 15364 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1606256979
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1606256979
transform 1 0 16652 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_184
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1606256979
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1606256979
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1606256979
transform 1 0 17388 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606256979
transform 1 0 17296 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606256979
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1606256979
transform 1 0 1656 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1606256979
transform 1 0 2852 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_12
timestamp 1606256979
transform 1 0 2208 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_18
timestamp 1606256979
transform 1 0 2760 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_25
timestamp 1606256979
transform 1 0 3404 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5888 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1606256979
transform 1 0 5520 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _13_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7728 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606256979
transform 1 0 8372 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1606256979
transform 1 0 7360 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1606256979
transform 1 0 8004 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606256979
transform 1 0 10028 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1606256979
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606256979
transform 1 0 11224 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1606256979
transform 1 0 10856 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1606256979
transform 1 0 12420 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1606256979
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606256979
transform 1 0 12788 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_2_140
timestamp 1606256979
transform 1 0 13984 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_144
timestamp 1606256979
transform 1 0 14352 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 15456 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1606256979
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1606256979
transform 1 0 16284 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606256979
transform 1 0 17848 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_2_
timestamp 1606256979
transform 1 0 16652 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_178
timestamp 1606256979
transform 1 0 17480 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1606256979
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1606256979
transform 1 0 1656 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1606256979
transform 1 0 2392 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606256979
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_12
timestamp 1606256979
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 1606256979
transform 1 0 2760 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1606256979
transform 1 0 3128 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3956 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_26
timestamp 1606256979
transform 1 0 3496 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_30
timestamp 1606256979
transform 1 0 3864 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1606256979
transform 1 0 4784 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1606256979
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_78
timestamp 1606256979
transform 1 0 8280 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606256979
transform 1 0 9108 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10304 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_86
timestamp 1606256979
transform 1 0 9016 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1606256979
transform 1 0 9936 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_116
timestamp 1606256979
transform 1 0 11776 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606256979
transform 1 0 12788 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606256979
transform 1 0 14352 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_3_140
timestamp 1606256979
transform 1 0 13984 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 16008 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_3_157
timestamp 1606256979
transform 1 0 15548 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_161
timestamp 1606256979
transform 1 0 15916 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_175
timestamp 1606256979
transform 1 0 17204 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_184
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1606256979
transform 1 0 1656 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1606256979
transform 1 0 2392 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1606256979
transform 1 0 2024 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_18
timestamp 1606256979
transform 1 0 2760 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1606256979
transform 1 0 3128 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4416 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_26
timestamp 1606256979
transform 1 0 3496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1606256979
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 5612 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1606256979
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1606256979
transform 1 0 6440 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_62
timestamp 1606256979
transform 1 0 6808 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1606256979
transform 1 0 6900 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7636 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_67
timestamp 1606256979
transform 1 0 7268 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606256979
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1606256979
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1606256979
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1606256979
transform 1 0 10028 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 11868 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_4_110
timestamp 1606256979
transform 1 0 11224 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_116
timestamp 1606256979
transform 1 0 11776 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 13616 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_4_130
timestamp 1606256979
transform 1 0 13064 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1606256979
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_167
timestamp 1606256979
transform 1 0 16468 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_180
timestamp 1606256979
transform 1 0 17664 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1606256979
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1606256979
transform 1 0 1656 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2576 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_10
timestamp 1606256979
transform 1 0 2024 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4876 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 3680 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_22
timestamp 1606256979
transform 1 0 3128 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1606256979
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1606256979
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8096 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_71
timestamp 1606256979
transform 1 0 7636 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_75
timestamp 1606256979
transform 1 0 8004 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10212 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9936 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_92
timestamp 1606256979
transform 1 0 9568 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1606256979
transform 1 0 12512 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1606256979
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1606256979
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_123
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606256979
transform 1 0 13248 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_5_128
timestamp 1606256979
transform 1 0 12880 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1606256979
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _15_
timestamp 1606256979
transform 1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15456 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_152
timestamp 1606256979
transform 1 0 15088 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_165
timestamp 1606256979
transform 1 0 16284 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1606256979
transform 1 0 16652 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1606256979
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1606256979
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_184
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_10
timestamp 1606256979
transform 1 0 2024 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1656 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1606256979
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_12
timestamp 1606256979
transform 1 0 2208 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2760 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2392 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4600 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_41
timestamp 1606256979
transform 1 0 4876 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_30
timestamp 1606256979
transform 1 0 3864 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606256979
transform 1 0 5520 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6256 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_47
timestamp 1606256979
transform 1 0 5428 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1606256979
transform 1 0 5888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_54
timestamp 1606256979
transform 1 0 6072 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606256979
transform 1 0 8372 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8004 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_6_72
timestamp 1606256979
transform 1 0 7728 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_78
timestamp 1606256979
transform 1 0 8280 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_71
timestamp 1606256979
transform 1 0 7636 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9200 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1606256979
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_84
timestamp 1606256979
transform 1 0 8832 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_104
timestamp 1606256979
transform 1 0 10672 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 11500 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1606256979
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1606256979
transform 1 0 11132 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_108
timestamp 1606256979
transform 1 0 11040 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606256979
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13340 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 14076 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_129
timestamp 1606256979
transform 1 0 12972 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1606256979
transform 1 0 13616 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_140
timestamp 1606256979
transform 1 0 13984 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1606256979
transform 1 0 15364 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1606256979
transform 1 0 16100 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1606256979
transform 1 0 15916 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1606256979
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_154
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_159
timestamp 1606256979
transform 1 0 15732 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_157
timestamp 1606256979
transform 1 0 15548 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606256979
transform 1 0 17204 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1606256979
transform 1 0 17296 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_172
timestamp 1606256979
transform 1 0 16928 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_185
timestamp 1606256979
transform 1 0 18124 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_170
timestamp 1606256979
transform 1 0 16744 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_174
timestamp 1606256979
transform 1 0 17112 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1606256979
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_184
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_189
timestamp 1606256979
transform 1 0 18492 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1606256979
transform 1 0 1656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2760 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_10
timestamp 1606256979
transform 1 0 2024 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 5888 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_48
timestamp 1606256979
transform 1 0 5520 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1606256979
transform 1 0 6716 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 7084 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 8372 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_74
timestamp 1606256979
transform 1 0 7912 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_78
timestamp 1606256979
transform 1 0 8280 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10396 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1606256979
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp 1606256979
transform 1 0 10028 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1606256979
transform 1 0 11592 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_110
timestamp 1606256979
transform 1 0 11224 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_123
timestamp 1606256979
transform 1 0 12420 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12788 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13984 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1606256979
transform 1 0 13616 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1606256979
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_163
timestamp 1606256979
transform 1 0 16100 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606256979
transform 1 0 17848 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16652 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1606256979
transform 1 0 17480 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1606256979
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1606256979
transform 1 0 1472 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2208 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1606256979
transform 1 0 1840 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1606256979
transform 1 0 3404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4324 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_21
timestamp 1606256979
transform 1 0 3036 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_29
timestamp 1606256979
transform 1 0 3772 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5520 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_44
timestamp 1606256979
transform 1 0 5152 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1606256979
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8372 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1606256979
transform 1 0 7176 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_75
timestamp 1606256979
transform 1 0 8004 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10304 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1606256979
transform 1 0 9844 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 1606256979
transform 1 0 10212 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_116
timestamp 1606256979
transform 1 0 11776 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 13708 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1606256979
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_136
timestamp 1606256979
transform 1 0 13616 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15548 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1606256979
transform 1 0 15180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_173
timestamp 1606256979
transform 1 0 17020 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1606256979
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_184
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1606256979
transform 1 0 2668 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1472 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1606256979
transform 1 0 2300 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4508 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_26
timestamp 1606256979
transform 1 0 3496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1606256979
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1606256979
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5704 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1606256979
transform 1 0 5336 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1606256979
transform 1 0 8740 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1606256979
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_66
timestamp 1606256979
transform 1 0 7176 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1606256979
transform 1 0 8372 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1606256979
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1606256979
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11684 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_109
timestamp 1606256979
transform 1 0 11132 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1606256979
transform 1 0 12512 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606256979
transform 1 0 14444 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12880 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_137
timestamp 1606256979
transform 1 0 13708 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15732 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1606256979
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1606256979
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1606256979
transform 1 0 16928 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_168
timestamp 1606256979
transform 1 0 16560 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_181
timestamp 1606256979
transform 1 0 17756 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1606256979
transform 1 0 18492 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1606256979
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_17
timestamp 1606256979
transform 1 0 2668 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 4232 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1606256979
transform 1 0 3036 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1606256979
transform 1 0 3864 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5520 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_43
timestamp 1606256979
transform 1 0 5060 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_47
timestamp 1606256979
transform 1 0 5428 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1606256979
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7360 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 8556 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1606256979
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1606256979
transform 1 0 8188 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10396 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1606256979
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1606256979
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12880 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_127
timestamp 1606256979
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_137
timestamp 1606256979
transform 1 0 13708 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_145
timestamp 1606256979
transform 1 0 14444 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 14536 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_162
timestamp 1606256979
transform 1 0 16008 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_175
timestamp 1606256979
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1564 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_21
timestamp 1606256979
transform 1 0 3036 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1606256979
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5888 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_48
timestamp 1606256979
transform 1 0 5520 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 1606256979
transform 1 0 6716 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 8372 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_74
timestamp 1606256979
transform 1 0 7912 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_78
timestamp 1606256979
transform 1 0 8280 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1606256979
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1606256979
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10948 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1606256979
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_123
timestamp 1606256979
transform 1 0 12420 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606256979
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12880 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 14076 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_127
timestamp 1606256979
transform 1 0 12788 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_137
timestamp 1606256979
transform 1 0 13708 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_144
timestamp 1606256979
transform 1 0 14352 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1606256979
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1606256979
transform 1 0 17112 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1606256979
transform 1 0 16744 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_183
timestamp 1606256979
transform 1 0 17940 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1606256979
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1840 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 2760 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1606256979
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1606256979
transform 1 0 2392 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_24
timestamp 1606256979
transform 1 0 3312 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_37
timestamp 1606256979
transform 1 0 4508 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606256979
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_38
timestamp 1606256979
transform 1 0 4600 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_51
timestamp 1606256979
transform 1 0 5796 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_43
timestamp 1606256979
transform 1 0 5060 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 5152 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4968 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5428 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1606256979
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_56
timestamp 1606256979
transform 1 0 6256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1606256979
transform 1 0 6164 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7544 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6992 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_80
timestamp 1606256979
transform 1 0 8464 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_64
timestamp 1606256979
transform 1 0 6992 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_86
timestamp 1606256979
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_93
timestamp 1606256979
transform 1 0 9660 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8832 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_103
timestamp 1606256979
transform 1 0 10580 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_103
timestamp 1606256979
transform 1 0 10580 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1606256979
transform 1 0 9752 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9752 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10672 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12144 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1606256979
transform 1 0 10948 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1606256979
transform 1 0 11500 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1606256979
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_116
timestamp 1606256979
transform 1 0 11776 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _14_
timestamp 1606256979
transform 1 0 13616 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 14260 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13340 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1606256979
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_139
timestamp 1606256979
transform 1 0 13892 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_129
timestamp 1606256979
transform 1 0 12972 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_142
timestamp 1606256979
transform 1 0 14168 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1606256979
transform 1 0 16100 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606256979
transform 1 0 14536 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15824 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_159
timestamp 1606256979
transform 1 0 15732 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_166
timestamp 1606256979
transform 1 0 16376 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1606256979
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_154
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1606256979
transform 1 0 16744 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1606256979
transform 1 0 17204 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1606256979
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_184
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_169
timestamp 1606256979
transform 1 0 16652 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_184
timestamp 1606256979
transform 1 0 18032 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1606256979
transform 1 0 1656 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2392 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_10
timestamp 1606256979
transform 1 0 2024 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4600 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 4324 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1606256979
transform 1 0 3864 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_34
timestamp 1606256979
transform 1 0 4232 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1606256979
transform 1 0 5428 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1606256979
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606256979
transform 1 0 8004 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1606256979
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_79
timestamp 1606256979
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_83
timestamp 1606256979
transform 1 0 8740 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 8832 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1606256979
transform 1 0 10672 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_100
timestamp 1606256979
transform 1 0 10304 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1606256979
transform 1 0 11500 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1606256979
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606256979
transform 1 0 12788 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13524 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_131
timestamp 1606256979
transform 1 0 13156 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15364 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_151
timestamp 1606256979
transform 1 0 14996 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606256979
transform 1 0 17204 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_171
timestamp 1606256979
transform 1 0 16836 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1606256979
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_184
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1606256979
transform 1 0 2668 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1472 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1606256979
transform 1 0 2300 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_26
timestamp 1606256979
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1606256979
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 1606256979
transform 1 0 4876 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606256979
transform 1 0 6716 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1606256979
transform 1 0 5336 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_45
timestamp 1606256979
transform 1 0 5244 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_55
timestamp 1606256979
transform 1 0 6164 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7452 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_65
timestamp 1606256979
transform 1 0 7084 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _09_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10488 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1606256979
transform 1 0 8924 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1606256979
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_96
timestamp 1606256979
transform 1 0 9936 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12512 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_16_118
timestamp 1606256979
transform 1 0 11960 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606256979
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_140
timestamp 1606256979
transform 1 0 13984 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_144
timestamp 1606256979
transform 1 0 14352 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1606256979
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1606256979
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606256979
transform 1 0 17848 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1606256979
transform 1 0 16468 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_176
timestamp 1606256979
transform 1 0 17296 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_186
timestamp 1606256979
transform 1 0 18216 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1606256979
transform 1 0 1564 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 2300 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1606256979
transform 1 0 1932 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 3588 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_22
timestamp 1606256979
transform 1 0 3128 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_26
timestamp 1606256979
transform 1 0 3496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5428 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_43
timestamp 1606256979
transform 1 0 5060 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_56
timestamp 1606256979
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1606256979
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8648 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1606256979
transform 1 0 8280 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_91 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9476 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_103
timestamp 1606256979
transform 1 0 10580 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_115
timestamp 1606256979
transform 1 0 11684 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1606256979
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13616 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1606256979
transform 1 0 13248 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_145
timestamp 1606256979
transform 1 0 14444 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606256979
transform 1 0 15732 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606256979
transform 1 0 14996 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_155
timestamp 1606256979
transform 1 0 15364 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1606256979
transform 1 0 16100 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1606256979
transform 1 0 17204 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606256979
transform 1 0 16468 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_171
timestamp 1606256979
transform 1 0 16836 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1606256979
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1606256979
transform 1 0 1564 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2300 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_9
timestamp 1606256979
transform 1 0 1932 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4600 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_22
timestamp 1606256979
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1606256979
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_32
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6440 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1606256979
transform 1 0 6072 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1606256979
transform 1 0 8280 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1606256979
transform 1 0 7912 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1606256979
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1606256979
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606256979
transform 1 0 12420 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1606256979
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_117
timestamp 1606256979
transform 1 0 11868 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606256979
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606256979
transform 1 0 13340 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_126
timestamp 1606256979
transform 1 0 12696 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_132
timestamp 1606256979
transform 1 0 13248 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_136
timestamp 1606256979
transform 1 0 13616 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_144
timestamp 1606256979
transform 1 0 14352 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606256979
transform 1 0 16376 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606256979
transform 1 0 15640 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1606256979
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_162
timestamp 1606256979
transform 1 0 16008 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1606256979
transform 1 0 17112 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606256979
transform 1 0 17848 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_170
timestamp 1606256979
transform 1 0 16744 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_178
timestamp 1606256979
transform 1 0 17480 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1606256979
transform 1 0 18216 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_9
timestamp 1606256979
transform 1 0 1932 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606256979
transform 1 0 1564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_14
timestamp 1606256979
transform 1 0 2392 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1606256979
transform 1 0 2300 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2760 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _10_
timestamp 1606256979
transform 1 0 4600 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_34
timestamp 1606256979
transform 1 0 4232 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_41
timestamp 1606256979
transform 1 0 4876 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_22
timestamp 1606256979
transform 1 0 3128 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1606256979
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_35
timestamp 1606256979
transform 1 0 4324 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _12_
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1606256979
transform 1 0 5520 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606256979
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_45
timestamp 1606256979
transform 1 0 5244 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1606256979
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_47
timestamp 1606256979
transform 1 0 5428 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_59
timestamp 1606256979
transform 1 0 6532 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7728 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_65
timestamp 1606256979
transform 1 0 7084 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_71
timestamp 1606256979
transform 1 0 7636 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_71
timestamp 1606256979
transform 1 0 7636 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_83
timestamp 1606256979
transform 1 0 8740 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_84
timestamp 1606256979
transform 1 0 8832 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_96
timestamp 1606256979
transform 1 0 9936 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606256979
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_108
timestamp 1606256979
transform 1 0 11040 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1606256979
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1606256979
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1606256979
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606256979
transform 1 0 12788 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606256979
transform 1 0 14168 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_130
timestamp 1606256979
transform 1 0 13064 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1606256979
transform 1 0 14444 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1606256979
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1606256979
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606256979
transform 1 0 15548 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606256979
transform 1 0 14904 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606256979
transform 1 0 15364 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_149
timestamp 1606256979
transform 1 0 14812 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1606256979
transform 1 0 15180 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1606256979
transform 1 0 15916 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_154
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_158
timestamp 1606256979
transform 1 0 15640 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606256979
transform 1 0 17848 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606256979
transform 1 0 17204 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606256979
transform 1 0 16468 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_171
timestamp 1606256979
transform 1 0 16836 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1606256979
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_170
timestamp 1606256979
transform 1 0 16744 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1606256979
transform 1 0 18216 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606256979
transform 1 0 1840 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1606256979
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_12
timestamp 1606256979
transform 1 0 2208 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_20
timestamp 1606256979
transform 1 0 2944 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1606256979
transform 1 0 3036 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_25
timestamp 1606256979
transform 1 0 3404 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_37
timestamp 1606256979
transform 1 0 4508 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1606256979
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_49
timestamp 1606256979
transform 1 0 5612 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1606256979
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_66
timestamp 1606256979
transform 1 0 7176 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_78
timestamp 1606256979
transform 1 0 8280 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_90
timestamp 1606256979
transform 1 0 9384 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_102
timestamp 1606256979
transform 1 0 10488 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1606256979
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606256979
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606256979
transform 1 0 14444 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1606256979
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1606256979
transform 1 0 13984 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_144
timestamp 1606256979
transform 1 0 14352 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606256979
transform 1 0 15640 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1606256979
transform 1 0 14812 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_157
timestamp 1606256979
transform 1 0 15548 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_162
timestamp 1606256979
transform 1 0 16008 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_174
timestamp 1606256979
transform 1 0 17112 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1606256979
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_184
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606256979
transform 1 0 1656 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606256979
transform 1 0 2484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_10
timestamp 1606256979
transform 1 0 2024 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_14
timestamp 1606256979
transform 1 0 2392 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_19
timestamp 1606256979
transform 1 0 2852 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1606256979
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1606256979
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1606256979
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1606256979
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1606256979
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1606256979
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1606256979
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1606256979
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1606256979
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1606256979
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606256979
transform 1 0 15456 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1606256979
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_160
timestamp 1606256979
transform 1 0 15824 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_172
timestamp 1606256979
transform 1 0 16928 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_184
timestamp 1606256979
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1606256979
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 7378 16520 7434 17000 6 IO_ISOL_N
port 0 nsew default input
rlabel metal2 s 5630 0 5686 480 6 SC_IN_BOT
port 1 nsew default input
rlabel metal2 s 6090 16520 6146 17000 6 SC_IN_TOP
port 2 nsew default input
rlabel metal2 s 6182 0 6238 480 6 SC_OUT_BOT
port 3 nsew default tristate
rlabel metal2 s 6734 16520 6790 17000 6 SC_OUT_TOP
port 4 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_grid_pin_0_
port 5 nsew default tristate
rlabel metal2 s 2686 0 2742 480 6 bottom_grid_pin_10_
port 6 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 bottom_grid_pin_12_
port 7 nsew default tristate
rlabel metal2 s 3606 0 3662 480 6 bottom_grid_pin_14_
port 8 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 bottom_grid_pin_16_
port 9 nsew default tristate
rlabel metal2 s 662 0 718 480 6 bottom_grid_pin_2_
port 10 nsew default tristate
rlabel metal2 s 1122 0 1178 480 6 bottom_grid_pin_4_
port 11 nsew default tristate
rlabel metal2 s 1674 0 1730 480 6 bottom_grid_pin_6_
port 12 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 bottom_grid_pin_8_
port 13 nsew default tristate
rlabel metal2 s 4618 0 4674 480 6 ccff_head
port 14 nsew default input
rlabel metal2 s 5170 0 5226 480 6 ccff_tail
port 15 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[0]
port 16 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[10]
port 17 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[11]
port 18 nsew default input
rlabel metal3 s 0 13744 480 13864 6 chanx_left_in[12]
port 19 nsew default input
rlabel metal3 s 0 14152 480 14272 6 chanx_left_in[13]
port 20 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[14]
port 21 nsew default input
rlabel metal3 s 0 14968 480 15088 6 chanx_left_in[15]
port 22 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[16]
port 23 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[17]
port 24 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_in[18]
port 25 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_in[19]
port 26 nsew default input
rlabel metal3 s 0 9256 480 9376 6 chanx_left_in[1]
port 27 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[2]
port 28 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[3]
port 29 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[4]
port 30 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[5]
port 31 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[6]
port 32 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[7]
port 33 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_left_in[8]
port 34 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[9]
port 35 nsew default input
rlabel metal3 s 0 552 480 672 6 chanx_left_out[0]
port 36 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 chanx_left_out[10]
port 37 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[11]
port 38 nsew default tristate
rlabel metal3 s 0 5448 480 5568 6 chanx_left_out[12]
port 39 nsew default tristate
rlabel metal3 s 0 5856 480 5976 6 chanx_left_out[13]
port 40 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[14]
port 41 nsew default tristate
rlabel metal3 s 0 6672 480 6792 6 chanx_left_out[15]
port 42 nsew default tristate
rlabel metal3 s 0 7080 480 7200 6 chanx_left_out[16]
port 43 nsew default tristate
rlabel metal3 s 0 7488 480 7608 6 chanx_left_out[17]
port 44 nsew default tristate
rlabel metal3 s 0 7896 480 8016 6 chanx_left_out[18]
port 45 nsew default tristate
rlabel metal3 s 0 8304 480 8424 6 chanx_left_out[19]
port 46 nsew default tristate
rlabel metal3 s 0 960 480 1080 6 chanx_left_out[1]
port 47 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 48 nsew default tristate
rlabel metal3 s 0 1776 480 1896 6 chanx_left_out[3]
port 49 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[4]
port 50 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[5]
port 51 nsew default tristate
rlabel metal3 s 0 3000 480 3120 6 chanx_left_out[6]
port 52 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[7]
port 53 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[8]
port 54 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_out[9]
port 55 nsew default tristate
rlabel metal3 s 19520 8576 20000 8696 6 chanx_right_in[0]
port 56 nsew default input
rlabel metal3 s 19520 12792 20000 12912 6 chanx_right_in[10]
port 57 nsew default input
rlabel metal3 s 19520 13200 20000 13320 6 chanx_right_in[11]
port 58 nsew default input
rlabel metal3 s 19520 13744 20000 13864 6 chanx_right_in[12]
port 59 nsew default input
rlabel metal3 s 19520 14152 20000 14272 6 chanx_right_in[13]
port 60 nsew default input
rlabel metal3 s 19520 14560 20000 14680 6 chanx_right_in[14]
port 61 nsew default input
rlabel metal3 s 19520 14968 20000 15088 6 chanx_right_in[15]
port 62 nsew default input
rlabel metal3 s 19520 15376 20000 15496 6 chanx_right_in[16]
port 63 nsew default input
rlabel metal3 s 19520 15784 20000 15904 6 chanx_right_in[17]
port 64 nsew default input
rlabel metal3 s 19520 16192 20000 16312 6 chanx_right_in[18]
port 65 nsew default input
rlabel metal3 s 19520 16600 20000 16720 6 chanx_right_in[19]
port 66 nsew default input
rlabel metal3 s 19520 8984 20000 9104 6 chanx_right_in[1]
port 67 nsew default input
rlabel metal3 s 19520 9392 20000 9512 6 chanx_right_in[2]
port 68 nsew default input
rlabel metal3 s 19520 9800 20000 9920 6 chanx_right_in[3]
port 69 nsew default input
rlabel metal3 s 19520 10344 20000 10464 6 chanx_right_in[4]
port 70 nsew default input
rlabel metal3 s 19520 10752 20000 10872 6 chanx_right_in[5]
port 71 nsew default input
rlabel metal3 s 19520 11160 20000 11280 6 chanx_right_in[6]
port 72 nsew default input
rlabel metal3 s 19520 11568 20000 11688 6 chanx_right_in[7]
port 73 nsew default input
rlabel metal3 s 19520 11976 20000 12096 6 chanx_right_in[8]
port 74 nsew default input
rlabel metal3 s 19520 12384 20000 12504 6 chanx_right_in[9]
port 75 nsew default input
rlabel metal3 s 19520 144 20000 264 6 chanx_right_out[0]
port 76 nsew default tristate
rlabel metal3 s 19520 4360 20000 4480 6 chanx_right_out[10]
port 77 nsew default tristate
rlabel metal3 s 19520 4768 20000 4888 6 chanx_right_out[11]
port 78 nsew default tristate
rlabel metal3 s 19520 5176 20000 5296 6 chanx_right_out[12]
port 79 nsew default tristate
rlabel metal3 s 19520 5584 20000 5704 6 chanx_right_out[13]
port 80 nsew default tristate
rlabel metal3 s 19520 5992 20000 6112 6 chanx_right_out[14]
port 81 nsew default tristate
rlabel metal3 s 19520 6400 20000 6520 6 chanx_right_out[15]
port 82 nsew default tristate
rlabel metal3 s 19520 6944 20000 7064 6 chanx_right_out[16]
port 83 nsew default tristate
rlabel metal3 s 19520 7352 20000 7472 6 chanx_right_out[17]
port 84 nsew default tristate
rlabel metal3 s 19520 7760 20000 7880 6 chanx_right_out[18]
port 85 nsew default tristate
rlabel metal3 s 19520 8168 20000 8288 6 chanx_right_out[19]
port 86 nsew default tristate
rlabel metal3 s 19520 552 20000 672 6 chanx_right_out[1]
port 87 nsew default tristate
rlabel metal3 s 19520 960 20000 1080 6 chanx_right_out[2]
port 88 nsew default tristate
rlabel metal3 s 19520 1368 20000 1488 6 chanx_right_out[3]
port 89 nsew default tristate
rlabel metal3 s 19520 1776 20000 1896 6 chanx_right_out[4]
port 90 nsew default tristate
rlabel metal3 s 19520 2184 20000 2304 6 chanx_right_out[5]
port 91 nsew default tristate
rlabel metal3 s 19520 2592 20000 2712 6 chanx_right_out[6]
port 92 nsew default tristate
rlabel metal3 s 19520 3000 20000 3120 6 chanx_right_out[7]
port 93 nsew default tristate
rlabel metal3 s 19520 3544 20000 3664 6 chanx_right_out[8]
port 94 nsew default tristate
rlabel metal3 s 19520 3952 20000 4072 6 chanx_right_out[9]
port 95 nsew default tristate
rlabel metal2 s 6642 0 6698 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 96 nsew default tristate
rlabel metal2 s 7102 0 7158 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 97 nsew default tristate
rlabel metal2 s 7654 0 7710 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 98 nsew default tristate
rlabel metal2 s 8114 0 8170 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 99 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 100 nsew default tristate
rlabel metal2 s 9126 0 9182 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 101 nsew default tristate
rlabel metal2 s 9678 0 9734 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 102 nsew default tristate
rlabel metal2 s 10138 0 10194 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 103 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 104 nsew default tristate
rlabel metal2 s 11150 0 11206 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 105 nsew default input
rlabel metal2 s 11610 0 11666 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 106 nsew default input
rlabel metal2 s 12162 0 12218 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 107 nsew default input
rlabel metal2 s 12622 0 12678 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 108 nsew default input
rlabel metal2 s 13174 0 13230 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 109 nsew default input
rlabel metal2 s 13634 0 13690 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 110 nsew default input
rlabel metal2 s 14094 0 14150 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 111 nsew default input
rlabel metal2 s 14646 0 14702 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 112 nsew default input
rlabel metal2 s 15106 0 15162 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 113 nsew default input
rlabel metal2 s 15658 0 15714 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 114 nsew default tristate
rlabel metal2 s 16118 0 16174 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 115 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 116 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 117 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 118 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 119 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 120 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 121 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 122 nsew default tristate
rlabel metal2 s 8022 16520 8078 17000 6 prog_clk_0_N_in
port 123 nsew default input
rlabel metal3 s 0 144 480 264 6 prog_clk_0_W_out
port 124 nsew default tristate
rlabel metal2 s 8666 16520 8722 17000 6 top_width_0_height_0__pin_0_
port 125 nsew default input
rlabel metal2 s 11886 16520 11942 17000 6 top_width_0_height_0__pin_10_
port 126 nsew default input
rlabel metal2 s 14462 16520 14518 17000 6 top_width_0_height_0__pin_11_lower
port 127 nsew default tristate
rlabel metal2 s 3514 16520 3570 17000 6 top_width_0_height_0__pin_11_upper
port 128 nsew default tristate
rlabel metal2 s 12530 16520 12586 17000 6 top_width_0_height_0__pin_12_
port 129 nsew default input
rlabel metal2 s 15106 16520 15162 17000 6 top_width_0_height_0__pin_13_lower
port 130 nsew default tristate
rlabel metal2 s 4158 16520 4214 17000 6 top_width_0_height_0__pin_13_upper
port 131 nsew default tristate
rlabel metal2 s 13174 16520 13230 17000 6 top_width_0_height_0__pin_14_
port 132 nsew default input
rlabel metal2 s 15750 16520 15806 17000 6 top_width_0_height_0__pin_15_lower
port 133 nsew default tristate
rlabel metal2 s 4802 16520 4858 17000 6 top_width_0_height_0__pin_15_upper
port 134 nsew default tristate
rlabel metal2 s 13818 16520 13874 17000 6 top_width_0_height_0__pin_16_
port 135 nsew default input
rlabel metal2 s 16394 16520 16450 17000 6 top_width_0_height_0__pin_17_lower
port 136 nsew default tristate
rlabel metal2 s 5446 16520 5502 17000 6 top_width_0_height_0__pin_17_upper
port 137 nsew default tristate
rlabel metal2 s 17038 16520 17094 17000 6 top_width_0_height_0__pin_1_lower
port 138 nsew default tristate
rlabel metal2 s 294 16520 350 17000 6 top_width_0_height_0__pin_1_upper
port 139 nsew default tristate
rlabel metal2 s 9310 16520 9366 17000 6 top_width_0_height_0__pin_2_
port 140 nsew default input
rlabel metal2 s 17682 16520 17738 17000 6 top_width_0_height_0__pin_3_lower
port 141 nsew default tristate
rlabel metal2 s 938 16520 994 17000 6 top_width_0_height_0__pin_3_upper
port 142 nsew default tristate
rlabel metal2 s 9954 16520 10010 17000 6 top_width_0_height_0__pin_4_
port 143 nsew default input
rlabel metal2 s 18326 16520 18382 17000 6 top_width_0_height_0__pin_5_lower
port 144 nsew default tristate
rlabel metal2 s 1582 16520 1638 17000 6 top_width_0_height_0__pin_5_upper
port 145 nsew default tristate
rlabel metal2 s 10598 16520 10654 17000 6 top_width_0_height_0__pin_6_
port 146 nsew default input
rlabel metal2 s 18970 16520 19026 17000 6 top_width_0_height_0__pin_7_lower
port 147 nsew default tristate
rlabel metal2 s 2226 16520 2282 17000 6 top_width_0_height_0__pin_7_upper
port 148 nsew default tristate
rlabel metal2 s 11242 16520 11298 17000 6 top_width_0_height_0__pin_8_
port 149 nsew default input
rlabel metal2 s 19614 16520 19670 17000 6 top_width_0_height_0__pin_9_lower
port 150 nsew default tristate
rlabel metal2 s 2870 16520 2926 17000 6 top_width_0_height_0__pin_9_upper
port 151 nsew default tristate
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 152 nsew default input
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 153 nsew default input
<< properties >>
string FIXED_BBOX 0 0 20000 17000
<< end >>
