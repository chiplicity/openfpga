magic
tech EFS8A
magscale 1 2
timestamp 1602527948
<< locali >>
rect 10091 24225 10218 24259
rect 24627 23137 24662 23171
rect 7331 20961 7366 20995
rect 2455 18785 2490 18819
rect 18291 17833 18337 17867
rect 24627 17697 24662 17731
rect 12771 15113 12909 15147
rect 7791 14501 7836 14535
rect 14415 13753 14599 13787
rect 9597 11679 9631 11781
rect 14559 11543 14593 11611
rect 14559 11509 14565 11543
rect 24627 11169 24662 11203
rect 7665 9911 7699 10217
rect 2547 8993 2582 9027
rect 22787 8993 22914 9027
rect 7573 7259 7607 7429
rect 24731 4233 24869 4267
rect 11799 3689 11805 3723
rect 11799 3621 11833 3689
rect 9919 3145 10057 3179
rect 7067 2601 7205 2635
<< viali >>
rect 6412 24225 6446 24259
rect 7456 24225 7490 24259
rect 8436 24225 8470 24259
rect 10057 24225 10091 24259
rect 6515 24021 6549 24055
rect 7527 24021 7561 24055
rect 8539 24021 8573 24055
rect 10287 24021 10321 24055
rect 2789 23817 2823 23851
rect 6377 23817 6411 23851
rect 7021 23817 7055 23851
rect 8309 23817 8343 23851
rect 10977 23817 11011 23851
rect 14013 23817 14047 23851
rect 19993 23817 20027 23851
rect 21925 23817 21959 23851
rect 25145 23817 25179 23851
rect 4629 23749 4663 23783
rect 7573 23681 7607 23715
rect 8493 23681 8527 23715
rect 2304 23613 2338 23647
rect 4236 23613 4270 23647
rect 6837 23613 6871 23647
rect 9873 23613 9907 23647
rect 10057 23613 10091 23647
rect 13829 23613 13863 23647
rect 14381 23613 14415 23647
rect 18128 23613 18162 23647
rect 19508 23613 19542 23647
rect 21440 23613 21474 23647
rect 24644 23613 24678 23647
rect 7941 23545 7975 23579
rect 8585 23545 8619 23579
rect 9137 23545 9171 23579
rect 9965 23545 9999 23579
rect 24731 23545 24765 23579
rect 2375 23477 2409 23511
rect 4307 23477 4341 23511
rect 18199 23477 18233 23511
rect 18613 23477 18647 23511
rect 19579 23477 19613 23511
rect 21511 23477 21545 23511
rect 6837 23273 6871 23307
rect 5549 23205 5583 23239
rect 8217 23205 8251 23239
rect 9873 23205 9907 23239
rect 1444 23137 1478 23171
rect 24593 23137 24627 23171
rect 5457 23069 5491 23103
rect 6101 23069 6135 23103
rect 7021 23069 7055 23103
rect 8125 23069 8159 23103
rect 8769 23069 8803 23103
rect 9781 23069 9815 23103
rect 7573 23001 7607 23035
rect 9137 23001 9171 23035
rect 10333 23001 10367 23035
rect 1547 22933 1581 22967
rect 24731 22933 24765 22967
rect 1593 22729 1627 22763
rect 9781 22729 9815 22763
rect 10149 22729 10183 22763
rect 12633 22729 12667 22763
rect 24685 22729 24719 22763
rect 5917 22593 5951 22627
rect 6193 22593 6227 22627
rect 7205 22593 7239 22627
rect 8585 22593 8619 22627
rect 8861 22593 8895 22627
rect 5089 22525 5123 22559
rect 5825 22525 5859 22559
rect 12449 22525 12483 22559
rect 13001 22525 13035 22559
rect 6929 22457 6963 22491
rect 7021 22457 7055 22491
rect 8677 22457 8711 22491
rect 6561 22389 6595 22423
rect 8033 22389 8067 22423
rect 5457 22185 5491 22219
rect 6929 22185 6963 22219
rect 7849 22185 7883 22219
rect 8033 22117 8067 22151
rect 8677 22049 8711 22083
rect 11320 22049 11354 22083
rect 12792 22049 12826 22083
rect 9045 21845 9079 21879
rect 11391 21845 11425 21879
rect 12541 21845 12575 21879
rect 12863 21845 12897 21879
rect 11023 21641 11057 21675
rect 11437 21641 11471 21675
rect 13553 21641 13587 21675
rect 12541 21505 12575 21539
rect 12817 21505 12851 21539
rect 10952 21437 10986 21471
rect 11713 21437 11747 21471
rect 12265 21369 12299 21403
rect 12633 21369 12667 21403
rect 8125 21301 8159 21335
rect 9689 21301 9723 21335
rect 11897 21029 11931 21063
rect 11989 21029 12023 21063
rect 7297 20961 7331 20995
rect 10333 20961 10367 20995
rect 12449 20825 12483 20859
rect 7435 20757 7469 20791
rect 8493 20757 8527 20791
rect 9965 20757 9999 20791
rect 7297 20553 7331 20587
rect 9597 20553 9631 20587
rect 9965 20553 9999 20587
rect 11069 20553 11103 20587
rect 11529 20553 11563 20587
rect 12725 20553 12759 20587
rect 8585 20417 8619 20451
rect 10149 20417 10183 20451
rect 10793 20417 10827 20451
rect 12541 20349 12575 20383
rect 8401 20281 8435 20315
rect 8677 20281 8711 20315
rect 9229 20281 9263 20315
rect 10241 20281 10275 20315
rect 11897 20213 11931 20247
rect 12173 20213 12207 20247
rect 5733 20009 5767 20043
rect 13093 20009 13127 20043
rect 6009 19941 6043 19975
rect 8217 19941 8251 19975
rect 9873 19941 9907 19975
rect 10425 19941 10459 19975
rect 11253 19941 11287 19975
rect 11345 19873 11379 19907
rect 12909 19873 12943 19907
rect 4813 19805 4847 19839
rect 5917 19805 5951 19839
rect 6193 19805 6227 19839
rect 8125 19805 8159 19839
rect 8769 19805 8803 19839
rect 9781 19805 9815 19839
rect 7849 19669 7883 19703
rect 6193 19465 6227 19499
rect 6561 19465 6595 19499
rect 8125 19465 8159 19499
rect 9689 19465 9723 19499
rect 10057 19465 10091 19499
rect 10333 19465 10367 19499
rect 11345 19465 11379 19499
rect 14657 19465 14691 19499
rect 12587 19397 12621 19431
rect 13277 19397 13311 19431
rect 5273 19329 5307 19363
rect 5549 19329 5583 19363
rect 6929 19261 6963 19295
rect 8769 19261 8803 19295
rect 12516 19261 12550 19295
rect 14172 19261 14206 19295
rect 5365 19193 5399 19227
rect 6837 19193 6871 19227
rect 9090 19193 9124 19227
rect 5089 19125 5123 19159
rect 8585 19125 8619 19159
rect 13001 19125 13035 19159
rect 14243 19125 14277 19159
rect 3157 18921 3191 18955
rect 4261 18921 4295 18955
rect 6469 18921 6503 18955
rect 8033 18921 8067 18955
rect 12173 18921 12207 18955
rect 5181 18853 5215 18887
rect 5911 18853 5945 18887
rect 11615 18853 11649 18887
rect 1476 18785 1510 18819
rect 2421 18785 2455 18819
rect 4077 18785 4111 18819
rect 7757 18785 7791 18819
rect 8217 18785 8251 18819
rect 5549 18717 5583 18751
rect 11253 18717 11287 18751
rect 13001 18717 13035 18751
rect 1547 18649 1581 18683
rect 2559 18581 2593 18615
rect 8769 18581 8803 18615
rect 10885 18581 10919 18615
rect 1961 18377 1995 18411
rect 2513 18377 2547 18411
rect 8953 18377 8987 18411
rect 18245 18377 18279 18411
rect 4261 18309 4295 18343
rect 3249 18241 3283 18275
rect 4721 18241 4755 18275
rect 5733 18241 5767 18275
rect 7205 18241 7239 18275
rect 8033 18241 8067 18275
rect 12541 18241 12575 18275
rect 1409 18173 1443 18207
rect 5089 18173 5123 18207
rect 5181 18173 5215 18207
rect 5641 18173 5675 18207
rect 11437 18173 11471 18207
rect 18061 18173 18095 18207
rect 18613 18173 18647 18207
rect 23740 18173 23774 18207
rect 24133 18173 24167 18207
rect 3065 18105 3099 18139
rect 3341 18105 3375 18139
rect 3893 18105 3927 18139
rect 8354 18105 8388 18139
rect 11529 18105 11563 18139
rect 12173 18105 12207 18139
rect 12633 18105 12667 18139
rect 13185 18105 13219 18139
rect 1593 18037 1627 18071
rect 6193 18037 6227 18071
rect 7573 18037 7607 18071
rect 7849 18037 7883 18071
rect 10701 18037 10735 18071
rect 11805 18037 11839 18071
rect 23811 18037 23845 18071
rect 1685 17833 1719 17867
rect 6561 17833 6595 17867
rect 11805 17833 11839 17867
rect 12541 17833 12575 17867
rect 14335 17833 14369 17867
rect 18337 17833 18371 17867
rect 2513 17765 2547 17799
rect 2605 17765 2639 17799
rect 4077 17765 4111 17799
rect 5962 17765 5996 17799
rect 8769 17765 8803 17799
rect 11206 17765 11240 17799
rect 12817 17765 12851 17799
rect 4629 17697 4663 17731
rect 8033 17697 8067 17731
rect 8493 17697 8527 17731
rect 14264 17697 14298 17731
rect 18220 17697 18254 17731
rect 24593 17697 24627 17731
rect 3157 17629 3191 17663
rect 5641 17629 5675 17663
rect 10885 17629 10919 17663
rect 12725 17629 12759 17663
rect 13185 17629 13219 17663
rect 5273 17493 5307 17527
rect 7757 17493 7791 17527
rect 10609 17493 10643 17527
rect 24731 17493 24765 17527
rect 2789 17289 2823 17323
rect 4629 17289 4663 17323
rect 4905 17289 4939 17323
rect 6009 17289 6043 17323
rect 8953 17289 8987 17323
rect 13461 17289 13495 17323
rect 24685 17289 24719 17323
rect 2513 17221 2547 17255
rect 7481 17221 7515 17255
rect 10425 17153 10459 17187
rect 12541 17153 12575 17187
rect 12909 17153 12943 17187
rect 14013 17153 14047 17187
rect 3709 17085 3743 17119
rect 8033 17085 8067 17119
rect 9229 17085 9263 17119
rect 10609 17085 10643 17119
rect 13921 17085 13955 17119
rect 14105 17085 14139 17119
rect 18153 17085 18187 17119
rect 3617 17017 3651 17051
rect 4030 17017 4064 17051
rect 5641 17017 5675 17051
rect 7849 17017 7883 17051
rect 8354 17017 8388 17051
rect 10930 17017 10964 17051
rect 12633 17017 12667 17051
rect 18061 17017 18095 17051
rect 7113 16949 7147 16983
rect 10149 16949 10183 16983
rect 11529 16949 11563 16983
rect 12265 16949 12299 16983
rect 15025 16949 15059 16983
rect 17509 16949 17543 16983
rect 17877 16949 17911 16983
rect 4721 16745 4755 16779
rect 5825 16745 5859 16779
rect 8769 16745 8803 16779
rect 12541 16745 12575 16779
rect 8170 16677 8204 16711
rect 10425 16677 10459 16711
rect 10885 16677 10919 16711
rect 11437 16677 11471 16711
rect 13829 16677 13863 16711
rect 14381 16677 14415 16711
rect 17693 16677 17727 16711
rect 5549 16609 5583 16643
rect 6101 16609 6135 16643
rect 9689 16609 9723 16643
rect 10241 16609 10275 16643
rect 11989 16609 12023 16643
rect 12817 16609 12851 16643
rect 7849 16541 7883 16575
rect 11345 16541 11379 16575
rect 13737 16541 13771 16575
rect 17601 16541 17635 16575
rect 19073 16541 19107 16575
rect 18153 16473 18187 16507
rect 3249 16405 3283 16439
rect 3709 16405 3743 16439
rect 7757 16405 7791 16439
rect 14749 16405 14783 16439
rect 18521 16405 18555 16439
rect 7757 16201 7791 16235
rect 11345 16201 11379 16235
rect 17233 16201 17267 16235
rect 17601 16201 17635 16235
rect 25145 16201 25179 16235
rect 3709 16065 3743 16099
rect 4813 16065 4847 16099
rect 5273 16065 5307 16099
rect 8861 16065 8895 16099
rect 10333 16065 10367 16099
rect 13277 16065 13311 16099
rect 14105 16065 14139 16099
rect 14657 16065 14691 16099
rect 18429 16065 18463 16099
rect 3065 15997 3099 16031
rect 3433 15997 3467 16031
rect 3617 15997 3651 16031
rect 7849 15997 7883 16031
rect 8401 15997 8435 16031
rect 10057 15997 10091 16031
rect 10241 15997 10275 16031
rect 24660 15997 24694 16031
rect 4905 15929 4939 15963
rect 14381 15929 14415 15963
rect 14473 15929 14507 15963
rect 18153 15929 18187 15963
rect 18245 15929 18279 15963
rect 4537 15861 4571 15895
rect 5733 15861 5767 15895
rect 6193 15861 6227 15895
rect 7297 15861 7331 15895
rect 7941 15861 7975 15895
rect 9229 15861 9263 15895
rect 9597 15861 9631 15895
rect 11621 15861 11655 15895
rect 13829 15861 13863 15895
rect 19073 15861 19107 15895
rect 24731 15861 24765 15895
rect 6469 15657 6503 15691
rect 8217 15657 8251 15691
rect 13921 15657 13955 15691
rect 14657 15657 14691 15691
rect 17141 15657 17175 15691
rect 4950 15589 4984 15623
rect 16542 15589 16576 15623
rect 18153 15589 18187 15623
rect 18705 15589 18739 15623
rect 24317 15589 24351 15623
rect 24869 15589 24903 15623
rect 5549 15521 5583 15555
rect 6653 15521 6687 15555
rect 6929 15521 6963 15555
rect 8217 15521 8251 15555
rect 8493 15521 8527 15555
rect 9873 15521 9907 15555
rect 11596 15521 11630 15555
rect 13737 15521 13771 15555
rect 2973 15453 3007 15487
rect 4629 15453 4663 15487
rect 7849 15453 7883 15487
rect 10517 15453 10551 15487
rect 16221 15453 16255 15487
rect 18061 15453 18095 15487
rect 24225 15453 24259 15487
rect 7481 15317 7515 15351
rect 10333 15317 10367 15351
rect 11667 15317 11701 15351
rect 6469 15113 6503 15147
rect 8493 15113 8527 15147
rect 12909 15113 12943 15147
rect 13185 15113 13219 15147
rect 14565 15113 14599 15147
rect 19073 15113 19107 15147
rect 25053 15113 25087 15147
rect 5917 15045 5951 15079
rect 8125 15045 8159 15079
rect 13461 15045 13495 15079
rect 15945 15045 15979 15079
rect 18705 15045 18739 15079
rect 4997 14977 5031 15011
rect 5273 14977 5307 15011
rect 7573 14977 7607 15011
rect 10333 14977 10367 15011
rect 17325 14977 17359 15011
rect 19441 14977 19475 15011
rect 24409 14977 24443 15011
rect 24685 14977 24719 15011
rect 3249 14909 3283 14943
rect 3985 14909 4019 14943
rect 9229 14909 9263 14943
rect 12265 14909 12299 14943
rect 12668 14909 12702 14943
rect 13645 14909 13679 14943
rect 14841 14909 14875 14943
rect 16129 14909 16163 14943
rect 23489 14909 23523 14943
rect 24041 14909 24075 14943
rect 4077 14841 4111 14875
rect 5089 14841 5123 14875
rect 7665 14841 7699 14875
rect 10425 14841 10459 14875
rect 10977 14841 11011 14875
rect 13966 14841 14000 14875
rect 16450 14841 16484 14875
rect 18153 14841 18187 14875
rect 18245 14841 18279 14875
rect 4629 14773 4663 14807
rect 7113 14773 7147 14807
rect 8861 14773 8895 14807
rect 9413 14773 9447 14807
rect 9689 14773 9723 14807
rect 10149 14773 10183 14807
rect 11621 14773 11655 14807
rect 15577 14773 15611 14807
rect 17049 14773 17083 14807
rect 17877 14773 17911 14807
rect 1593 14569 1627 14603
rect 5089 14569 5123 14603
rect 5549 14569 5583 14603
rect 8401 14569 8435 14603
rect 12449 14569 12483 14603
rect 16129 14569 16163 14603
rect 17969 14569 18003 14603
rect 7297 14501 7331 14535
rect 7757 14501 7791 14535
rect 10010 14501 10044 14535
rect 11621 14501 11655 14535
rect 13921 14501 13955 14535
rect 16910 14501 16944 14535
rect 18337 14501 18371 14535
rect 24225 14501 24259 14535
rect 24777 14501 24811 14535
rect 1409 14433 1443 14467
rect 4721 14433 4755 14467
rect 6009 14433 6043 14467
rect 6653 14433 6687 14467
rect 13185 14433 13219 14467
rect 13737 14433 13771 14467
rect 14197 14433 14231 14467
rect 18429 14433 18463 14467
rect 7481 14365 7515 14399
rect 9689 14365 9723 14399
rect 11529 14365 11563 14399
rect 11805 14365 11839 14399
rect 16589 14365 16623 14399
rect 24133 14365 24167 14399
rect 4353 14229 4387 14263
rect 9045 14229 9079 14263
rect 10609 14229 10643 14263
rect 15485 14229 15519 14263
rect 17509 14229 17543 14263
rect 1685 14025 1719 14059
rect 2927 14025 2961 14059
rect 6009 14025 6043 14059
rect 8861 14025 8895 14059
rect 10057 14025 10091 14059
rect 11989 14025 12023 14059
rect 16681 14025 16715 14059
rect 18429 14025 18463 14059
rect 6653 13957 6687 13991
rect 8125 13957 8159 13991
rect 2697 13889 2731 13923
rect 4629 13889 4663 13923
rect 11345 13889 11379 13923
rect 11621 13889 11655 13923
rect 14289 13889 14323 13923
rect 16957 13889 16991 13923
rect 2824 13821 2858 13855
rect 9045 13821 9079 13855
rect 9597 13821 9631 13855
rect 10517 13821 10551 13855
rect 10701 13821 10735 13855
rect 12449 13821 12483 13855
rect 13553 13821 13587 13855
rect 14013 13821 14047 13855
rect 15117 13821 15151 13855
rect 15577 13821 15611 13855
rect 15853 13821 15887 13855
rect 3433 13753 3467 13787
rect 4353 13753 4387 13787
rect 4445 13753 4479 13787
rect 7297 13753 7331 13787
rect 7573 13753 7607 13787
rect 7665 13753 7699 13787
rect 9781 13753 9815 13787
rect 14381 13753 14415 13787
rect 3801 13685 3835 13719
rect 4169 13685 4203 13719
rect 8493 13685 8527 13719
rect 12633 13685 12667 13719
rect 13185 13685 13219 13719
rect 14933 13685 14967 13719
rect 24041 13685 24075 13719
rect 24501 13685 24535 13719
rect 7573 13481 7607 13515
rect 7849 13481 7883 13515
rect 9873 13481 9907 13515
rect 15577 13481 15611 13515
rect 4261 13413 4295 13447
rect 7205 13413 7239 13447
rect 11161 13413 11195 13447
rect 12173 13413 12207 13447
rect 12725 13413 12759 13447
rect 6285 13345 6319 13379
rect 8033 13345 8067 13379
rect 8309 13345 8343 13379
rect 11069 13345 11103 13379
rect 13645 13345 13679 13379
rect 15301 13345 15335 13379
rect 15761 13345 15795 13379
rect 2973 13277 3007 13311
rect 4169 13277 4203 13311
rect 4445 13277 4479 13311
rect 6745 13277 6779 13311
rect 12081 13277 12115 13311
rect 8861 13141 8895 13175
rect 11897 13141 11931 13175
rect 13185 13141 13219 13175
rect 13829 13141 13863 13175
rect 3617 12937 3651 12971
rect 4997 12937 5031 12971
rect 5917 12937 5951 12971
rect 6285 12937 6319 12971
rect 6653 12937 6687 12971
rect 8861 12937 8895 12971
rect 10425 12937 10459 12971
rect 11989 12937 12023 12971
rect 13553 12937 13587 12971
rect 13829 12937 13863 12971
rect 15301 12937 15335 12971
rect 8677 12869 8711 12903
rect 1869 12801 1903 12835
rect 5549 12801 5583 12835
rect 6929 12801 6963 12835
rect 7205 12801 7239 12835
rect 8769 12801 8803 12835
rect 9413 12801 9447 12835
rect 12817 12801 12851 12835
rect 14105 12801 14139 12835
rect 14381 12801 14415 12835
rect 1476 12733 1510 12767
rect 3249 12733 3283 12767
rect 4077 12733 4111 12767
rect 8548 12733 8582 12767
rect 10609 12733 10643 12767
rect 3985 12665 4019 12699
rect 4439 12665 4473 12699
rect 7021 12665 7055 12699
rect 8401 12665 8435 12699
rect 10149 12665 10183 12699
rect 10930 12665 10964 12699
rect 12541 12665 12575 12699
rect 12633 12665 12667 12699
rect 14197 12665 14231 12699
rect 1547 12597 1581 12631
rect 7849 12597 7883 12631
rect 8217 12597 8251 12631
rect 11529 12597 11563 12631
rect 15669 12597 15703 12631
rect 4261 12393 4295 12427
rect 6377 12393 6411 12427
rect 11805 12393 11839 12427
rect 12265 12393 12299 12427
rect 12633 12393 12667 12427
rect 14565 12393 14599 12427
rect 18153 12393 18187 12427
rect 5778 12325 5812 12359
rect 7389 12325 7423 12359
rect 10425 12325 10459 12359
rect 11069 12325 11103 12359
rect 13093 12325 13127 12359
rect 9689 12257 9723 12291
rect 10241 12257 10275 12291
rect 15393 12257 15427 12291
rect 5457 12189 5491 12223
rect 7297 12189 7331 12223
rect 7573 12189 7607 12223
rect 13001 12189 13035 12223
rect 13553 12121 13587 12155
rect 6929 12053 6963 12087
rect 8401 12053 8435 12087
rect 8769 12053 8803 12087
rect 10701 12053 10735 12087
rect 14289 12053 14323 12087
rect 15761 12053 15795 12087
rect 5641 11849 5675 11883
rect 7297 11849 7331 11883
rect 7849 11849 7883 11883
rect 8539 11849 8573 11883
rect 9045 11849 9079 11883
rect 9689 11849 9723 11883
rect 10130 11849 10164 11883
rect 10977 11849 11011 11883
rect 12173 11849 12207 11883
rect 13369 11849 13403 11883
rect 13645 11849 13679 11883
rect 15117 11849 15151 11883
rect 15761 11849 15795 11883
rect 7002 11781 7036 11815
rect 8677 11781 8711 11815
rect 9597 11781 9631 11815
rect 10241 11781 10275 11815
rect 4537 11713 4571 11747
rect 6653 11713 6687 11747
rect 7205 11713 7239 11747
rect 8309 11713 8343 11747
rect 8769 11713 8803 11747
rect 10333 11713 10367 11747
rect 16313 11713 16347 11747
rect 18153 11713 18187 11747
rect 18429 11713 18463 11747
rect 1752 11645 1786 11679
rect 4905 11645 4939 11679
rect 5181 11645 5215 11679
rect 6285 11645 6319 11679
rect 7067 11645 7101 11679
rect 9597 11645 9631 11679
rect 12449 11645 12483 11679
rect 14197 11645 14231 11679
rect 6837 11577 6871 11611
rect 8401 11577 8435 11611
rect 9965 11577 9999 11611
rect 10701 11577 10735 11611
rect 11345 11577 11379 11611
rect 12770 11577 12804 11611
rect 16037 11577 16071 11611
rect 16129 11577 16163 11611
rect 18245 11577 18279 11611
rect 1823 11509 1857 11543
rect 2237 11509 2271 11543
rect 4721 11509 4755 11543
rect 11805 11509 11839 11543
rect 14105 11509 14139 11543
rect 14565 11509 14599 11543
rect 15393 11509 15427 11543
rect 17785 11509 17819 11543
rect 5365 11305 5399 11339
rect 6101 11305 6135 11339
rect 7389 11305 7423 11339
rect 9965 11305 9999 11339
rect 10241 11305 10275 11339
rect 12541 11305 12575 11339
rect 13001 11305 13035 11339
rect 14197 11305 14231 11339
rect 15485 11305 15519 11339
rect 17785 11305 17819 11339
rect 7481 11237 7515 11271
rect 16123 11237 16157 11271
rect 1409 11169 1443 11203
rect 5181 11169 5215 11203
rect 5641 11169 5675 11203
rect 9781 11169 9815 11203
rect 10793 11169 10827 11203
rect 11437 11169 11471 11203
rect 12357 11169 12391 11203
rect 16681 11169 16715 11203
rect 17601 11169 17635 11203
rect 24593 11169 24627 11203
rect 4721 11101 4755 11135
rect 7849 11101 7883 11135
rect 15761 11101 15795 11135
rect 1593 11033 1627 11067
rect 7941 11033 7975 11067
rect 8953 11033 8987 11067
rect 13369 11033 13403 11067
rect 6469 10965 6503 10999
rect 6929 10965 6963 10999
rect 7619 10965 7653 10999
rect 7757 10965 7791 10999
rect 8493 10965 8527 10999
rect 9229 10965 9263 10999
rect 10609 10965 10643 10999
rect 13645 10965 13679 10999
rect 24731 10965 24765 10999
rect 1593 10761 1627 10795
rect 5181 10761 5215 10795
rect 5549 10761 5583 10795
rect 7849 10761 7883 10795
rect 8585 10761 8619 10795
rect 9781 10761 9815 10795
rect 11897 10761 11931 10795
rect 14381 10761 14415 10795
rect 15209 10761 15243 10795
rect 17601 10761 17635 10795
rect 24685 10761 24719 10795
rect 6653 10693 6687 10727
rect 8677 10625 8711 10659
rect 9045 10625 9079 10659
rect 15393 10625 15427 10659
rect 16773 10625 16807 10659
rect 7297 10557 7331 10591
rect 8456 10557 8490 10591
rect 10425 10557 10459 10591
rect 11069 10557 11103 10591
rect 11253 10557 11287 10591
rect 13185 10557 13219 10591
rect 13461 10557 13495 10591
rect 13737 10557 13771 10591
rect 14105 10557 14139 10591
rect 16037 10557 16071 10591
rect 8309 10489 8343 10523
rect 12173 10489 12207 10523
rect 15485 10489 15519 10523
rect 7113 10421 7147 10455
rect 7481 10421 7515 10455
rect 8217 10421 8251 10455
rect 9413 10421 9447 10455
rect 10241 10421 10275 10455
rect 10701 10421 10735 10455
rect 12725 10421 12759 10455
rect 14841 10421 14875 10455
rect 16313 10421 16347 10455
rect 6837 10217 6871 10251
rect 7665 10217 7699 10251
rect 9137 10217 9171 10251
rect 12541 10217 12575 10251
rect 14289 10217 14323 10251
rect 23949 10217 23983 10251
rect 6193 10149 6227 10183
rect 6340 10081 6374 10115
rect 7481 10081 7515 10115
rect 6561 10013 6595 10047
rect 6469 9945 6503 9979
rect 8493 10149 8527 10183
rect 17325 10149 17359 10183
rect 17877 10149 17911 10183
rect 7757 10081 7791 10115
rect 9689 10081 9723 10115
rect 10241 10081 10275 10115
rect 11253 10081 11287 10115
rect 13461 10081 13495 10115
rect 13645 10081 13679 10115
rect 14013 10081 14047 10115
rect 15393 10081 15427 10115
rect 15853 10081 15887 10115
rect 8125 10013 8159 10047
rect 10149 10013 10183 10047
rect 16129 10013 16163 10047
rect 17233 10013 17267 10047
rect 7922 9945 7956 9979
rect 11437 9945 11471 9979
rect 7665 9877 7699 9911
rect 8033 9877 8067 9911
rect 8769 9877 8803 9911
rect 10885 9877 10919 9911
rect 16957 9877 16991 9911
rect 7481 9673 7515 9707
rect 8401 9673 8435 9707
rect 9321 9673 9355 9707
rect 9643 9673 9677 9707
rect 10885 9673 10919 9707
rect 11805 9673 11839 9707
rect 13461 9673 13495 9707
rect 13921 9673 13955 9707
rect 14473 9673 14507 9707
rect 15669 9673 15703 9707
rect 17509 9673 17543 9707
rect 6285 9605 6319 9639
rect 6653 9605 6687 9639
rect 7113 9605 7147 9639
rect 8106 9605 8140 9639
rect 8217 9605 8251 9639
rect 8953 9605 8987 9639
rect 9781 9605 9815 9639
rect 10149 9605 10183 9639
rect 5917 9537 5951 9571
rect 8309 9537 8343 9571
rect 9873 9537 9907 9571
rect 12541 9537 12575 9571
rect 12817 9537 12851 9571
rect 16221 9537 16255 9571
rect 23949 9537 23983 9571
rect 5549 9469 5583 9503
rect 6929 9469 6963 9503
rect 7941 9469 7975 9503
rect 10517 9469 10551 9503
rect 14657 9469 14691 9503
rect 15117 9469 15151 9503
rect 17141 9469 17175 9503
rect 17877 9469 17911 9503
rect 18705 9469 18739 9503
rect 9505 9401 9539 9435
rect 12265 9401 12299 9435
rect 12633 9401 12667 9435
rect 15393 9401 15427 9435
rect 16583 9401 16617 9435
rect 18061 9401 18095 9435
rect 24041 9401 24075 9435
rect 24593 9401 24627 9435
rect 7849 9333 7883 9367
rect 11345 9333 11379 9367
rect 16129 9333 16163 9367
rect 23397 9333 23431 9367
rect 6193 9129 6227 9163
rect 7205 9129 7239 9163
rect 9413 9129 9447 9163
rect 9873 9129 9907 9163
rect 10241 9129 10275 9163
rect 16313 9129 16347 9163
rect 25559 9129 25593 9163
rect 8033 9061 8067 9095
rect 12862 9061 12896 9095
rect 13737 9061 13771 9095
rect 17227 9061 17261 9095
rect 18705 9061 18739 9095
rect 18797 9061 18831 9095
rect 24041 9061 24075 9095
rect 1409 8993 1443 9027
rect 2513 8993 2547 9027
rect 6009 8993 6043 9027
rect 7021 8993 7055 9027
rect 7849 8993 7883 9027
rect 9045 8993 9079 9027
rect 10609 8993 10643 9027
rect 11161 8993 11195 9027
rect 11437 8993 11471 9027
rect 15301 8993 15335 9027
rect 15761 8993 15795 9027
rect 16865 8993 16899 9027
rect 22753 8993 22787 9027
rect 24593 8993 24627 9027
rect 25488 8993 25522 9027
rect 6929 8925 6963 8959
rect 8401 8925 8435 8959
rect 8769 8925 8803 8959
rect 11713 8925 11747 8959
rect 12541 8925 12575 8959
rect 16037 8925 16071 8959
rect 18981 8925 19015 8959
rect 23949 8925 23983 8959
rect 1593 8857 1627 8891
rect 8309 8857 8343 8891
rect 17785 8857 17819 8891
rect 2651 8789 2685 8823
rect 6561 8789 6595 8823
rect 8171 8789 8205 8823
rect 13461 8789 13495 8823
rect 14657 8789 14691 8823
rect 15025 8789 15059 8823
rect 18153 8789 18187 8823
rect 22983 8789 23017 8823
rect 1685 8585 1719 8619
rect 7021 8585 7055 8619
rect 7389 8585 7423 8619
rect 7757 8585 7791 8619
rect 8493 8585 8527 8619
rect 9229 8585 9263 8619
rect 9965 8585 9999 8619
rect 10609 8585 10643 8619
rect 13461 8585 13495 8619
rect 14381 8585 14415 8619
rect 15209 8585 15243 8619
rect 16773 8585 16807 8619
rect 17417 8585 17451 8619
rect 17877 8585 17911 8619
rect 19073 8585 19107 8619
rect 19533 8585 19567 8619
rect 22937 8585 22971 8619
rect 23397 8585 23431 8619
rect 25513 8585 25547 8619
rect 8585 8449 8619 8483
rect 9597 8449 9631 8483
rect 11529 8449 11563 8483
rect 16957 8449 16991 8483
rect 18153 8449 18187 8483
rect 18797 8449 18831 8483
rect 24409 8449 24443 8483
rect 24685 8449 24719 8483
rect 7205 8381 7239 8415
rect 8364 8381 8398 8415
rect 9781 8381 9815 8415
rect 10241 8381 10275 8415
rect 10885 8381 10919 8415
rect 11345 8381 11379 8415
rect 11805 8381 11839 8415
rect 12633 8381 12667 8415
rect 14197 8381 14231 8415
rect 14657 8381 14691 8415
rect 15301 8381 15335 8415
rect 15761 8381 15795 8415
rect 16313 8381 16347 8415
rect 23765 8381 23799 8415
rect 6653 8313 6687 8347
rect 8217 8313 8251 8347
rect 8953 8313 8987 8347
rect 12449 8313 12483 8347
rect 16037 8313 16071 8347
rect 18245 8313 18279 8347
rect 25053 8313 25087 8347
rect 2605 8245 2639 8279
rect 6101 8245 6135 8279
rect 8033 8245 8067 8279
rect 12173 8245 12207 8279
rect 7205 8041 7239 8075
rect 8769 8041 8803 8075
rect 9873 8041 9907 8075
rect 11345 8041 11379 8075
rect 12817 8041 12851 8075
rect 15577 8041 15611 8075
rect 24271 8041 24305 8075
rect 11989 7973 12023 8007
rect 15853 7973 15887 8007
rect 16634 7973 16668 8007
rect 6193 7905 6227 7939
rect 7849 7905 7883 7939
rect 9689 7905 9723 7939
rect 10701 7905 10735 7939
rect 12541 7905 12575 7939
rect 13461 7905 13495 7939
rect 16313 7905 16347 7939
rect 17233 7905 17267 7939
rect 18245 7905 18279 7939
rect 24200 7905 24234 7939
rect 6561 7837 6595 7871
rect 8493 7837 8527 7871
rect 11897 7837 11931 7871
rect 13369 7837 13403 7871
rect 6358 7769 6392 7803
rect 6469 7701 6503 7735
rect 6837 7701 6871 7735
rect 7573 7701 7607 7735
rect 9137 7701 9171 7735
rect 10977 7701 11011 7735
rect 18337 7701 18371 7735
rect 23765 7701 23799 7735
rect 9321 7497 9355 7531
rect 10701 7497 10735 7531
rect 11897 7497 11931 7531
rect 12173 7497 12207 7531
rect 13461 7497 13495 7531
rect 16681 7497 16715 7531
rect 17417 7497 17451 7531
rect 6285 7429 6319 7463
rect 7573 7429 7607 7463
rect 1547 7361 1581 7395
rect 1444 7293 1478 7327
rect 1869 7293 1903 7327
rect 6561 7293 6595 7327
rect 13645 7361 13679 7395
rect 14105 7361 14139 7395
rect 18153 7361 18187 7395
rect 18521 7361 18555 7395
rect 23765 7361 23799 7395
rect 24041 7361 24075 7395
rect 7941 7293 7975 7327
rect 8401 7293 8435 7327
rect 9505 7293 9539 7327
rect 9965 7293 9999 7327
rect 10793 7293 10827 7327
rect 11253 7293 11287 7327
rect 15117 7293 15151 7327
rect 15577 7293 15611 7327
rect 5917 7225 5951 7259
rect 7389 7225 7423 7259
rect 7573 7225 7607 7259
rect 7849 7225 7883 7259
rect 11529 7225 11563 7259
rect 13737 7225 13771 7259
rect 14657 7225 14691 7259
rect 18245 7225 18279 7259
rect 23857 7225 23891 7259
rect 7021 7157 7055 7191
rect 9689 7157 9723 7191
rect 13093 7157 13127 7191
rect 14933 7157 14967 7191
rect 15393 7157 15427 7191
rect 16313 7157 16347 7191
rect 17877 7157 17911 7191
rect 23489 7157 23523 7191
rect 24777 7157 24811 7191
rect 8677 6953 8711 6987
rect 10333 6953 10367 6987
rect 11253 6953 11287 6987
rect 13185 6953 13219 6987
rect 13645 6953 13679 6987
rect 15577 6953 15611 6987
rect 18153 6953 18187 6987
rect 12586 6885 12620 6919
rect 17002 6885 17036 6919
rect 18521 6885 18555 6919
rect 18613 6885 18647 6919
rect 22937 6885 22971 6919
rect 23029 6885 23063 6919
rect 24409 6885 24443 6919
rect 6193 6817 6227 6851
rect 6837 6817 6871 6851
rect 7665 6817 7699 6851
rect 8217 6817 8251 6851
rect 9689 6817 9723 6851
rect 16681 6817 16715 6851
rect 17601 6817 17635 6851
rect 24685 6817 24719 6851
rect 7205 6749 7239 6783
rect 7573 6749 7607 6783
rect 8033 6749 8067 6783
rect 10057 6749 10091 6783
rect 12265 6749 12299 6783
rect 14013 6749 14047 6783
rect 19165 6749 19199 6783
rect 23581 6749 23615 6783
rect 9965 6681 9999 6715
rect 9827 6613 9861 6647
rect 10885 6613 10919 6647
rect 23857 6613 23891 6647
rect 8290 6409 8324 6443
rect 10425 6409 10459 6443
rect 11805 6409 11839 6443
rect 13369 6409 13403 6443
rect 17141 6409 17175 6443
rect 19625 6409 19659 6443
rect 24685 6409 24719 6443
rect 25421 6409 25455 6443
rect 8401 6341 8435 6375
rect 12633 6341 12667 6375
rect 14105 6341 14139 6375
rect 16497 6341 16531 6375
rect 19257 6341 19291 6375
rect 21833 6341 21867 6375
rect 8493 6273 8527 6307
rect 10057 6273 10091 6307
rect 15577 6273 15611 6307
rect 17877 6273 17911 6307
rect 18705 6273 18739 6307
rect 20177 6273 20211 6307
rect 22753 6273 22787 6307
rect 23489 6273 23523 6307
rect 23765 6273 23799 6307
rect 24041 6273 24075 6307
rect 7113 6205 7147 6239
rect 8125 6205 8159 6239
rect 9137 6205 9171 6239
rect 10793 6205 10827 6239
rect 11253 6205 11287 6239
rect 12449 6205 12483 6239
rect 22109 6205 22143 6239
rect 23029 6205 23063 6239
rect 25237 6205 25271 6239
rect 25789 6205 25823 6239
rect 7665 6137 7699 6171
rect 8861 6137 8895 6171
rect 13553 6137 13587 6171
rect 13645 6137 13679 6171
rect 15898 6137 15932 6171
rect 16773 6137 16807 6171
rect 18797 6137 18831 6171
rect 23857 6137 23891 6171
rect 6193 6069 6227 6103
rect 7297 6069 7331 6103
rect 9689 6069 9723 6103
rect 11069 6069 11103 6103
rect 12173 6069 12207 6103
rect 13001 6069 13035 6103
rect 15485 6069 15519 6103
rect 18429 6069 18463 6103
rect 6837 5865 6871 5899
rect 7573 5865 7607 5899
rect 7941 5865 7975 5899
rect 9505 5865 9539 5899
rect 13553 5865 13587 5899
rect 16589 5865 16623 5899
rect 22109 5865 22143 5899
rect 22845 5865 22879 5899
rect 24823 5865 24857 5899
rect 8033 5797 8067 5831
rect 10194 5797 10228 5831
rect 11805 5797 11839 5831
rect 15990 5797 16024 5831
rect 18429 5797 18463 5831
rect 23305 5797 23339 5831
rect 23857 5797 23891 5831
rect 6561 5729 6595 5763
rect 6745 5729 6779 5763
rect 9873 5729 9907 5763
rect 13645 5729 13679 5763
rect 14197 5729 14231 5763
rect 24720 5729 24754 5763
rect 8401 5661 8435 5695
rect 8769 5661 8803 5695
rect 11713 5661 11747 5695
rect 12173 5661 12207 5695
rect 14381 5661 14415 5695
rect 15669 5661 15703 5695
rect 18337 5661 18371 5695
rect 18613 5661 18647 5695
rect 19257 5661 19291 5695
rect 23213 5661 23247 5695
rect 8171 5593 8205 5627
rect 8309 5593 8343 5627
rect 9045 5525 9079 5559
rect 10793 5525 10827 5559
rect 11069 5525 11103 5559
rect 8309 5321 8343 5355
rect 8677 5321 8711 5355
rect 9413 5321 9447 5355
rect 11161 5321 11195 5355
rect 12725 5321 12759 5355
rect 13093 5321 13127 5355
rect 13461 5321 13495 5355
rect 16221 5321 16255 5355
rect 16589 5321 16623 5355
rect 18429 5321 18463 5355
rect 22707 5321 22741 5355
rect 23949 5321 23983 5355
rect 25421 5321 25455 5355
rect 10793 5253 10827 5287
rect 14749 5253 14783 5287
rect 17877 5253 17911 5287
rect 23397 5253 23431 5287
rect 7389 5185 7423 5219
rect 8769 5185 8803 5219
rect 11621 5185 11655 5219
rect 12081 5185 12115 5219
rect 7021 5117 7055 5151
rect 7665 5117 7699 5151
rect 8548 5117 8582 5151
rect 13645 5117 13679 5151
rect 14105 5117 14139 5151
rect 15025 5117 15059 5151
rect 15209 5117 15243 5151
rect 15669 5117 15703 5151
rect 18245 5117 18279 5151
rect 19752 5117 19786 5151
rect 20177 5117 20211 5151
rect 22636 5117 22670 5151
rect 24660 5117 24694 5151
rect 6837 5049 6871 5083
rect 8401 5049 8435 5083
rect 9137 5049 9171 5083
rect 10241 5049 10275 5083
rect 10333 5049 10367 5083
rect 14381 5049 14415 5083
rect 23121 5049 23155 5083
rect 25145 5049 25179 5083
rect 6193 4981 6227 5015
rect 6561 4981 6595 5015
rect 9873 4981 9907 5015
rect 15301 4981 15335 5015
rect 19855 4981 19889 5015
rect 24731 4981 24765 5015
rect 7297 4777 7331 4811
rect 7757 4777 7791 4811
rect 8401 4777 8435 4811
rect 10793 4777 10827 4811
rect 13921 4777 13955 4811
rect 18245 4777 18279 4811
rect 8125 4709 8159 4743
rect 11431 4709 11465 4743
rect 15622 4709 15656 4743
rect 17233 4709 17267 4743
rect 1476 4641 1510 4675
rect 6285 4641 6319 4675
rect 6837 4641 6871 4675
rect 11069 4641 11103 4675
rect 13277 4641 13311 4675
rect 15301 4641 15335 4675
rect 18613 4641 18647 4675
rect 19717 4641 19751 4675
rect 6653 4573 6687 4607
rect 8769 4573 8803 4607
rect 17141 4573 17175 4607
rect 1547 4505 1581 4539
rect 13461 4505 13495 4539
rect 17693 4505 17727 4539
rect 10149 4437 10183 4471
rect 11989 4437 12023 4471
rect 16221 4437 16255 4471
rect 19901 4437 19935 4471
rect 1593 4233 1627 4267
rect 7113 4233 7147 4267
rect 8125 4233 8159 4267
rect 10241 4233 10275 4267
rect 10701 4233 10735 4267
rect 18199 4233 18233 4267
rect 18613 4233 18647 4267
rect 19809 4233 19843 4267
rect 24869 4233 24903 4267
rect 6285 4165 6319 4199
rect 17785 4165 17819 4199
rect 9965 4097 9999 4131
rect 14289 4097 14323 4131
rect 6929 4029 6963 4063
rect 9137 4029 9171 4063
rect 9873 4029 9907 4063
rect 10793 4029 10827 4063
rect 11253 4029 11287 4063
rect 12265 4029 12299 4063
rect 13093 4029 13127 4063
rect 14473 4029 14507 4063
rect 16221 4029 16255 4063
rect 16497 4029 16531 4063
rect 18128 4029 18162 4063
rect 24660 4029 24694 4063
rect 11529 3961 11563 3995
rect 12449 3961 12483 3995
rect 14794 3961 14828 3995
rect 15669 3961 15703 3995
rect 17049 3961 17083 3995
rect 17325 3961 17359 3995
rect 5917 3893 5951 3927
rect 11805 3893 11839 3927
rect 13461 3893 13495 3927
rect 15393 3893 15427 3927
rect 25145 3893 25179 3927
rect 6837 3689 6871 3723
rect 11069 3689 11103 3723
rect 11805 3689 11839 3723
rect 14473 3689 14507 3723
rect 15761 3689 15795 3723
rect 13277 3621 13311 3655
rect 13369 3621 13403 3655
rect 16497 3621 16531 3655
rect 17049 3621 17083 3655
rect 5952 3553 5986 3587
rect 18521 3553 18555 3587
rect 10425 3485 10459 3519
rect 11437 3485 11471 3519
rect 13553 3485 13587 3519
rect 15301 3485 15335 3519
rect 16405 3485 16439 3519
rect 17877 3485 17911 3519
rect 6055 3349 6089 3383
rect 12357 3349 12391 3383
rect 12633 3349 12667 3383
rect 6009 3145 6043 3179
rect 7159 3145 7193 3179
rect 8907 3145 8941 3179
rect 10057 3145 10091 3179
rect 12265 3145 12299 3179
rect 13461 3145 13495 3179
rect 16497 3145 16531 3179
rect 18521 3145 18555 3179
rect 14197 3077 14231 3111
rect 14657 3077 14691 3111
rect 18199 3077 18233 3111
rect 13185 3009 13219 3043
rect 15025 3009 15059 3043
rect 15577 3009 15611 3043
rect 7088 2941 7122 2975
rect 8815 2941 8849 2975
rect 9229 2941 9263 2975
rect 9848 2941 9882 2975
rect 10701 2941 10735 2975
rect 10885 2941 10919 2975
rect 13829 2941 13863 2975
rect 14013 2941 14047 2975
rect 16221 2941 16255 2975
rect 18128 2941 18162 2975
rect 18889 2941 18923 2975
rect 19108 2941 19142 2975
rect 19533 2941 19567 2975
rect 10793 2873 10827 2907
rect 12541 2873 12575 2907
rect 12633 2873 12667 2907
rect 15669 2873 15703 2907
rect 7573 2805 7607 2839
rect 10333 2805 10367 2839
rect 11805 2805 11839 2839
rect 15393 2805 15427 2839
rect 16957 2805 16991 2839
rect 19211 2805 19245 2839
rect 7205 2601 7239 2635
rect 8815 2601 8849 2635
rect 10793 2601 10827 2635
rect 11989 2601 12023 2635
rect 12357 2601 12391 2635
rect 13645 2601 13679 2635
rect 15209 2601 15243 2635
rect 17371 2601 17405 2635
rect 19579 2601 19613 2635
rect 10517 2533 10551 2567
rect 11069 2533 11103 2567
rect 11161 2533 11195 2567
rect 12817 2533 12851 2567
rect 14933 2533 14967 2567
rect 15577 2533 15611 2567
rect 15669 2533 15703 2567
rect 16221 2533 16255 2567
rect 6996 2465 7030 2499
rect 8744 2465 8778 2499
rect 9597 2465 9631 2499
rect 9873 2465 9907 2499
rect 14289 2465 14323 2499
rect 17300 2465 17334 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 19508 2465 19542 2499
rect 19901 2465 19935 2499
rect 21256 2465 21290 2499
rect 9229 2397 9263 2431
rect 12725 2397 12759 2431
rect 13001 2397 13035 2431
rect 14197 2397 14231 2431
rect 10057 2329 10091 2363
rect 11621 2329 11655 2363
rect 14473 2329 14507 2363
rect 18521 2329 18555 2363
rect 7481 2261 7515 2295
rect 17785 2261 17819 2295
rect 21327 2261 21361 2295
rect 21741 2261 21775 2295
<< metal1 >>
rect 23750 27480 23756 27532
rect 23808 27520 23814 27532
rect 25130 27520 25136 27532
rect 23808 27492 25136 27520
rect 23808 27480 23814 27492
rect 25130 27480 25136 27492
rect 25188 27480 25194 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 6270 24216 6276 24268
rect 6328 24256 6334 24268
rect 6400 24259 6458 24265
rect 6400 24256 6412 24259
rect 6328 24228 6412 24256
rect 6328 24216 6334 24228
rect 6400 24225 6412 24228
rect 6446 24225 6458 24259
rect 6400 24219 6458 24225
rect 7444 24259 7502 24265
rect 7444 24225 7456 24259
rect 7490 24256 7502 24259
rect 7558 24256 7564 24268
rect 7490 24228 7564 24256
rect 7490 24225 7502 24228
rect 7444 24219 7502 24225
rect 7558 24216 7564 24228
rect 7616 24216 7622 24268
rect 8294 24216 8300 24268
rect 8352 24256 8358 24268
rect 8424 24259 8482 24265
rect 8424 24256 8436 24259
rect 8352 24228 8436 24256
rect 8352 24216 8358 24228
rect 8424 24225 8436 24228
rect 8470 24225 8482 24259
rect 8424 24219 8482 24225
rect 10045 24259 10103 24265
rect 10045 24225 10057 24259
rect 10091 24256 10103 24259
rect 10134 24256 10140 24268
rect 10091 24228 10140 24256
rect 10091 24225 10103 24228
rect 10045 24219 10103 24225
rect 10134 24216 10140 24228
rect 10192 24216 10198 24268
rect 6362 24012 6368 24064
rect 6420 24052 6426 24064
rect 6503 24055 6561 24061
rect 6503 24052 6515 24055
rect 6420 24024 6515 24052
rect 6420 24012 6426 24024
rect 6503 24021 6515 24024
rect 6549 24021 6561 24055
rect 6503 24015 6561 24021
rect 6822 24012 6828 24064
rect 6880 24052 6886 24064
rect 7515 24055 7573 24061
rect 7515 24052 7527 24055
rect 6880 24024 7527 24052
rect 6880 24012 6886 24024
rect 7515 24021 7527 24024
rect 7561 24021 7573 24055
rect 7515 24015 7573 24021
rect 8527 24055 8585 24061
rect 8527 24021 8539 24055
rect 8573 24052 8585 24055
rect 8662 24052 8668 24064
rect 8573 24024 8668 24052
rect 8573 24021 8585 24024
rect 8527 24015 8585 24021
rect 8662 24012 8668 24024
rect 8720 24012 8726 24064
rect 10042 24012 10048 24064
rect 10100 24052 10106 24064
rect 10275 24055 10333 24061
rect 10275 24052 10287 24055
rect 10100 24024 10287 24052
rect 10100 24012 10106 24024
rect 10275 24021 10287 24024
rect 10321 24021 10333 24055
rect 10275 24015 10333 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2774 23848 2780 23860
rect 2735 23820 2780 23848
rect 2774 23808 2780 23820
rect 2832 23808 2838 23860
rect 6270 23808 6276 23860
rect 6328 23848 6334 23860
rect 6365 23851 6423 23857
rect 6365 23848 6377 23851
rect 6328 23820 6377 23848
rect 6328 23808 6334 23820
rect 6365 23817 6377 23820
rect 6411 23817 6423 23851
rect 6365 23811 6423 23817
rect 6454 23808 6460 23860
rect 6512 23848 6518 23860
rect 7009 23851 7067 23857
rect 7009 23848 7021 23851
rect 6512 23820 7021 23848
rect 6512 23808 6518 23820
rect 7009 23817 7021 23820
rect 7055 23817 7067 23851
rect 8294 23848 8300 23860
rect 8255 23820 8300 23848
rect 7009 23811 7067 23817
rect 8294 23808 8300 23820
rect 8352 23808 8358 23860
rect 10134 23808 10140 23860
rect 10192 23848 10198 23860
rect 10965 23851 11023 23857
rect 10965 23848 10977 23851
rect 10192 23820 10977 23848
rect 10192 23808 10198 23820
rect 10965 23817 10977 23820
rect 11011 23817 11023 23851
rect 10965 23811 11023 23817
rect 14001 23851 14059 23857
rect 14001 23817 14013 23851
rect 14047 23848 14059 23851
rect 15838 23848 15844 23860
rect 14047 23820 15844 23848
rect 14047 23817 14059 23820
rect 14001 23811 14059 23817
rect 15838 23808 15844 23820
rect 15896 23808 15902 23860
rect 19981 23851 20039 23857
rect 19981 23817 19993 23851
rect 20027 23848 20039 23851
rect 21358 23848 21364 23860
rect 20027 23820 21364 23848
rect 20027 23817 20039 23820
rect 19981 23811 20039 23817
rect 934 23740 940 23792
rect 992 23780 998 23792
rect 4617 23783 4675 23789
rect 4617 23780 4629 23783
rect 992 23752 4629 23780
rect 992 23740 998 23752
rect 2292 23647 2350 23653
rect 2292 23613 2304 23647
rect 2338 23644 2350 23647
rect 2774 23644 2780 23656
rect 2338 23616 2780 23644
rect 2338 23613 2350 23616
rect 2292 23607 2350 23613
rect 2774 23604 2780 23616
rect 2832 23604 2838 23656
rect 4239 23653 4267 23752
rect 4617 23749 4629 23752
rect 4663 23749 4675 23783
rect 4617 23743 4675 23749
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23712 7619 23715
rect 8481 23715 8539 23721
rect 8481 23712 8493 23715
rect 7607 23684 8493 23712
rect 7607 23681 7619 23684
rect 7561 23675 7619 23681
rect 8481 23681 8493 23684
rect 8527 23712 8539 23715
rect 8662 23712 8668 23724
rect 8527 23684 8668 23712
rect 8527 23681 8539 23684
rect 8481 23675 8539 23681
rect 8662 23672 8668 23684
rect 8720 23672 8726 23724
rect 4224 23647 4282 23653
rect 4224 23613 4236 23647
rect 4270 23613 4282 23647
rect 6822 23644 6828 23656
rect 6783 23616 6828 23644
rect 4224 23607 4282 23613
rect 6822 23604 6828 23616
rect 6880 23604 6886 23656
rect 9861 23647 9919 23653
rect 9861 23644 9873 23647
rect 9232 23616 9873 23644
rect 7929 23579 7987 23585
rect 7929 23545 7941 23579
rect 7975 23576 7987 23579
rect 8573 23579 8631 23585
rect 8573 23576 8585 23579
rect 7975 23548 8585 23576
rect 7975 23545 7987 23548
rect 7929 23539 7987 23545
rect 8573 23545 8585 23548
rect 8619 23545 8631 23579
rect 9122 23576 9128 23588
rect 9083 23548 9128 23576
rect 8573 23539 8631 23545
rect 2363 23511 2421 23517
rect 2363 23477 2375 23511
rect 2409 23508 2421 23511
rect 2498 23508 2504 23520
rect 2409 23480 2504 23508
rect 2409 23477 2421 23480
rect 2363 23471 2421 23477
rect 2498 23468 2504 23480
rect 2556 23468 2562 23520
rect 4295 23511 4353 23517
rect 4295 23477 4307 23511
rect 4341 23508 4353 23511
rect 4522 23508 4528 23520
rect 4341 23480 4528 23508
rect 4341 23477 4353 23480
rect 4295 23471 4353 23477
rect 4522 23468 4528 23480
rect 4580 23468 4586 23520
rect 8588 23508 8616 23539
rect 9122 23536 9128 23548
rect 9180 23536 9186 23588
rect 8846 23508 8852 23520
rect 8588 23480 8852 23508
rect 8846 23468 8852 23480
rect 8904 23508 8910 23520
rect 9232 23508 9260 23616
rect 9861 23613 9873 23616
rect 9907 23644 9919 23647
rect 10045 23647 10103 23653
rect 10045 23644 10057 23647
rect 9907 23616 10057 23644
rect 9907 23613 9919 23616
rect 9861 23607 9919 23613
rect 10045 23613 10057 23616
rect 10091 23613 10103 23647
rect 10045 23607 10103 23613
rect 12802 23604 12808 23656
rect 12860 23644 12866 23656
rect 13817 23647 13875 23653
rect 13817 23644 13829 23647
rect 12860 23616 13829 23644
rect 12860 23604 12866 23616
rect 13817 23613 13829 23616
rect 13863 23644 13875 23647
rect 14369 23647 14427 23653
rect 14369 23644 14381 23647
rect 13863 23616 14381 23644
rect 13863 23613 13875 23616
rect 13817 23607 13875 23613
rect 14369 23613 14381 23616
rect 14415 23613 14427 23647
rect 14369 23607 14427 23613
rect 18116 23647 18174 23653
rect 18116 23613 18128 23647
rect 18162 23644 18174 23647
rect 18598 23644 18604 23656
rect 18162 23616 18604 23644
rect 18162 23613 18174 23616
rect 18116 23607 18174 23613
rect 18598 23604 18604 23616
rect 18656 23604 18662 23656
rect 19496 23647 19554 23653
rect 19496 23613 19508 23647
rect 19542 23644 19554 23647
rect 19996 23644 20024 23811
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 21913 23851 21971 23857
rect 21913 23817 21925 23851
rect 21959 23848 21971 23851
rect 23290 23848 23296 23860
rect 21959 23820 23296 23848
rect 21959 23817 21971 23820
rect 21913 23811 21971 23817
rect 19542 23616 20024 23644
rect 21428 23647 21486 23653
rect 19542 23613 19554 23616
rect 19496 23607 19554 23613
rect 21428 23613 21440 23647
rect 21474 23644 21486 23647
rect 21928 23644 21956 23811
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 21474 23616 21956 23644
rect 24632 23647 24690 23653
rect 21474 23613 21486 23616
rect 21428 23607 21486 23613
rect 24632 23613 24644 23647
rect 24678 23644 24690 23647
rect 25130 23644 25136 23656
rect 24678 23616 25136 23644
rect 24678 23613 24690 23616
rect 24632 23607 24690 23613
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 9950 23576 9956 23588
rect 9911 23548 9956 23576
rect 9950 23536 9956 23548
rect 10008 23536 10014 23588
rect 21726 23536 21732 23588
rect 21784 23576 21790 23588
rect 24719 23579 24777 23585
rect 24719 23576 24731 23579
rect 21784 23548 24731 23576
rect 21784 23536 21790 23548
rect 24719 23545 24731 23548
rect 24765 23545 24777 23579
rect 24719 23539 24777 23545
rect 8904 23480 9260 23508
rect 8904 23468 8910 23480
rect 17770 23468 17776 23520
rect 17828 23508 17834 23520
rect 18187 23511 18245 23517
rect 18187 23508 18199 23511
rect 17828 23480 18199 23508
rect 17828 23468 17834 23480
rect 18187 23477 18199 23480
rect 18233 23477 18245 23511
rect 18598 23508 18604 23520
rect 18559 23480 18604 23508
rect 18187 23471 18245 23477
rect 18598 23468 18604 23480
rect 18656 23468 18662 23520
rect 18690 23468 18696 23520
rect 18748 23508 18754 23520
rect 19567 23511 19625 23517
rect 19567 23508 19579 23511
rect 18748 23480 19579 23508
rect 18748 23468 18754 23480
rect 19567 23477 19579 23480
rect 19613 23477 19625 23511
rect 19567 23471 19625 23477
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 21499 23511 21557 23517
rect 21499 23508 21511 23511
rect 20036 23480 21511 23508
rect 20036 23468 20042 23480
rect 21499 23477 21511 23480
rect 21545 23477 21557 23511
rect 21499 23471 21557 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 6822 23304 6828 23316
rect 6783 23276 6828 23304
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 5534 23236 5540 23248
rect 5495 23208 5540 23236
rect 5534 23196 5540 23208
rect 5592 23196 5598 23248
rect 8110 23196 8116 23248
rect 8168 23236 8174 23248
rect 8205 23239 8263 23245
rect 8205 23236 8217 23239
rect 8168 23208 8217 23236
rect 8168 23196 8174 23208
rect 8205 23205 8217 23208
rect 8251 23205 8263 23239
rect 8205 23199 8263 23205
rect 9766 23196 9772 23248
rect 9824 23236 9830 23248
rect 9861 23239 9919 23245
rect 9861 23236 9873 23239
rect 9824 23208 9873 23236
rect 9824 23196 9830 23208
rect 9861 23205 9873 23208
rect 9907 23236 9919 23239
rect 9950 23236 9956 23248
rect 9907 23208 9956 23236
rect 9907 23205 9919 23208
rect 9861 23199 9919 23205
rect 9950 23196 9956 23208
rect 10008 23196 10014 23248
rect 1210 23128 1216 23180
rect 1268 23168 1274 23180
rect 1432 23171 1490 23177
rect 1432 23168 1444 23171
rect 1268 23140 1444 23168
rect 1268 23128 1274 23140
rect 1432 23137 1444 23140
rect 1478 23137 1490 23171
rect 1432 23131 1490 23137
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 4522 23060 4528 23112
rect 4580 23100 4586 23112
rect 5442 23100 5448 23112
rect 4580 23072 5448 23100
rect 4580 23060 4586 23072
rect 5442 23060 5448 23072
rect 5500 23060 5506 23112
rect 6089 23103 6147 23109
rect 6089 23069 6101 23103
rect 6135 23100 6147 23103
rect 6270 23100 6276 23112
rect 6135 23072 6276 23100
rect 6135 23069 6147 23072
rect 6089 23063 6147 23069
rect 6270 23060 6276 23072
rect 6328 23060 6334 23112
rect 7009 23103 7067 23109
rect 7009 23069 7021 23103
rect 7055 23100 7067 23103
rect 7834 23100 7840 23112
rect 7055 23072 7840 23100
rect 7055 23069 7067 23072
rect 7009 23063 7067 23069
rect 7834 23060 7840 23072
rect 7892 23100 7898 23112
rect 8113 23103 8171 23109
rect 8113 23100 8125 23103
rect 7892 23072 8125 23100
rect 7892 23060 7898 23072
rect 8113 23069 8125 23072
rect 8159 23069 8171 23103
rect 8754 23100 8760 23112
rect 8715 23072 8760 23100
rect 8113 23063 8171 23069
rect 8754 23060 8760 23072
rect 8812 23060 8818 23112
rect 9769 23103 9827 23109
rect 9769 23069 9781 23103
rect 9815 23100 9827 23103
rect 10134 23100 10140 23112
rect 9815 23072 10140 23100
rect 9815 23069 9827 23072
rect 9769 23063 9827 23069
rect 10134 23060 10140 23072
rect 10192 23100 10198 23112
rect 18690 23100 18696 23112
rect 10192 23072 18696 23100
rect 10192 23060 10198 23072
rect 18690 23060 18696 23072
rect 18748 23060 18754 23112
rect 7558 23032 7564 23044
rect 7471 23004 7564 23032
rect 7558 22992 7564 23004
rect 7616 23032 7622 23044
rect 8772 23032 8800 23060
rect 9122 23032 9128 23044
rect 7616 23004 8800 23032
rect 9035 23004 9128 23032
rect 7616 22992 7622 23004
rect 9122 22992 9128 23004
rect 9180 23032 9186 23044
rect 10321 23035 10379 23041
rect 10321 23032 10333 23035
rect 9180 23004 10333 23032
rect 9180 22992 9186 23004
rect 10321 23001 10333 23004
rect 10367 23001 10379 23035
rect 10321 22995 10379 23001
rect 1535 22967 1593 22973
rect 1535 22933 1547 22967
rect 1581 22964 1593 22967
rect 2314 22964 2320 22976
rect 1581 22936 2320 22964
rect 1581 22933 1593 22936
rect 1535 22927 1593 22933
rect 2314 22924 2320 22936
rect 2372 22924 2378 22976
rect 22186 22924 22192 22976
rect 22244 22964 22250 22976
rect 24719 22967 24777 22973
rect 24719 22964 24731 22967
rect 22244 22936 24731 22964
rect 22244 22924 22250 22936
rect 24719 22933 24731 22936
rect 24765 22933 24777 22967
rect 24719 22927 24777 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1210 22720 1216 22772
rect 1268 22760 1274 22772
rect 1581 22763 1639 22769
rect 1581 22760 1593 22763
rect 1268 22732 1593 22760
rect 1268 22720 1274 22732
rect 1581 22729 1593 22732
rect 1627 22729 1639 22763
rect 9766 22760 9772 22772
rect 9727 22732 9772 22760
rect 1581 22723 1639 22729
rect 9766 22720 9772 22732
rect 9824 22720 9830 22772
rect 10134 22760 10140 22772
rect 10095 22732 10140 22760
rect 10134 22720 10140 22732
rect 10192 22720 10198 22772
rect 12621 22763 12679 22769
rect 12621 22729 12633 22763
rect 12667 22760 12679 22763
rect 17678 22760 17684 22772
rect 12667 22732 17684 22760
rect 12667 22729 12679 22732
rect 12621 22723 12679 22729
rect 17678 22720 17684 22732
rect 17736 22720 17742 22772
rect 24670 22760 24676 22772
rect 24631 22732 24676 22760
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 9122 22692 9128 22704
rect 8588 22664 9128 22692
rect 5534 22584 5540 22636
rect 5592 22624 5598 22636
rect 5905 22627 5963 22633
rect 5905 22624 5917 22627
rect 5592 22596 5917 22624
rect 5592 22584 5598 22596
rect 5905 22593 5917 22596
rect 5951 22624 5963 22627
rect 6181 22627 6239 22633
rect 6181 22624 6193 22627
rect 5951 22596 6193 22624
rect 5951 22593 5963 22596
rect 5905 22587 5963 22593
rect 6181 22593 6193 22596
rect 6227 22593 6239 22627
rect 6181 22587 6239 22593
rect 6270 22584 6276 22636
rect 6328 22624 6334 22636
rect 8588 22633 8616 22664
rect 9122 22652 9128 22664
rect 9180 22652 9186 22704
rect 7193 22627 7251 22633
rect 7193 22624 7205 22627
rect 6328 22596 7205 22624
rect 6328 22584 6334 22596
rect 7193 22593 7205 22596
rect 7239 22593 7251 22627
rect 7193 22587 7251 22593
rect 8573 22627 8631 22633
rect 8573 22593 8585 22627
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 8754 22584 8760 22636
rect 8812 22624 8818 22636
rect 8849 22627 8907 22633
rect 8849 22624 8861 22627
rect 8812 22596 8861 22624
rect 8812 22584 8818 22596
rect 8849 22593 8861 22596
rect 8895 22593 8907 22627
rect 8849 22587 8907 22593
rect 5077 22559 5135 22565
rect 5077 22525 5089 22559
rect 5123 22556 5135 22559
rect 5813 22559 5871 22565
rect 5813 22556 5825 22559
rect 5123 22528 5825 22556
rect 5123 22525 5135 22528
rect 5077 22519 5135 22525
rect 5813 22525 5825 22528
rect 5859 22556 5871 22559
rect 5859 22528 6592 22556
rect 5859 22525 5871 22528
rect 5813 22519 5871 22525
rect 6564 22432 6592 22528
rect 11238 22516 11244 22568
rect 11296 22556 11302 22568
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 11296 22528 12449 22556
rect 11296 22516 11302 22528
rect 12437 22525 12449 22528
rect 12483 22556 12495 22559
rect 12989 22559 13047 22565
rect 12989 22556 13001 22559
rect 12483 22528 13001 22556
rect 12483 22525 12495 22528
rect 12437 22519 12495 22525
rect 12989 22525 13001 22528
rect 13035 22525 13047 22559
rect 12989 22519 13047 22525
rect 6914 22488 6920 22500
rect 6875 22460 6920 22488
rect 6914 22448 6920 22460
rect 6972 22448 6978 22500
rect 7009 22491 7067 22497
rect 7009 22457 7021 22491
rect 7055 22457 7067 22491
rect 7009 22451 7067 22457
rect 8665 22491 8723 22497
rect 8665 22457 8677 22491
rect 8711 22488 8723 22491
rect 8938 22488 8944 22500
rect 8711 22460 8944 22488
rect 8711 22457 8723 22460
rect 8665 22451 8723 22457
rect 6546 22420 6552 22432
rect 6507 22392 6552 22420
rect 6546 22380 6552 22392
rect 6604 22420 6610 22432
rect 7024 22420 7052 22451
rect 8938 22448 8944 22460
rect 8996 22448 9002 22500
rect 8018 22420 8024 22432
rect 6604 22392 7052 22420
rect 7979 22392 8024 22420
rect 6604 22380 6610 22392
rect 8018 22380 8024 22392
rect 8076 22380 8082 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 5442 22216 5448 22228
rect 5403 22188 5448 22216
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 6914 22216 6920 22228
rect 6875 22188 6920 22216
rect 6914 22176 6920 22188
rect 6972 22176 6978 22228
rect 7834 22216 7840 22228
rect 7795 22188 7840 22216
rect 7834 22176 7840 22188
rect 7892 22176 7898 22228
rect 8018 22148 8024 22160
rect 7979 22120 8024 22148
rect 8018 22108 8024 22120
rect 8076 22108 8082 22160
rect 8665 22083 8723 22089
rect 8665 22049 8677 22083
rect 8711 22080 8723 22083
rect 8938 22080 8944 22092
rect 8711 22052 8944 22080
rect 8711 22049 8723 22052
rect 8665 22043 8723 22049
rect 8938 22040 8944 22052
rect 8996 22040 9002 22092
rect 11308 22083 11366 22089
rect 11308 22049 11320 22083
rect 11354 22080 11366 22083
rect 11422 22080 11428 22092
rect 11354 22052 11428 22080
rect 11354 22049 11366 22052
rect 11308 22043 11366 22049
rect 11422 22040 11428 22052
rect 11480 22080 11486 22092
rect 12066 22080 12072 22092
rect 11480 22052 12072 22080
rect 11480 22040 11486 22052
rect 12066 22040 12072 22052
rect 12124 22040 12130 22092
rect 12780 22083 12838 22089
rect 12780 22049 12792 22083
rect 12826 22080 12838 22083
rect 13538 22080 13544 22092
rect 12826 22052 13544 22080
rect 12826 22049 12838 22052
rect 12780 22043 12838 22049
rect 13538 22040 13544 22052
rect 13596 22040 13602 22092
rect 8938 21836 8944 21888
rect 8996 21876 9002 21888
rect 9033 21879 9091 21885
rect 9033 21876 9045 21879
rect 8996 21848 9045 21876
rect 8996 21836 9002 21848
rect 9033 21845 9045 21848
rect 9079 21845 9091 21879
rect 9033 21839 9091 21845
rect 11379 21879 11437 21885
rect 11379 21845 11391 21879
rect 11425 21876 11437 21879
rect 11882 21876 11888 21888
rect 11425 21848 11888 21876
rect 11425 21845 11437 21848
rect 11379 21839 11437 21845
rect 11882 21836 11888 21848
rect 11940 21836 11946 21888
rect 12526 21876 12532 21888
rect 12439 21848 12532 21876
rect 12526 21836 12532 21848
rect 12584 21876 12590 21888
rect 12851 21879 12909 21885
rect 12851 21876 12863 21879
rect 12584 21848 12863 21876
rect 12584 21836 12590 21848
rect 12851 21845 12863 21848
rect 12897 21845 12909 21879
rect 12851 21839 12909 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 11011 21675 11069 21681
rect 11011 21641 11023 21675
rect 11057 21672 11069 21675
rect 11238 21672 11244 21684
rect 11057 21644 11244 21672
rect 11057 21641 11069 21644
rect 11011 21635 11069 21641
rect 11238 21632 11244 21644
rect 11296 21632 11302 21684
rect 11422 21672 11428 21684
rect 11383 21644 11428 21672
rect 11422 21632 11428 21644
rect 11480 21632 11486 21684
rect 13538 21672 13544 21684
rect 13499 21644 13544 21672
rect 13538 21632 13544 21644
rect 13596 21632 13602 21684
rect 12434 21564 12440 21616
rect 12492 21604 12498 21616
rect 12492 21576 12848 21604
rect 12492 21564 12498 21576
rect 12526 21536 12532 21548
rect 12487 21508 12532 21536
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 12820 21545 12848 21576
rect 12805 21539 12863 21545
rect 12805 21505 12817 21539
rect 12851 21505 12863 21539
rect 12805 21499 12863 21505
rect 10778 21428 10784 21480
rect 10836 21468 10842 21480
rect 10940 21471 10998 21477
rect 10940 21468 10952 21471
rect 10836 21440 10952 21468
rect 10836 21428 10842 21440
rect 10940 21437 10952 21440
rect 10986 21468 10998 21471
rect 11701 21471 11759 21477
rect 11701 21468 11713 21471
rect 10986 21440 11713 21468
rect 10986 21437 10998 21440
rect 10940 21431 10998 21437
rect 11701 21437 11713 21440
rect 11747 21437 11759 21471
rect 11701 21431 11759 21437
rect 12253 21403 12311 21409
rect 12253 21369 12265 21403
rect 12299 21400 12311 21403
rect 12618 21400 12624 21412
rect 12299 21372 12624 21400
rect 12299 21369 12311 21372
rect 12253 21363 12311 21369
rect 12618 21360 12624 21372
rect 12676 21360 12682 21412
rect 8113 21335 8171 21341
rect 8113 21301 8125 21335
rect 8159 21332 8171 21335
rect 8938 21332 8944 21344
rect 8159 21304 8944 21332
rect 8159 21301 8171 21304
rect 8113 21295 8171 21301
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 9674 21332 9680 21344
rect 9635 21304 9680 21332
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 11882 21060 11888 21072
rect 11843 21032 11888 21060
rect 11882 21020 11888 21032
rect 11940 21020 11946 21072
rect 11977 21063 12035 21069
rect 11977 21029 11989 21063
rect 12023 21060 12035 21063
rect 12158 21060 12164 21072
rect 12023 21032 12164 21060
rect 12023 21029 12035 21032
rect 11977 21023 12035 21029
rect 12158 21020 12164 21032
rect 12216 21020 12222 21072
rect 7282 20992 7288 21004
rect 7243 20964 7288 20992
rect 7282 20952 7288 20964
rect 7340 20952 7346 21004
rect 10318 20992 10324 21004
rect 10279 20964 10324 20992
rect 10318 20952 10324 20964
rect 10376 20952 10382 21004
rect 12434 20856 12440 20868
rect 12395 20828 12440 20856
rect 12434 20816 12440 20828
rect 12492 20816 12498 20868
rect 7423 20791 7481 20797
rect 7423 20757 7435 20791
rect 7469 20788 7481 20791
rect 8481 20791 8539 20797
rect 8481 20788 8493 20791
rect 7469 20760 8493 20788
rect 7469 20757 7481 20760
rect 7423 20751 7481 20757
rect 8481 20757 8493 20760
rect 8527 20788 8539 20791
rect 8570 20788 8576 20800
rect 8527 20760 8576 20788
rect 8527 20757 8539 20760
rect 8481 20751 8539 20757
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 9950 20788 9956 20800
rect 9911 20760 9956 20788
rect 9950 20748 9956 20760
rect 10008 20748 10014 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 7282 20584 7288 20596
rect 7243 20556 7288 20584
rect 7282 20544 7288 20556
rect 7340 20544 7346 20596
rect 9585 20587 9643 20593
rect 9585 20553 9597 20587
rect 9631 20584 9643 20587
rect 9674 20584 9680 20596
rect 9631 20556 9680 20584
rect 9631 20553 9643 20556
rect 9585 20547 9643 20553
rect 9674 20544 9680 20556
rect 9732 20544 9738 20596
rect 9950 20584 9956 20596
rect 9911 20556 9956 20584
rect 9950 20544 9956 20556
rect 10008 20544 10014 20596
rect 10318 20544 10324 20596
rect 10376 20584 10382 20596
rect 11057 20587 11115 20593
rect 11057 20584 11069 20587
rect 10376 20556 11069 20584
rect 10376 20544 10382 20556
rect 11057 20553 11069 20556
rect 11103 20553 11115 20587
rect 11057 20547 11115 20553
rect 11517 20587 11575 20593
rect 11517 20553 11529 20587
rect 11563 20584 11575 20587
rect 11882 20584 11888 20596
rect 11563 20556 11888 20584
rect 11563 20553 11575 20556
rect 11517 20547 11575 20553
rect 11882 20544 11888 20556
rect 11940 20544 11946 20596
rect 12618 20544 12624 20596
rect 12676 20584 12682 20596
rect 12713 20587 12771 20593
rect 12713 20584 12725 20587
rect 12676 20556 12725 20584
rect 12676 20544 12682 20556
rect 12713 20553 12725 20556
rect 12759 20553 12771 20587
rect 12713 20547 12771 20553
rect 8570 20448 8576 20460
rect 8531 20420 8576 20448
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 9692 20448 9720 20544
rect 10137 20451 10195 20457
rect 10137 20448 10149 20451
rect 9692 20420 10149 20448
rect 10137 20417 10149 20420
rect 10183 20417 10195 20451
rect 10778 20448 10784 20460
rect 10739 20420 10784 20448
rect 10137 20411 10195 20417
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 12529 20383 12587 20389
rect 12529 20380 12541 20383
rect 12176 20352 12541 20380
rect 8389 20315 8447 20321
rect 8389 20281 8401 20315
rect 8435 20312 8447 20315
rect 8662 20312 8668 20324
rect 8435 20284 8668 20312
rect 8435 20281 8447 20284
rect 8389 20275 8447 20281
rect 8662 20272 8668 20284
rect 8720 20272 8726 20324
rect 9214 20312 9220 20324
rect 9175 20284 9220 20312
rect 9214 20272 9220 20284
rect 9272 20272 9278 20324
rect 10229 20315 10287 20321
rect 10229 20281 10241 20315
rect 10275 20281 10287 20315
rect 10229 20275 10287 20281
rect 9950 20204 9956 20256
rect 10008 20244 10014 20256
rect 10244 20244 10272 20275
rect 12176 20256 12204 20352
rect 12529 20349 12541 20352
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 10008 20216 10272 20244
rect 11885 20247 11943 20253
rect 10008 20204 10014 20216
rect 11885 20213 11897 20247
rect 11931 20244 11943 20247
rect 12158 20244 12164 20256
rect 11931 20216 12164 20244
rect 11931 20213 11943 20216
rect 11885 20207 11943 20213
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 5721 20043 5779 20049
rect 5721 20009 5733 20043
rect 5767 20040 5779 20043
rect 6270 20040 6276 20052
rect 5767 20012 6276 20040
rect 5767 20009 5779 20012
rect 5721 20003 5779 20009
rect 4798 19836 4804 19848
rect 4759 19808 4804 19836
rect 4798 19796 4804 19808
rect 4856 19796 4862 19848
rect 5736 19836 5764 20003
rect 6270 20000 6276 20012
rect 6328 20000 6334 20052
rect 13081 20043 13139 20049
rect 8220 20012 10916 20040
rect 5994 19972 6000 19984
rect 5955 19944 6000 19972
rect 5994 19932 6000 19944
rect 6052 19932 6058 19984
rect 8110 19932 8116 19984
rect 8168 19972 8174 19984
rect 8220 19981 8248 20012
rect 8205 19975 8263 19981
rect 8205 19972 8217 19975
rect 8168 19944 8217 19972
rect 8168 19932 8174 19944
rect 8205 19941 8217 19944
rect 8251 19941 8263 19975
rect 8205 19935 8263 19941
rect 9861 19975 9919 19981
rect 9861 19941 9873 19975
rect 9907 19972 9919 19975
rect 10134 19972 10140 19984
rect 9907 19944 10140 19972
rect 9907 19941 9919 19944
rect 9861 19935 9919 19941
rect 10134 19932 10140 19944
rect 10192 19932 10198 19984
rect 10413 19975 10471 19981
rect 10413 19941 10425 19975
rect 10459 19972 10471 19975
rect 10778 19972 10784 19984
rect 10459 19944 10784 19972
rect 10459 19941 10471 19944
rect 10413 19935 10471 19941
rect 10778 19932 10784 19944
rect 10836 19932 10842 19984
rect 10888 19972 10916 20012
rect 13081 20009 13093 20043
rect 13127 20040 13139 20043
rect 13906 20040 13912 20052
rect 13127 20012 13912 20040
rect 13127 20009 13139 20012
rect 13081 20003 13139 20009
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 11241 19975 11299 19981
rect 11241 19972 11253 19975
rect 10888 19944 11253 19972
rect 11241 19941 11253 19944
rect 11287 19941 11299 19975
rect 11241 19935 11299 19941
rect 11330 19904 11336 19916
rect 11291 19876 11336 19904
rect 11330 19864 11336 19876
rect 11388 19864 11394 19916
rect 12894 19904 12900 19916
rect 12855 19876 12900 19904
rect 12894 19864 12900 19876
rect 12952 19864 12958 19916
rect 5905 19839 5963 19845
rect 5905 19836 5917 19839
rect 5736 19808 5917 19836
rect 5905 19805 5917 19808
rect 5951 19805 5963 19839
rect 5905 19799 5963 19805
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19805 6239 19839
rect 6181 19799 6239 19805
rect 8113 19839 8171 19845
rect 8113 19805 8125 19839
rect 8159 19805 8171 19839
rect 8113 19799 8171 19805
rect 8757 19839 8815 19845
rect 8757 19805 8769 19839
rect 8803 19836 8815 19839
rect 9214 19836 9220 19848
rect 8803 19808 9220 19836
rect 8803 19805 8815 19808
rect 8757 19799 8815 19805
rect 5442 19728 5448 19780
rect 5500 19768 5506 19780
rect 6196 19768 6224 19799
rect 5500 19740 6224 19768
rect 5500 19728 5506 19740
rect 7466 19660 7472 19712
rect 7524 19700 7530 19712
rect 7837 19703 7895 19709
rect 7837 19700 7849 19703
rect 7524 19672 7849 19700
rect 7524 19660 7530 19672
rect 7837 19669 7849 19672
rect 7883 19700 7895 19703
rect 8128 19700 8156 19799
rect 9214 19796 9220 19808
rect 9272 19836 9278 19848
rect 9769 19839 9827 19845
rect 9769 19836 9781 19839
rect 9272 19808 9781 19836
rect 9272 19796 9278 19808
rect 9769 19805 9781 19808
rect 9815 19836 9827 19839
rect 10226 19836 10232 19848
rect 9815 19808 10232 19836
rect 9815 19805 9827 19808
rect 9769 19799 9827 19805
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 8662 19728 8668 19780
rect 8720 19768 8726 19780
rect 11330 19768 11336 19780
rect 8720 19740 11336 19768
rect 8720 19728 8726 19740
rect 11330 19728 11336 19740
rect 11388 19728 11394 19780
rect 7883 19672 8156 19700
rect 7883 19669 7895 19672
rect 7837 19663 7895 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 5994 19456 6000 19508
rect 6052 19496 6058 19508
rect 6181 19499 6239 19505
rect 6181 19496 6193 19499
rect 6052 19468 6193 19496
rect 6052 19456 6058 19468
rect 6181 19465 6193 19468
rect 6227 19496 6239 19499
rect 6454 19496 6460 19508
rect 6227 19468 6460 19496
rect 6227 19465 6239 19468
rect 6181 19459 6239 19465
rect 6454 19456 6460 19468
rect 6512 19496 6518 19508
rect 6549 19499 6607 19505
rect 6549 19496 6561 19499
rect 6512 19468 6561 19496
rect 6512 19456 6518 19468
rect 6549 19465 6561 19468
rect 6595 19465 6607 19499
rect 8110 19496 8116 19508
rect 8071 19468 8116 19496
rect 6549 19459 6607 19465
rect 8110 19456 8116 19468
rect 8168 19456 8174 19508
rect 9677 19499 9735 19505
rect 9677 19465 9689 19499
rect 9723 19496 9735 19499
rect 10045 19499 10103 19505
rect 10045 19496 10057 19499
rect 9723 19468 10057 19496
rect 9723 19465 9735 19468
rect 9677 19459 9735 19465
rect 10045 19465 10057 19468
rect 10091 19496 10103 19499
rect 10134 19496 10140 19508
rect 10091 19468 10140 19496
rect 10091 19465 10103 19468
rect 10045 19459 10103 19465
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 10226 19456 10232 19508
rect 10284 19496 10290 19508
rect 10321 19499 10379 19505
rect 10321 19496 10333 19499
rect 10284 19468 10333 19496
rect 10284 19456 10290 19468
rect 10321 19465 10333 19468
rect 10367 19465 10379 19499
rect 11330 19496 11336 19508
rect 11291 19468 11336 19496
rect 10321 19459 10379 19465
rect 11330 19456 11336 19468
rect 11388 19456 11394 19508
rect 14642 19496 14648 19508
rect 14603 19468 14648 19496
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 12575 19431 12633 19437
rect 12575 19397 12587 19431
rect 12621 19428 12633 19431
rect 12894 19428 12900 19440
rect 12621 19400 12900 19428
rect 12621 19397 12633 19400
rect 12575 19391 12633 19397
rect 12894 19388 12900 19400
rect 12952 19428 12958 19440
rect 13265 19431 13323 19437
rect 13265 19428 13277 19431
rect 12952 19400 13277 19428
rect 12952 19388 12958 19400
rect 13265 19397 13277 19400
rect 13311 19397 13323 19431
rect 13265 19391 13323 19397
rect 3970 19320 3976 19372
rect 4028 19360 4034 19372
rect 4798 19360 4804 19372
rect 4028 19332 4804 19360
rect 4028 19320 4034 19332
rect 4798 19320 4804 19332
rect 4856 19360 4862 19372
rect 5261 19363 5319 19369
rect 5261 19360 5273 19363
rect 4856 19332 5273 19360
rect 4856 19320 4862 19332
rect 5261 19329 5273 19332
rect 5307 19329 5319 19363
rect 5261 19323 5319 19329
rect 5442 19320 5448 19372
rect 5500 19360 5506 19372
rect 5537 19363 5595 19369
rect 5537 19360 5549 19363
rect 5500 19332 5549 19360
rect 5500 19320 5506 19332
rect 5537 19329 5549 19332
rect 5583 19329 5595 19363
rect 5537 19323 5595 19329
rect 6454 19252 6460 19304
rect 6512 19292 6518 19304
rect 6917 19295 6975 19301
rect 6917 19292 6929 19295
rect 6512 19264 6929 19292
rect 6512 19252 6518 19264
rect 6917 19261 6929 19264
rect 6963 19261 6975 19295
rect 8754 19292 8760 19304
rect 8715 19264 8760 19292
rect 6917 19255 6975 19261
rect 8754 19252 8760 19264
rect 8812 19252 8818 19304
rect 12504 19295 12562 19301
rect 12504 19261 12516 19295
rect 12550 19292 12562 19295
rect 14160 19295 14218 19301
rect 12550 19264 13032 19292
rect 12550 19261 12562 19264
rect 12504 19255 12562 19261
rect 5353 19227 5411 19233
rect 5353 19193 5365 19227
rect 5399 19193 5411 19227
rect 6825 19227 6883 19233
rect 6825 19224 6837 19227
rect 5353 19187 5411 19193
rect 6012 19196 6837 19224
rect 5077 19159 5135 19165
rect 5077 19125 5089 19159
rect 5123 19156 5135 19159
rect 5368 19156 5396 19187
rect 6012 19156 6040 19196
rect 6825 19193 6837 19196
rect 6871 19193 6883 19227
rect 9078 19227 9136 19233
rect 9078 19224 9090 19227
rect 6825 19187 6883 19193
rect 8588 19196 9090 19224
rect 8588 19168 8616 19196
rect 9078 19193 9090 19196
rect 9124 19193 9136 19227
rect 9078 19187 9136 19193
rect 8570 19156 8576 19168
rect 5123 19128 6040 19156
rect 8531 19128 8576 19156
rect 5123 19125 5135 19128
rect 5077 19119 5135 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 13004 19165 13032 19264
rect 14160 19261 14172 19295
rect 14206 19292 14218 19295
rect 14642 19292 14648 19304
rect 14206 19264 14648 19292
rect 14206 19261 14218 19264
rect 14160 19255 14218 19261
rect 14642 19252 14648 19264
rect 14700 19252 14706 19304
rect 12989 19159 13047 19165
rect 12989 19125 13001 19159
rect 13035 19156 13047 19159
rect 13170 19156 13176 19168
rect 13035 19128 13176 19156
rect 13035 19125 13047 19128
rect 12989 19119 13047 19125
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 14090 19116 14096 19168
rect 14148 19156 14154 19168
rect 14231 19159 14289 19165
rect 14231 19156 14243 19159
rect 14148 19128 14243 19156
rect 14148 19116 14154 19128
rect 14231 19125 14243 19128
rect 14277 19125 14289 19159
rect 14231 19119 14289 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2498 18912 2504 18964
rect 2556 18952 2562 18964
rect 3145 18955 3203 18961
rect 3145 18952 3157 18955
rect 2556 18924 3157 18952
rect 2556 18912 2562 18924
rect 3145 18921 3157 18924
rect 3191 18952 3203 18955
rect 3234 18952 3240 18964
rect 3191 18924 3240 18952
rect 3191 18921 3203 18924
rect 3145 18915 3203 18921
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 4246 18952 4252 18964
rect 4207 18924 4252 18952
rect 4246 18912 4252 18924
rect 4304 18912 4310 18964
rect 6454 18952 6460 18964
rect 6415 18924 6460 18952
rect 6454 18912 6460 18924
rect 6512 18912 6518 18964
rect 8018 18952 8024 18964
rect 7979 18924 8024 18952
rect 8018 18912 8024 18924
rect 8076 18912 8082 18964
rect 12158 18952 12164 18964
rect 12119 18924 12164 18952
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 3970 18844 3976 18896
rect 4028 18884 4034 18896
rect 5169 18887 5227 18893
rect 5169 18884 5181 18887
rect 4028 18856 5181 18884
rect 4028 18844 4034 18856
rect 5169 18853 5181 18856
rect 5215 18853 5227 18887
rect 5169 18847 5227 18853
rect 5899 18887 5957 18893
rect 5899 18853 5911 18887
rect 5945 18884 5957 18887
rect 6086 18884 6092 18896
rect 5945 18856 6092 18884
rect 5945 18853 5957 18856
rect 5899 18847 5957 18853
rect 6086 18844 6092 18856
rect 6144 18844 6150 18896
rect 11603 18887 11661 18893
rect 11603 18853 11615 18887
rect 11649 18884 11661 18887
rect 11698 18884 11704 18896
rect 11649 18856 11704 18884
rect 11649 18853 11661 18856
rect 11603 18847 11661 18853
rect 11698 18844 11704 18856
rect 11756 18844 11762 18896
rect 1464 18819 1522 18825
rect 1464 18785 1476 18819
rect 1510 18816 1522 18819
rect 1946 18816 1952 18828
rect 1510 18788 1952 18816
rect 1510 18785 1522 18788
rect 1464 18779 1522 18785
rect 1946 18776 1952 18788
rect 2004 18776 2010 18828
rect 2409 18819 2467 18825
rect 2409 18785 2421 18819
rect 2455 18816 2467 18819
rect 2498 18816 2504 18828
rect 2455 18788 2504 18816
rect 2455 18785 2467 18788
rect 2409 18779 2467 18785
rect 2498 18776 2504 18788
rect 2556 18776 2562 18828
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 4246 18816 4252 18828
rect 4111 18788 4252 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4246 18776 4252 18788
rect 4304 18776 4310 18828
rect 7558 18776 7564 18828
rect 7616 18816 7622 18828
rect 7745 18819 7803 18825
rect 7745 18816 7757 18819
rect 7616 18788 7757 18816
rect 7616 18776 7622 18788
rect 7745 18785 7757 18788
rect 7791 18785 7803 18819
rect 8202 18816 8208 18828
rect 8163 18788 8208 18816
rect 7745 18779 7803 18785
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 5534 18748 5540 18760
rect 5495 18720 5540 18748
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 10778 18708 10784 18760
rect 10836 18748 10842 18760
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 10836 18720 11253 18748
rect 10836 18708 10842 18720
rect 11241 18717 11253 18720
rect 11287 18717 11299 18751
rect 12986 18748 12992 18760
rect 12947 18720 12992 18748
rect 11241 18711 11299 18717
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 1535 18683 1593 18689
rect 1535 18649 1547 18683
rect 1581 18680 1593 18683
rect 2222 18680 2228 18692
rect 1581 18652 2228 18680
rect 1581 18649 1593 18652
rect 1535 18643 1593 18649
rect 2222 18640 2228 18652
rect 2280 18640 2286 18692
rect 1670 18572 1676 18624
rect 1728 18612 1734 18624
rect 2547 18615 2605 18621
rect 2547 18612 2559 18615
rect 1728 18584 2559 18612
rect 1728 18572 1734 18584
rect 2547 18581 2559 18584
rect 2593 18581 2605 18615
rect 8754 18612 8760 18624
rect 8715 18584 8760 18612
rect 2547 18575 2605 18581
rect 8754 18572 8760 18584
rect 8812 18572 8818 18624
rect 10873 18615 10931 18621
rect 10873 18581 10885 18615
rect 10919 18612 10931 18615
rect 11422 18612 11428 18624
rect 10919 18584 11428 18612
rect 10919 18581 10931 18584
rect 10873 18575 10931 18581
rect 11422 18572 11428 18584
rect 11480 18572 11486 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2498 18408 2504 18420
rect 2411 18380 2504 18408
rect 2498 18368 2504 18380
rect 2556 18408 2562 18420
rect 5442 18408 5448 18420
rect 2556 18380 5448 18408
rect 2556 18368 2562 18380
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 8662 18368 8668 18420
rect 8720 18408 8726 18420
rect 8941 18411 8999 18417
rect 8941 18408 8953 18411
rect 8720 18380 8953 18408
rect 8720 18368 8726 18380
rect 8941 18377 8953 18380
rect 8987 18377 8999 18411
rect 8941 18371 8999 18377
rect 18233 18411 18291 18417
rect 18233 18377 18245 18411
rect 18279 18408 18291 18411
rect 19518 18408 19524 18420
rect 18279 18380 19524 18408
rect 18279 18377 18291 18380
rect 18233 18371 18291 18377
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 4246 18340 4252 18352
rect 4159 18312 4252 18340
rect 4246 18300 4252 18312
rect 4304 18340 4310 18352
rect 12618 18340 12624 18352
rect 4304 18312 12624 18340
rect 4304 18300 4310 18312
rect 12618 18300 12624 18312
rect 12676 18300 12682 18352
rect 3234 18272 3240 18284
rect 3195 18244 3240 18272
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18272 4767 18275
rect 5534 18272 5540 18284
rect 4755 18244 5540 18272
rect 4755 18241 4767 18244
rect 4709 18235 4767 18241
rect 5534 18232 5540 18244
rect 5592 18272 5598 18284
rect 5721 18275 5779 18281
rect 5721 18272 5733 18275
rect 5592 18244 5733 18272
rect 5592 18232 5598 18244
rect 5721 18241 5733 18244
rect 5767 18241 5779 18275
rect 5721 18235 5779 18241
rect 7193 18275 7251 18281
rect 7193 18241 7205 18275
rect 7239 18272 7251 18275
rect 8018 18272 8024 18284
rect 7239 18244 8024 18272
rect 7239 18241 7251 18244
rect 7193 18235 7251 18241
rect 8018 18232 8024 18244
rect 8076 18232 8082 18284
rect 12526 18272 12532 18284
rect 12439 18244 12532 18272
rect 12526 18232 12532 18244
rect 12584 18272 12590 18284
rect 12986 18272 12992 18284
rect 12584 18244 12992 18272
rect 12584 18232 12590 18244
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 1670 18204 1676 18216
rect 1443 18176 1676 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 1670 18164 1676 18176
rect 1728 18164 1734 18216
rect 5077 18207 5135 18213
rect 5077 18173 5089 18207
rect 5123 18204 5135 18207
rect 5166 18204 5172 18216
rect 5123 18176 5172 18204
rect 5123 18173 5135 18176
rect 5077 18167 5135 18173
rect 5166 18164 5172 18176
rect 5224 18164 5230 18216
rect 5629 18207 5687 18213
rect 5629 18173 5641 18207
rect 5675 18204 5687 18207
rect 6178 18204 6184 18216
rect 5675 18176 6184 18204
rect 5675 18173 5687 18176
rect 5629 18167 5687 18173
rect 6178 18164 6184 18176
rect 6236 18164 6242 18216
rect 11422 18204 11428 18216
rect 11383 18176 11428 18204
rect 11422 18164 11428 18176
rect 11480 18164 11486 18216
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 18322 18204 18328 18216
rect 18095 18176 18328 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 18322 18164 18328 18176
rect 18380 18204 18386 18216
rect 23750 18213 23756 18216
rect 18601 18207 18659 18213
rect 18601 18204 18613 18207
rect 18380 18176 18613 18204
rect 18380 18164 18386 18176
rect 18601 18173 18613 18176
rect 18647 18173 18659 18207
rect 23728 18207 23756 18213
rect 23728 18204 23740 18207
rect 23663 18176 23740 18204
rect 18601 18167 18659 18173
rect 23728 18173 23740 18176
rect 23808 18204 23814 18216
rect 24121 18207 24179 18213
rect 24121 18204 24133 18207
rect 23808 18176 24133 18204
rect 23728 18167 23756 18173
rect 23750 18164 23756 18167
rect 23808 18164 23814 18176
rect 24121 18173 24133 18176
rect 24167 18173 24179 18207
rect 24121 18167 24179 18173
rect 3053 18139 3111 18145
rect 3053 18105 3065 18139
rect 3099 18136 3111 18139
rect 3326 18136 3332 18148
rect 3099 18108 3332 18136
rect 3099 18105 3111 18108
rect 3053 18099 3111 18105
rect 3326 18096 3332 18108
rect 3384 18096 3390 18148
rect 3878 18136 3884 18148
rect 3839 18108 3884 18136
rect 3878 18096 3884 18108
rect 3936 18096 3942 18148
rect 8342 18139 8400 18145
rect 8342 18136 8354 18139
rect 7852 18108 8354 18136
rect 106 18028 112 18080
rect 164 18068 170 18080
rect 1581 18071 1639 18077
rect 1581 18068 1593 18071
rect 164 18040 1593 18068
rect 164 18028 170 18040
rect 1581 18037 1593 18040
rect 1627 18037 1639 18071
rect 1581 18031 1639 18037
rect 6086 18028 6092 18080
rect 6144 18068 6150 18080
rect 6181 18071 6239 18077
rect 6181 18068 6193 18071
rect 6144 18040 6193 18068
rect 6144 18028 6150 18040
rect 6181 18037 6193 18040
rect 6227 18037 6239 18071
rect 7558 18068 7564 18080
rect 7519 18040 7564 18068
rect 6181 18031 6239 18037
rect 7558 18028 7564 18040
rect 7616 18028 7622 18080
rect 7742 18028 7748 18080
rect 7800 18068 7806 18080
rect 7852 18077 7880 18108
rect 8342 18105 8354 18108
rect 8388 18136 8400 18139
rect 8570 18136 8576 18148
rect 8388 18108 8576 18136
rect 8388 18105 8400 18108
rect 8342 18099 8400 18105
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 11517 18139 11575 18145
rect 11517 18105 11529 18139
rect 11563 18136 11575 18139
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 11563 18108 12173 18136
rect 11563 18105 11575 18108
rect 11517 18099 11575 18105
rect 12161 18105 12173 18108
rect 12207 18105 12219 18139
rect 12161 18099 12219 18105
rect 12621 18139 12679 18145
rect 12621 18105 12633 18139
rect 12667 18105 12679 18139
rect 13170 18136 13176 18148
rect 13131 18108 13176 18136
rect 12621 18099 12679 18105
rect 7837 18071 7895 18077
rect 7837 18068 7849 18071
rect 7800 18040 7849 18068
rect 7800 18028 7806 18040
rect 7837 18037 7849 18040
rect 7883 18037 7895 18071
rect 7837 18031 7895 18037
rect 10689 18071 10747 18077
rect 10689 18037 10701 18071
rect 10735 18068 10747 18071
rect 10778 18068 10784 18080
rect 10735 18040 10784 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11698 18028 11704 18080
rect 11756 18068 11762 18080
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 11756 18040 11805 18068
rect 11756 18028 11762 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 12176 18068 12204 18099
rect 12636 18068 12664 18099
rect 13170 18096 13176 18108
rect 13228 18096 13234 18148
rect 12176 18040 12664 18068
rect 11793 18031 11851 18037
rect 17494 18028 17500 18080
rect 17552 18068 17558 18080
rect 23799 18071 23857 18077
rect 23799 18068 23811 18071
rect 17552 18040 23811 18068
rect 17552 18028 17558 18040
rect 23799 18037 23811 18040
rect 23845 18037 23857 18071
rect 23799 18031 23857 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1670 17864 1676 17876
rect 1631 17836 1676 17864
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 6546 17864 6552 17876
rect 6507 17836 6552 17864
rect 6546 17824 6552 17836
rect 6604 17824 6610 17876
rect 11422 17824 11428 17876
rect 11480 17864 11486 17876
rect 11793 17867 11851 17873
rect 11793 17864 11805 17867
rect 11480 17836 11805 17864
rect 11480 17824 11486 17836
rect 11793 17833 11805 17836
rect 11839 17833 11851 17867
rect 12526 17864 12532 17876
rect 12487 17836 12532 17864
rect 11793 17827 11851 17833
rect 2222 17756 2228 17808
rect 2280 17796 2286 17808
rect 2501 17799 2559 17805
rect 2501 17796 2513 17799
rect 2280 17768 2513 17796
rect 2280 17756 2286 17768
rect 2501 17765 2513 17768
rect 2547 17765 2559 17799
rect 2501 17759 2559 17765
rect 2590 17756 2596 17808
rect 2648 17796 2654 17808
rect 2648 17768 3188 17796
rect 2648 17756 2654 17768
rect 3160 17728 3188 17768
rect 3326 17756 3332 17808
rect 3384 17796 3390 17808
rect 4065 17799 4123 17805
rect 4065 17796 4077 17799
rect 3384 17768 4077 17796
rect 3384 17756 3390 17768
rect 4065 17765 4077 17768
rect 4111 17765 4123 17799
rect 4065 17759 4123 17765
rect 5534 17756 5540 17808
rect 5592 17796 5598 17808
rect 5950 17799 6008 17805
rect 5950 17796 5962 17799
rect 5592 17768 5962 17796
rect 5592 17756 5598 17768
rect 5950 17765 5962 17768
rect 5996 17796 6008 17799
rect 6086 17796 6092 17808
rect 5996 17768 6092 17796
rect 5996 17765 6008 17768
rect 5950 17759 6008 17765
rect 6086 17756 6092 17768
rect 6144 17756 6150 17808
rect 8754 17796 8760 17808
rect 8715 17768 8760 17796
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 10502 17756 10508 17808
rect 10560 17796 10566 17808
rect 11194 17799 11252 17805
rect 11194 17796 11206 17799
rect 10560 17768 11206 17796
rect 10560 17756 10566 17768
rect 11194 17765 11206 17768
rect 11240 17796 11252 17799
rect 11698 17796 11704 17808
rect 11240 17768 11704 17796
rect 11240 17765 11252 17768
rect 11194 17759 11252 17765
rect 11698 17756 11704 17768
rect 11756 17756 11762 17808
rect 11808 17796 11836 17827
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 14323 17867 14381 17873
rect 14323 17864 14335 17867
rect 12676 17836 14335 17864
rect 12676 17824 12682 17836
rect 14323 17833 14335 17836
rect 14369 17833 14381 17867
rect 18322 17864 18328 17876
rect 18283 17836 18328 17864
rect 14323 17827 14381 17833
rect 18322 17824 18328 17836
rect 18380 17824 18386 17876
rect 12805 17799 12863 17805
rect 12805 17796 12817 17799
rect 11808 17768 12817 17796
rect 12805 17765 12817 17768
rect 12851 17796 12863 17799
rect 13446 17796 13452 17808
rect 12851 17768 13452 17796
rect 12851 17765 12863 17768
rect 12805 17759 12863 17765
rect 13446 17756 13452 17768
rect 13504 17756 13510 17808
rect 4614 17728 4620 17740
rect 3160 17700 4620 17728
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 8018 17728 8024 17740
rect 7979 17700 8024 17728
rect 8018 17688 8024 17700
rect 8076 17688 8082 17740
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17697 8539 17731
rect 8481 17691 8539 17697
rect 14252 17731 14310 17737
rect 14252 17697 14264 17731
rect 14298 17728 14310 17731
rect 14366 17728 14372 17740
rect 14298 17700 14372 17728
rect 14298 17697 14310 17700
rect 14252 17691 14310 17697
rect 3145 17663 3203 17669
rect 3145 17629 3157 17663
rect 3191 17660 3203 17663
rect 3878 17660 3884 17672
rect 3191 17632 3884 17660
rect 3191 17629 3203 17632
rect 3145 17623 3203 17629
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 5629 17663 5687 17669
rect 5629 17629 5641 17663
rect 5675 17660 5687 17663
rect 5994 17660 6000 17672
rect 5675 17632 6000 17660
rect 5675 17629 5687 17632
rect 5629 17623 5687 17629
rect 5994 17620 6000 17632
rect 6052 17620 6058 17672
rect 8202 17660 8208 17672
rect 7760 17632 8208 17660
rect 5261 17527 5319 17533
rect 5261 17493 5273 17527
rect 5307 17524 5319 17527
rect 6178 17524 6184 17536
rect 5307 17496 6184 17524
rect 5307 17493 5319 17496
rect 5261 17487 5319 17493
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 6822 17484 6828 17536
rect 6880 17524 6886 17536
rect 7760 17533 7788 17632
rect 8202 17620 8208 17632
rect 8260 17660 8266 17672
rect 8496 17660 8524 17691
rect 14366 17688 14372 17700
rect 14424 17688 14430 17740
rect 18208 17731 18266 17737
rect 18208 17697 18220 17731
rect 18254 17728 18266 17731
rect 18414 17728 18420 17740
rect 18254 17700 18420 17728
rect 18254 17697 18266 17700
rect 18208 17691 18266 17697
rect 18414 17688 18420 17700
rect 18472 17688 18478 17740
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24670 17728 24676 17740
rect 24627 17700 24676 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 10870 17660 10876 17672
rect 8260 17632 8524 17660
rect 10831 17632 10876 17660
rect 8260 17620 8266 17632
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17660 12771 17663
rect 12894 17660 12900 17672
rect 12759 17632 12900 17660
rect 12759 17629 12771 17632
rect 12713 17623 12771 17629
rect 12894 17620 12900 17632
rect 12952 17620 12958 17672
rect 13170 17660 13176 17672
rect 13131 17632 13176 17660
rect 13170 17620 13176 17632
rect 13228 17620 13234 17672
rect 7745 17527 7803 17533
rect 7745 17524 7757 17527
rect 6880 17496 7757 17524
rect 6880 17484 6886 17496
rect 7745 17493 7757 17496
rect 7791 17493 7803 17527
rect 7745 17487 7803 17493
rect 10502 17484 10508 17536
rect 10560 17524 10566 17536
rect 10597 17527 10655 17533
rect 10597 17524 10609 17527
rect 10560 17496 10609 17524
rect 10560 17484 10566 17496
rect 10597 17493 10609 17496
rect 10643 17493 10655 17527
rect 10597 17487 10655 17493
rect 22278 17484 22284 17536
rect 22336 17524 22342 17536
rect 24719 17527 24777 17533
rect 24719 17524 24731 17527
rect 22336 17496 24731 17524
rect 22336 17484 22342 17496
rect 24719 17493 24731 17496
rect 24765 17493 24777 17527
rect 24719 17487 24777 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2222 17280 2228 17332
rect 2280 17320 2286 17332
rect 2777 17323 2835 17329
rect 2777 17320 2789 17323
rect 2280 17292 2789 17320
rect 2280 17280 2286 17292
rect 2777 17289 2789 17292
rect 2823 17289 2835 17323
rect 4614 17320 4620 17332
rect 4527 17292 4620 17320
rect 2777 17283 2835 17289
rect 4614 17280 4620 17292
rect 4672 17320 4678 17332
rect 4893 17323 4951 17329
rect 4893 17320 4905 17323
rect 4672 17292 4905 17320
rect 4672 17280 4678 17292
rect 4893 17289 4905 17292
rect 4939 17289 4951 17323
rect 5994 17320 6000 17332
rect 5955 17292 6000 17320
rect 4893 17283 4951 17289
rect 5994 17280 6000 17292
rect 6052 17280 6058 17332
rect 8938 17320 8944 17332
rect 8899 17292 8944 17320
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 13446 17320 13452 17332
rect 13407 17292 13452 17320
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 24670 17320 24676 17332
rect 24631 17292 24676 17320
rect 24670 17280 24676 17292
rect 24728 17280 24734 17332
rect 2501 17255 2559 17261
rect 2501 17221 2513 17255
rect 2547 17252 2559 17255
rect 2590 17252 2596 17264
rect 2547 17224 2596 17252
rect 2547 17221 2559 17224
rect 2501 17215 2559 17221
rect 2590 17212 2596 17224
rect 2648 17212 2654 17264
rect 5166 17212 5172 17264
rect 5224 17252 5230 17264
rect 6638 17252 6644 17264
rect 5224 17224 6644 17252
rect 5224 17212 5230 17224
rect 6638 17212 6644 17224
rect 6696 17252 6702 17264
rect 7469 17255 7527 17261
rect 7469 17252 7481 17255
rect 6696 17224 7481 17252
rect 6696 17212 6702 17224
rect 7469 17221 7481 17224
rect 7515 17252 7527 17255
rect 8018 17252 8024 17264
rect 7515 17224 8024 17252
rect 7515 17221 7527 17224
rect 7469 17215 7527 17221
rect 8018 17212 8024 17224
rect 8076 17212 8082 17264
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 11480 17224 13676 17252
rect 11480 17212 11486 17224
rect 10413 17187 10471 17193
rect 10413 17184 10425 17187
rect 9324 17156 10425 17184
rect 3694 17116 3700 17128
rect 3655 17088 3700 17116
rect 3694 17076 3700 17088
rect 3752 17076 3758 17128
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17116 8079 17119
rect 8202 17116 8208 17128
rect 8067 17088 8208 17116
rect 8067 17085 8079 17088
rect 8021 17079 8079 17085
rect 8202 17076 8208 17088
rect 8260 17116 8266 17128
rect 9217 17119 9275 17125
rect 9217 17116 9229 17119
rect 8260 17088 9229 17116
rect 8260 17076 8266 17088
rect 9217 17085 9229 17088
rect 9263 17085 9275 17119
rect 9217 17079 9275 17085
rect 3605 17051 3663 17057
rect 3605 17017 3617 17051
rect 3651 17048 3663 17051
rect 4018 17051 4076 17057
rect 4018 17048 4030 17051
rect 3651 17020 4030 17048
rect 3651 17017 3663 17020
rect 3605 17011 3663 17017
rect 4018 17017 4030 17020
rect 4064 17048 4076 17051
rect 4614 17048 4620 17060
rect 4064 17020 4620 17048
rect 4064 17017 4076 17020
rect 4018 17011 4076 17017
rect 4614 17008 4620 17020
rect 4672 17048 4678 17060
rect 5534 17048 5540 17060
rect 4672 17020 5540 17048
rect 4672 17008 4678 17020
rect 5534 17008 5540 17020
rect 5592 17048 5598 17060
rect 5629 17051 5687 17057
rect 5629 17048 5641 17051
rect 5592 17020 5641 17048
rect 5592 17008 5598 17020
rect 5629 17017 5641 17020
rect 5675 17048 5687 17051
rect 7742 17048 7748 17060
rect 5675 17020 7748 17048
rect 5675 17017 5687 17020
rect 5629 17011 5687 17017
rect 7742 17008 7748 17020
rect 7800 17048 7806 17060
rect 7837 17051 7895 17057
rect 7837 17048 7849 17051
rect 7800 17020 7849 17048
rect 7800 17008 7806 17020
rect 7837 17017 7849 17020
rect 7883 17048 7895 17051
rect 8342 17051 8400 17057
rect 8342 17048 8354 17051
rect 7883 17020 8354 17048
rect 7883 17017 7895 17020
rect 7837 17011 7895 17017
rect 8342 17017 8354 17020
rect 8388 17048 8400 17051
rect 9324 17048 9352 17156
rect 10413 17153 10425 17156
rect 10459 17184 10471 17187
rect 10502 17184 10508 17196
rect 10459 17156 10508 17184
rect 10459 17153 10471 17156
rect 10413 17147 10471 17153
rect 10502 17144 10508 17156
rect 10560 17184 10566 17196
rect 12526 17184 12532 17196
rect 10560 17156 10961 17184
rect 12487 17156 12532 17184
rect 10560 17144 10566 17156
rect 10597 17119 10655 17125
rect 10597 17116 10609 17119
rect 8388 17020 9352 17048
rect 10152 17088 10609 17116
rect 8388 17017 8400 17020
rect 8342 17011 8400 17017
rect 10152 16992 10180 17088
rect 10597 17085 10609 17088
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 10933 17057 10961 17156
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12894 17184 12900 17196
rect 12855 17156 12900 17184
rect 12894 17144 12900 17156
rect 12952 17144 12958 17196
rect 13648 17184 13676 17224
rect 14001 17187 14059 17193
rect 14001 17184 14013 17187
rect 13648 17156 14013 17184
rect 14001 17153 14013 17156
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13786 17088 13921 17116
rect 10918 17051 10976 17057
rect 10918 17017 10930 17051
rect 10964 17017 10976 17051
rect 10918 17011 10976 17017
rect 12621 17051 12679 17057
rect 12621 17017 12633 17051
rect 12667 17017 12679 17051
rect 13786 17048 13814 17088
rect 13909 17085 13921 17088
rect 13955 17116 13967 17119
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13955 17088 14105 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 18046 17048 18052 17060
rect 12621 17011 12679 17017
rect 13280 17020 13814 17048
rect 18007 17020 18052 17048
rect 6822 16940 6828 16992
rect 6880 16980 6886 16992
rect 7101 16983 7159 16989
rect 7101 16980 7113 16983
rect 6880 16952 7113 16980
rect 6880 16940 6886 16952
rect 7101 16949 7113 16952
rect 7147 16949 7159 16983
rect 10134 16980 10140 16992
rect 10095 16952 10140 16980
rect 7101 16943 7159 16949
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 11517 16983 11575 16989
rect 11517 16949 11529 16983
rect 11563 16980 11575 16983
rect 12253 16983 12311 16989
rect 12253 16980 12265 16983
rect 11563 16952 12265 16980
rect 11563 16949 11575 16952
rect 11517 16943 11575 16949
rect 12253 16949 12265 16952
rect 12299 16980 12311 16983
rect 12636 16980 12664 17011
rect 13280 16980 13308 17020
rect 18046 17008 18052 17020
rect 18104 17008 18110 17060
rect 12299 16952 13308 16980
rect 12299 16949 12311 16952
rect 12253 16943 12311 16949
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 15013 16983 15071 16989
rect 15013 16980 15025 16983
rect 14424 16952 15025 16980
rect 14424 16940 14430 16952
rect 15013 16949 15025 16952
rect 15059 16949 15071 16983
rect 17494 16980 17500 16992
rect 17455 16952 17500 16980
rect 15013 16943 15071 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 17865 16983 17923 16989
rect 17865 16949 17877 16983
rect 17911 16980 17923 16983
rect 18156 16980 18184 17079
rect 18230 16980 18236 16992
rect 17911 16952 18236 16980
rect 17911 16949 17923 16952
rect 17865 16943 17923 16949
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 3878 16736 3884 16788
rect 3936 16776 3942 16788
rect 4709 16779 4767 16785
rect 4709 16776 4721 16779
rect 3936 16748 4721 16776
rect 3936 16736 3942 16748
rect 4709 16745 4721 16748
rect 4755 16776 4767 16779
rect 4798 16776 4804 16788
rect 4755 16748 4804 16776
rect 4755 16745 4767 16748
rect 4709 16739 4767 16745
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 5813 16779 5871 16785
rect 5813 16745 5825 16779
rect 5859 16776 5871 16779
rect 5994 16776 6000 16788
rect 5859 16748 6000 16776
rect 5859 16745 5871 16748
rect 5813 16739 5871 16745
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 8846 16776 8852 16788
rect 8803 16748 8852 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 8846 16736 8852 16748
rect 8904 16736 8910 16788
rect 12526 16776 12532 16788
rect 12487 16748 12532 16776
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 7742 16668 7748 16720
rect 7800 16708 7806 16720
rect 8158 16711 8216 16717
rect 8158 16708 8170 16711
rect 7800 16680 8170 16708
rect 7800 16668 7806 16680
rect 8158 16677 8170 16680
rect 8204 16677 8216 16711
rect 8158 16671 8216 16677
rect 10413 16711 10471 16717
rect 10413 16677 10425 16711
rect 10459 16708 10471 16711
rect 10870 16708 10876 16720
rect 10459 16680 10876 16708
rect 10459 16677 10471 16680
rect 10413 16671 10471 16677
rect 10870 16668 10876 16680
rect 10928 16668 10934 16720
rect 11422 16708 11428 16720
rect 11383 16680 11428 16708
rect 11422 16668 11428 16680
rect 11480 16668 11486 16720
rect 13817 16711 13875 16717
rect 13817 16677 13829 16711
rect 13863 16708 13875 16711
rect 13906 16708 13912 16720
rect 13863 16680 13912 16708
rect 13863 16677 13875 16680
rect 13817 16671 13875 16677
rect 13906 16668 13912 16680
rect 13964 16668 13970 16720
rect 14366 16708 14372 16720
rect 14327 16680 14372 16708
rect 14366 16668 14372 16680
rect 14424 16668 14430 16720
rect 17586 16668 17592 16720
rect 17644 16708 17650 16720
rect 17681 16711 17739 16717
rect 17681 16708 17693 16711
rect 17644 16680 17693 16708
rect 17644 16668 17650 16680
rect 17681 16677 17693 16680
rect 17727 16708 17739 16711
rect 18046 16708 18052 16720
rect 17727 16680 18052 16708
rect 17727 16677 17739 16680
rect 17681 16671 17739 16677
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 5534 16640 5540 16652
rect 5495 16612 5540 16640
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 6089 16643 6147 16649
rect 6089 16609 6101 16643
rect 6135 16640 6147 16643
rect 6178 16640 6184 16652
rect 6135 16612 6184 16640
rect 6135 16609 6147 16612
rect 6089 16603 6147 16609
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 9456 16612 9689 16640
rect 9456 16600 9462 16612
rect 9677 16609 9689 16612
rect 9723 16609 9735 16643
rect 10226 16640 10232 16652
rect 10187 16612 10232 16640
rect 9677 16603 9735 16609
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 11977 16643 12035 16649
rect 11977 16609 11989 16643
rect 12023 16640 12035 16643
rect 12805 16643 12863 16649
rect 12805 16640 12817 16643
rect 12023 16612 12817 16640
rect 12023 16609 12035 16612
rect 11977 16603 12035 16609
rect 12805 16609 12817 16612
rect 12851 16640 12863 16643
rect 12894 16640 12900 16652
rect 12851 16612 12900 16640
rect 12851 16609 12863 16612
rect 12805 16603 12863 16609
rect 12894 16600 12900 16612
rect 12952 16600 12958 16652
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16541 7895 16575
rect 7837 16535 7895 16541
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16572 11391 16575
rect 11422 16572 11428 16584
rect 11379 16544 11428 16572
rect 11379 16541 11391 16544
rect 11333 16535 11391 16541
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 3510 16436 3516 16448
rect 3283 16408 3516 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 3510 16396 3516 16408
rect 3568 16396 3574 16448
rect 3694 16436 3700 16448
rect 3655 16408 3700 16436
rect 3694 16396 3700 16408
rect 3752 16396 3758 16448
rect 7745 16439 7803 16445
rect 7745 16405 7757 16439
rect 7791 16436 7803 16439
rect 7852 16436 7880 16535
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 13722 16572 13728 16584
rect 13683 16544 13728 16572
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 17218 16532 17224 16584
rect 17276 16572 17282 16584
rect 17589 16575 17647 16581
rect 17589 16572 17601 16575
rect 17276 16544 17601 16572
rect 17276 16532 17282 16544
rect 17589 16541 17601 16544
rect 17635 16572 17647 16575
rect 19061 16575 19119 16581
rect 19061 16572 19073 16575
rect 17635 16544 19073 16572
rect 17635 16541 17647 16544
rect 17589 16535 17647 16541
rect 19061 16541 19073 16544
rect 19107 16541 19119 16575
rect 19061 16535 19119 16541
rect 17494 16464 17500 16516
rect 17552 16504 17558 16516
rect 18141 16507 18199 16513
rect 18141 16504 18153 16507
rect 17552 16476 18153 16504
rect 17552 16464 17558 16476
rect 18141 16473 18153 16476
rect 18187 16504 18199 16507
rect 18414 16504 18420 16516
rect 18187 16476 18420 16504
rect 18187 16473 18199 16476
rect 18141 16467 18199 16473
rect 18414 16464 18420 16476
rect 18472 16464 18478 16516
rect 7926 16436 7932 16448
rect 7791 16408 7932 16436
rect 7791 16405 7803 16408
rect 7745 16399 7803 16405
rect 7926 16396 7932 16408
rect 7984 16396 7990 16448
rect 14734 16436 14740 16448
rect 14695 16408 14740 16436
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 18230 16396 18236 16448
rect 18288 16436 18294 16448
rect 18509 16439 18567 16445
rect 18509 16436 18521 16439
rect 18288 16408 18521 16436
rect 18288 16396 18294 16408
rect 18509 16405 18521 16408
rect 18555 16405 18567 16439
rect 18509 16399 18567 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 5166 16232 5172 16244
rect 4442 16204 5172 16232
rect 4442 16164 4470 16204
rect 5166 16192 5172 16204
rect 5224 16192 5230 16244
rect 7742 16232 7748 16244
rect 7703 16204 7748 16232
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 11330 16232 11336 16244
rect 11291 16204 11336 16232
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 17218 16232 17224 16244
rect 13780 16192 13814 16232
rect 17179 16204 17224 16232
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 17586 16232 17592 16244
rect 17547 16204 17592 16232
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 25130 16232 25136 16244
rect 25091 16204 25136 16232
rect 25130 16192 25136 16204
rect 25188 16192 25194 16244
rect 6914 16164 6920 16176
rect 3436 16136 4470 16164
rect 4632 16136 6920 16164
rect 3436 16037 3464 16136
rect 3694 16096 3700 16108
rect 3655 16068 3700 16096
rect 3694 16056 3700 16068
rect 3752 16056 3758 16108
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 16028 3111 16031
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 3099 16000 3433 16028
rect 3099 15997 3111 16000
rect 3053 15991 3111 15997
rect 3421 15997 3433 16000
rect 3467 15997 3479 16031
rect 3421 15991 3479 15997
rect 3510 15988 3516 16040
rect 3568 16028 3574 16040
rect 3605 16031 3663 16037
rect 3605 16028 3617 16031
rect 3568 16000 3617 16028
rect 3568 15988 3574 16000
rect 3605 15997 3617 16000
rect 3651 16028 3663 16031
rect 4632 16028 4660 16136
rect 6914 16124 6920 16136
rect 6972 16124 6978 16176
rect 10962 16164 10968 16176
rect 10060 16136 10968 16164
rect 4798 16096 4804 16108
rect 4759 16068 4804 16096
rect 4798 16056 4804 16068
rect 4856 16056 4862 16108
rect 5258 16096 5264 16108
rect 5219 16068 5264 16096
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 7558 16096 7564 16108
rect 5592 16068 7564 16096
rect 5592 16056 5598 16068
rect 7558 16056 7564 16068
rect 7616 16096 7622 16108
rect 8849 16099 8907 16105
rect 8849 16096 8861 16099
rect 7616 16068 8861 16096
rect 7616 16056 7622 16068
rect 8849 16065 8861 16068
rect 8895 16096 8907 16099
rect 10060 16096 10088 16136
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 8895 16068 10088 16096
rect 8895 16065 8907 16068
rect 8849 16059 8907 16065
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 3651 16000 4660 16028
rect 7300 16000 7849 16028
rect 3651 15997 3663 16000
rect 3605 15991 3663 15997
rect 4893 15963 4951 15969
rect 4893 15929 4905 15963
rect 4939 15929 4951 15963
rect 4893 15923 4951 15929
rect 4522 15892 4528 15904
rect 4483 15864 4528 15892
rect 4522 15852 4528 15864
rect 4580 15892 4586 15904
rect 4908 15892 4936 15923
rect 4580 15864 4936 15892
rect 4580 15852 4586 15864
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5534 15892 5540 15904
rect 5224 15864 5540 15892
rect 5224 15852 5230 15864
rect 5534 15852 5540 15864
rect 5592 15892 5598 15904
rect 5721 15895 5779 15901
rect 5721 15892 5733 15895
rect 5592 15864 5733 15892
rect 5592 15852 5598 15864
rect 5721 15861 5733 15864
rect 5767 15861 5779 15895
rect 6178 15892 6184 15904
rect 6139 15864 6184 15892
rect 5721 15855 5779 15861
rect 6178 15852 6184 15864
rect 6236 15852 6242 15904
rect 7190 15852 7196 15904
rect 7248 15892 7254 15904
rect 7300 15901 7328 16000
rect 7837 15997 7849 16000
rect 7883 15997 7895 16031
rect 8386 16028 8392 16040
rect 8347 16000 8392 16028
rect 7837 15991 7895 15997
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 10060 16037 10088 16068
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 10192 16068 10333 16096
rect 10192 16056 10198 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16096 13323 16099
rect 13786 16096 13814 16192
rect 14093 16099 14151 16105
rect 14093 16096 14105 16099
rect 13311 16068 14105 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 14093 16065 14105 16068
rect 14139 16065 14151 16099
rect 14093 16059 14151 16065
rect 14366 16056 14372 16108
rect 14424 16096 14430 16108
rect 14645 16099 14703 16105
rect 14645 16096 14657 16099
rect 14424 16068 14657 16096
rect 14424 16056 14430 16068
rect 14645 16065 14657 16068
rect 14691 16065 14703 16099
rect 18414 16096 18420 16108
rect 18375 16068 18420 16096
rect 14645 16059 14703 16065
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 10045 16031 10103 16037
rect 10045 15997 10057 16031
rect 10091 15997 10103 16031
rect 10226 16028 10232 16040
rect 10139 16000 10232 16028
rect 10045 15991 10103 15997
rect 10226 15988 10232 16000
rect 10284 15988 10290 16040
rect 24648 16031 24706 16037
rect 24648 15997 24660 16031
rect 24694 16028 24706 16031
rect 25130 16028 25136 16040
rect 24694 16000 25136 16028
rect 24694 15997 24706 16000
rect 24648 15991 24706 15997
rect 25130 15988 25136 16000
rect 25188 15988 25194 16040
rect 10244 15960 10272 15988
rect 9232 15932 10272 15960
rect 14369 15963 14427 15969
rect 7285 15895 7343 15901
rect 7285 15892 7297 15895
rect 7248 15864 7297 15892
rect 7248 15852 7254 15864
rect 7285 15861 7297 15864
rect 7331 15861 7343 15895
rect 7926 15892 7932 15904
rect 7887 15864 7932 15892
rect 7285 15855 7343 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 9030 15852 9036 15904
rect 9088 15892 9094 15904
rect 9232 15901 9260 15932
rect 14369 15929 14381 15963
rect 14415 15929 14427 15963
rect 14369 15923 14427 15929
rect 9217 15895 9275 15901
rect 9217 15892 9229 15895
rect 9088 15864 9229 15892
rect 9088 15852 9094 15864
rect 9217 15861 9229 15864
rect 9263 15861 9275 15895
rect 9217 15855 9275 15861
rect 9398 15852 9404 15904
rect 9456 15892 9462 15904
rect 9585 15895 9643 15901
rect 9585 15892 9597 15895
rect 9456 15864 9597 15892
rect 9456 15852 9462 15864
rect 9585 15861 9597 15864
rect 9631 15861 9643 15895
rect 9585 15855 9643 15861
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 11609 15895 11667 15901
rect 11609 15892 11621 15895
rect 11480 15864 11621 15892
rect 11480 15852 11486 15864
rect 11609 15861 11621 15864
rect 11655 15861 11667 15895
rect 11609 15855 11667 15861
rect 13817 15895 13875 15901
rect 13817 15861 13829 15895
rect 13863 15892 13875 15895
rect 13906 15892 13912 15904
rect 13863 15864 13912 15892
rect 13863 15861 13875 15864
rect 13817 15855 13875 15861
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 14384 15892 14412 15923
rect 14458 15920 14464 15972
rect 14516 15960 14522 15972
rect 18141 15963 18199 15969
rect 14516 15932 14561 15960
rect 14516 15920 14522 15932
rect 18141 15929 18153 15963
rect 18187 15929 18199 15963
rect 18141 15923 18199 15929
rect 14734 15892 14740 15904
rect 14384 15864 14740 15892
rect 14734 15852 14740 15864
rect 14792 15892 14798 15904
rect 15102 15892 15108 15904
rect 14792 15864 15108 15892
rect 14792 15852 14798 15864
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 18156 15892 18184 15923
rect 18230 15920 18236 15972
rect 18288 15960 18294 15972
rect 18288 15932 18333 15960
rect 18288 15920 18294 15932
rect 18690 15892 18696 15904
rect 18156 15864 18696 15892
rect 18690 15852 18696 15864
rect 18748 15892 18754 15904
rect 19061 15895 19119 15901
rect 19061 15892 19073 15895
rect 18748 15864 19073 15892
rect 18748 15852 18754 15864
rect 19061 15861 19073 15864
rect 19107 15861 19119 15895
rect 19061 15855 19119 15861
rect 24719 15895 24777 15901
rect 24719 15861 24731 15895
rect 24765 15892 24777 15895
rect 25038 15892 25044 15904
rect 24765 15864 25044 15892
rect 24765 15861 24777 15864
rect 24719 15855 24777 15861
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 6457 15691 6515 15697
rect 6457 15688 6469 15691
rect 5592 15660 6469 15688
rect 5592 15648 5598 15660
rect 6457 15657 6469 15660
rect 6503 15657 6515 15691
rect 8202 15688 8208 15700
rect 8163 15660 8208 15688
rect 6457 15651 6515 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 13906 15688 13912 15700
rect 13867 15660 13912 15688
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 14458 15648 14464 15700
rect 14516 15688 14522 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 14516 15660 14657 15688
rect 14516 15648 14522 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 14645 15651 14703 15657
rect 17129 15691 17187 15697
rect 17129 15657 17141 15691
rect 17175 15688 17187 15691
rect 18230 15688 18236 15700
rect 17175 15660 18236 15688
rect 17175 15657 17187 15660
rect 17129 15651 17187 15657
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 4614 15580 4620 15632
rect 4672 15620 4678 15632
rect 4938 15623 4996 15629
rect 4938 15620 4950 15623
rect 4672 15592 4950 15620
rect 4672 15580 4678 15592
rect 4938 15589 4950 15592
rect 4984 15589 4996 15623
rect 4938 15583 4996 15589
rect 4522 15512 4528 15564
rect 4580 15552 4586 15564
rect 5537 15555 5595 15561
rect 5537 15552 5549 15555
rect 4580 15524 5549 15552
rect 4580 15512 4586 15524
rect 5537 15521 5549 15524
rect 5583 15521 5595 15555
rect 6638 15552 6644 15564
rect 6599 15524 6644 15552
rect 5537 15515 5595 15521
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 6914 15552 6920 15564
rect 6875 15524 6920 15552
rect 6914 15512 6920 15524
rect 6972 15512 6978 15564
rect 8202 15552 8208 15564
rect 8163 15524 8208 15552
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8386 15512 8392 15564
rect 8444 15552 8450 15564
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 8444 15524 8493 15552
rect 8444 15512 8450 15524
rect 8481 15521 8493 15524
rect 8527 15552 8539 15555
rect 8846 15552 8852 15564
rect 8527 15524 8852 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 8846 15512 8852 15524
rect 8904 15512 8910 15564
rect 9030 15512 9036 15564
rect 9088 15552 9094 15564
rect 9861 15555 9919 15561
rect 9861 15552 9873 15555
rect 9088 15524 9873 15552
rect 9088 15512 9094 15524
rect 9861 15521 9873 15524
rect 9907 15521 9919 15555
rect 9861 15515 9919 15521
rect 11584 15555 11642 15561
rect 11584 15521 11596 15555
rect 11630 15552 11642 15555
rect 11790 15552 11796 15564
rect 11630 15524 11796 15552
rect 11630 15521 11642 15524
rect 11584 15515 11642 15521
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 13722 15552 13728 15564
rect 13683 15524 13728 15552
rect 13722 15512 13728 15524
rect 13780 15552 13786 15564
rect 14476 15552 14504 15648
rect 16114 15580 16120 15632
rect 16172 15620 16178 15632
rect 16530 15623 16588 15629
rect 16530 15620 16542 15623
rect 16172 15592 16542 15620
rect 16172 15580 16178 15592
rect 16530 15589 16542 15592
rect 16576 15589 16588 15623
rect 18138 15620 18144 15632
rect 18099 15592 18144 15620
rect 16530 15583 16588 15589
rect 18138 15580 18144 15592
rect 18196 15580 18202 15632
rect 18690 15620 18696 15632
rect 18651 15592 18696 15620
rect 18690 15580 18696 15592
rect 18748 15580 18754 15632
rect 24210 15580 24216 15632
rect 24268 15620 24274 15632
rect 24305 15623 24363 15629
rect 24305 15620 24317 15623
rect 24268 15592 24317 15620
rect 24268 15580 24274 15592
rect 24305 15589 24317 15592
rect 24351 15589 24363 15623
rect 24854 15620 24860 15632
rect 24815 15592 24860 15620
rect 24305 15583 24363 15589
rect 24854 15580 24860 15592
rect 24912 15580 24918 15632
rect 13780 15524 14504 15552
rect 13780 15512 13786 15524
rect 2958 15484 2964 15496
rect 2919 15456 2964 15484
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15484 7895 15487
rect 8404 15484 8432 15512
rect 7883 15456 8432 15484
rect 10505 15487 10563 15493
rect 7883 15453 7895 15456
rect 7837 15447 7895 15453
rect 10505 15453 10517 15487
rect 10551 15484 10563 15487
rect 11330 15484 11336 15496
rect 10551 15456 11336 15484
rect 10551 15453 10563 15456
rect 10505 15447 10563 15453
rect 4632 15416 4660 15447
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 15838 15444 15844 15496
rect 15896 15484 15902 15496
rect 16209 15487 16267 15493
rect 16209 15484 16221 15487
rect 15896 15456 16221 15484
rect 15896 15444 15902 15456
rect 16209 15453 16221 15456
rect 16255 15453 16267 15487
rect 16209 15447 16267 15453
rect 17770 15444 17776 15496
rect 17828 15484 17834 15496
rect 18049 15487 18107 15493
rect 18049 15484 18061 15487
rect 17828 15456 18061 15484
rect 17828 15444 17834 15456
rect 18049 15453 18061 15456
rect 18095 15453 18107 15487
rect 18049 15447 18107 15453
rect 24213 15487 24271 15493
rect 24213 15453 24225 15487
rect 24259 15484 24271 15487
rect 25038 15484 25044 15496
rect 24259 15456 25044 15484
rect 24259 15453 24271 15456
rect 24213 15447 24271 15453
rect 25038 15444 25044 15456
rect 25096 15444 25102 15496
rect 5534 15416 5540 15428
rect 4632 15388 5540 15416
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 7469 15351 7527 15357
rect 7469 15317 7481 15351
rect 7515 15348 7527 15351
rect 7650 15348 7656 15360
rect 7515 15320 7656 15348
rect 7515 15317 7527 15320
rect 7469 15311 7527 15317
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 10318 15348 10324 15360
rect 10279 15320 10324 15348
rect 10318 15308 10324 15320
rect 10376 15308 10382 15360
rect 11655 15351 11713 15357
rect 11655 15317 11667 15351
rect 11701 15348 11713 15351
rect 12434 15348 12440 15360
rect 11701 15320 12440 15348
rect 11701 15317 11713 15320
rect 11655 15311 11713 15317
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 6454 15144 6460 15156
rect 6367 15116 6460 15144
rect 6454 15104 6460 15116
rect 6512 15144 6518 15156
rect 6638 15144 6644 15156
rect 6512 15116 6644 15144
rect 6512 15104 6518 15116
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 8481 15147 8539 15153
rect 8481 15144 8493 15147
rect 8260 15116 8493 15144
rect 8260 15104 8266 15116
rect 8481 15113 8493 15116
rect 8527 15113 8539 15147
rect 8481 15107 8539 15113
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 12897 15147 12955 15153
rect 12897 15144 12909 15147
rect 12860 15116 12909 15144
rect 12860 15104 12866 15116
rect 12897 15113 12909 15116
rect 12943 15113 12955 15147
rect 12897 15107 12955 15113
rect 13173 15147 13231 15153
rect 13173 15113 13185 15147
rect 13219 15144 13231 15147
rect 13722 15144 13728 15156
rect 13219 15116 13728 15144
rect 13219 15113 13231 15116
rect 13173 15107 13231 15113
rect 13722 15104 13728 15116
rect 13780 15144 13786 15156
rect 14553 15147 14611 15153
rect 14553 15144 14565 15147
rect 13780 15116 14565 15144
rect 13780 15104 13786 15116
rect 14553 15113 14565 15116
rect 14599 15113 14611 15147
rect 14553 15107 14611 15113
rect 17770 15104 17776 15156
rect 17828 15144 17834 15156
rect 19061 15147 19119 15153
rect 19061 15144 19073 15147
rect 17828 15116 19073 15144
rect 17828 15104 17834 15116
rect 19061 15113 19073 15116
rect 19107 15113 19119 15147
rect 25038 15144 25044 15156
rect 24999 15116 25044 15144
rect 19061 15107 19119 15113
rect 25038 15104 25044 15116
rect 25096 15104 25102 15156
rect 5905 15079 5963 15085
rect 5905 15076 5917 15079
rect 5000 15048 5917 15076
rect 2958 14968 2964 15020
rect 3016 15008 3022 15020
rect 5000 15017 5028 15048
rect 5905 15045 5917 15048
rect 5951 15045 5963 15079
rect 8110 15076 8116 15088
rect 8071 15048 8116 15076
rect 5905 15039 5963 15045
rect 8110 15036 8116 15048
rect 8168 15036 8174 15088
rect 10042 15036 10048 15088
rect 10100 15076 10106 15088
rect 13449 15079 13507 15085
rect 13449 15076 13461 15079
rect 10100 15048 13461 15076
rect 10100 15036 10106 15048
rect 13449 15045 13461 15048
rect 13495 15045 13507 15079
rect 15933 15079 15991 15085
rect 15933 15076 15945 15079
rect 13449 15039 13507 15045
rect 15488 15048 15945 15076
rect 4985 15011 5043 15017
rect 4985 15008 4997 15011
rect 3016 14980 4997 15008
rect 3016 14968 3022 14980
rect 4985 14977 4997 14980
rect 5031 14977 5043 15011
rect 5258 15008 5264 15020
rect 5219 14980 5264 15008
rect 4985 14971 5043 14977
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 6362 14968 6368 15020
rect 6420 15008 6426 15020
rect 7282 15008 7288 15020
rect 6420 14980 7288 15008
rect 6420 14968 6426 14980
rect 7282 14968 7288 14980
rect 7340 15008 7346 15020
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 7340 14980 7573 15008
rect 7340 14968 7346 14980
rect 7561 14977 7573 14980
rect 7607 14977 7619 15011
rect 8128 15008 8156 15036
rect 10318 15008 10324 15020
rect 8128 14980 10324 15008
rect 7561 14971 7619 14977
rect 10318 14968 10324 14980
rect 10376 14968 10382 15020
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14940 3295 14943
rect 3973 14943 4031 14949
rect 3973 14940 3985 14943
rect 3283 14912 3985 14940
rect 3283 14909 3295 14912
rect 3237 14903 3295 14909
rect 3973 14909 3985 14912
rect 4019 14940 4031 14943
rect 4522 14940 4528 14952
rect 4019 14912 4528 14940
rect 4019 14909 4031 14912
rect 3973 14903 4031 14909
rect 4522 14900 4528 14912
rect 4580 14900 4586 14952
rect 12710 14949 12716 14952
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14940 9275 14943
rect 12253 14943 12311 14949
rect 9263 14912 9628 14940
rect 9263 14909 9275 14912
rect 9217 14903 9275 14909
rect 4062 14872 4068 14884
rect 4023 14844 4068 14872
rect 4062 14832 4068 14844
rect 4120 14832 4126 14884
rect 5074 14832 5080 14884
rect 5132 14872 5138 14884
rect 5132 14844 5177 14872
rect 5132 14832 5138 14844
rect 7650 14832 7656 14884
rect 7708 14872 7714 14884
rect 7708 14844 7753 14872
rect 7708 14832 7714 14844
rect 9600 14816 9628 14912
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12656 14943 12716 14949
rect 12656 14940 12668 14943
rect 12299 14912 12668 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12656 14909 12668 14912
rect 12702 14909 12716 14943
rect 12656 14903 12716 14909
rect 12710 14900 12716 14903
rect 12768 14900 12774 14952
rect 10413 14875 10471 14881
rect 10413 14841 10425 14875
rect 10459 14872 10471 14875
rect 10686 14872 10692 14884
rect 10459 14844 10692 14872
rect 10459 14841 10471 14844
rect 10413 14835 10471 14841
rect 4614 14804 4620 14816
rect 4575 14776 4620 14804
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 6914 14764 6920 14816
rect 6972 14804 6978 14816
rect 7101 14807 7159 14813
rect 7101 14804 7113 14807
rect 6972 14776 7113 14804
rect 6972 14764 6978 14776
rect 7101 14773 7113 14776
rect 7147 14804 7159 14807
rect 8662 14804 8668 14816
rect 7147 14776 8668 14804
rect 7147 14773 7159 14776
rect 7101 14767 7159 14773
rect 8662 14764 8668 14776
rect 8720 14764 8726 14816
rect 8846 14804 8852 14816
rect 8807 14776 8852 14804
rect 8846 14764 8852 14776
rect 8904 14764 8910 14816
rect 9398 14804 9404 14816
rect 9359 14776 9404 14804
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 9582 14764 9588 14816
rect 9640 14804 9646 14816
rect 9677 14807 9735 14813
rect 9677 14804 9689 14807
rect 9640 14776 9689 14804
rect 9640 14764 9646 14776
rect 9677 14773 9689 14776
rect 9723 14773 9735 14807
rect 9677 14767 9735 14773
rect 10137 14807 10195 14813
rect 10137 14773 10149 14807
rect 10183 14804 10195 14807
rect 10428 14804 10456 14835
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 10965 14875 11023 14881
rect 10965 14841 10977 14875
rect 11011 14841 11023 14875
rect 13464 14872 13492 15039
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13814 14940 13820 14952
rect 13679 14912 13820 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13814 14900 13820 14912
rect 13872 14940 13878 14952
rect 14829 14943 14887 14949
rect 14829 14940 14841 14943
rect 13872 14912 14841 14940
rect 13872 14900 13878 14912
rect 14829 14909 14841 14912
rect 14875 14909 14887 14943
rect 14829 14903 14887 14909
rect 13954 14875 14012 14881
rect 13954 14872 13966 14875
rect 13464 14844 13966 14872
rect 10965 14835 11023 14841
rect 13954 14841 13966 14844
rect 14000 14872 14012 14875
rect 15488 14872 15516 15048
rect 15933 15045 15945 15048
rect 15979 15076 15991 15079
rect 16114 15076 16120 15088
rect 15979 15048 16120 15076
rect 15979 15045 15991 15048
rect 15933 15039 15991 15045
rect 16114 15036 16120 15048
rect 16172 15036 16178 15088
rect 18690 15076 18696 15088
rect 18651 15048 18696 15076
rect 18690 15036 18696 15048
rect 18748 15036 18754 15088
rect 15838 14968 15844 15020
rect 15896 15008 15902 15020
rect 17313 15011 17371 15017
rect 17313 15008 17325 15011
rect 15896 14980 17325 15008
rect 15896 14968 15902 14980
rect 17313 14977 17325 14980
rect 17359 14977 17371 15011
rect 19429 15011 19487 15017
rect 19429 15008 19441 15011
rect 17313 14971 17371 14977
rect 17972 14980 19441 15008
rect 16117 14943 16175 14949
rect 16117 14940 16129 14943
rect 14000 14844 15516 14872
rect 15580 14912 16129 14940
rect 14000 14841 14012 14844
rect 13954 14835 14012 14841
rect 10183 14776 10456 14804
rect 10980 14804 11008 14835
rect 15580 14816 15608 14912
rect 16117 14909 16129 14912
rect 16163 14909 16175 14943
rect 16117 14903 16175 14909
rect 16206 14832 16212 14884
rect 16264 14872 16270 14884
rect 16438 14875 16496 14881
rect 16438 14872 16450 14875
rect 16264 14844 16450 14872
rect 16264 14832 16270 14844
rect 16438 14841 16450 14844
rect 16484 14841 16496 14875
rect 16438 14835 16496 14841
rect 16574 14832 16580 14884
rect 16632 14872 16638 14884
rect 17972 14872 18000 14980
rect 19429 14977 19441 14980
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 24210 14968 24216 15020
rect 24268 15008 24274 15020
rect 24397 15011 24455 15017
rect 24397 15008 24409 15011
rect 24268 14980 24409 15008
rect 24268 14968 24274 14980
rect 24397 14977 24409 14980
rect 24443 15008 24455 15011
rect 24673 15011 24731 15017
rect 24673 15008 24685 15011
rect 24443 14980 24685 15008
rect 24443 14977 24455 14980
rect 24397 14971 24455 14977
rect 24673 14977 24685 14980
rect 24719 14977 24731 15011
rect 24673 14971 24731 14977
rect 23477 14943 23535 14949
rect 23477 14909 23489 14943
rect 23523 14940 23535 14943
rect 24026 14940 24032 14952
rect 23523 14912 24032 14940
rect 23523 14909 23535 14912
rect 23477 14903 23535 14909
rect 24026 14900 24032 14912
rect 24084 14900 24090 14952
rect 18141 14875 18199 14881
rect 18141 14872 18153 14875
rect 16632 14844 18153 14872
rect 16632 14832 16638 14844
rect 18141 14841 18153 14844
rect 18187 14841 18199 14875
rect 18141 14835 18199 14841
rect 18230 14832 18236 14884
rect 18288 14872 18294 14884
rect 18288 14844 18333 14872
rect 18288 14832 18294 14844
rect 11609 14807 11667 14813
rect 11609 14804 11621 14807
rect 10980 14776 11621 14804
rect 10183 14773 10195 14776
rect 10137 14767 10195 14773
rect 11609 14773 11621 14776
rect 11655 14804 11667 14807
rect 11790 14804 11796 14816
rect 11655 14776 11796 14804
rect 11655 14773 11667 14776
rect 11609 14767 11667 14773
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 15562 14804 15568 14816
rect 15523 14776 15568 14804
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 17034 14804 17040 14816
rect 16995 14776 17040 14804
rect 17034 14764 17040 14776
rect 17092 14764 17098 14816
rect 17865 14807 17923 14813
rect 17865 14773 17877 14807
rect 17911 14804 17923 14807
rect 18248 14804 18276 14832
rect 17911 14776 18276 14804
rect 17911 14773 17923 14776
rect 17865 14767 17923 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 5074 14600 5080 14612
rect 4120 14572 5080 14600
rect 4120 14560 4126 14572
rect 5074 14560 5080 14572
rect 5132 14560 5138 14612
rect 5534 14600 5540 14612
rect 5495 14572 5540 14600
rect 5534 14560 5540 14572
rect 5592 14560 5598 14612
rect 7650 14600 7656 14612
rect 6012 14572 7656 14600
rect 6012 14476 6040 14572
rect 7650 14560 7656 14572
rect 7708 14600 7714 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 7708 14572 8401 14600
rect 7708 14560 7714 14572
rect 8389 14569 8401 14572
rect 8435 14569 8447 14603
rect 12434 14600 12440 14612
rect 12395 14572 12440 14600
rect 8389 14563 8447 14569
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 16114 14600 16120 14612
rect 13872 14572 13952 14600
rect 16075 14572 16120 14600
rect 13872 14560 13878 14572
rect 7282 14532 7288 14544
rect 7243 14504 7288 14532
rect 7282 14492 7288 14504
rect 7340 14492 7346 14544
rect 7742 14532 7748 14544
rect 7703 14504 7748 14532
rect 7742 14492 7748 14504
rect 7800 14532 7806 14544
rect 10042 14541 10048 14544
rect 9998 14535 10048 14541
rect 9998 14532 10010 14535
rect 7800 14504 10010 14532
rect 7800 14492 7806 14504
rect 9998 14501 10010 14504
rect 10044 14501 10048 14535
rect 9998 14495 10048 14501
rect 10042 14492 10048 14495
rect 10100 14492 10106 14544
rect 11606 14532 11612 14544
rect 11567 14504 11612 14532
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 13924 14541 13952 14572
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 17034 14560 17040 14612
rect 17092 14600 17098 14612
rect 17957 14603 18015 14609
rect 17957 14600 17969 14603
rect 17092 14572 17969 14600
rect 17092 14560 17098 14572
rect 17957 14569 17969 14572
rect 18003 14600 18015 14603
rect 18138 14600 18144 14612
rect 18003 14572 18144 14600
rect 18003 14569 18015 14572
rect 17957 14563 18015 14569
rect 18138 14560 18144 14572
rect 18196 14600 18202 14612
rect 18196 14572 18460 14600
rect 18196 14560 18202 14572
rect 13909 14535 13967 14541
rect 13909 14501 13921 14535
rect 13955 14501 13967 14535
rect 16132 14532 16160 14560
rect 16666 14532 16672 14544
rect 16132 14504 16672 14532
rect 13909 14495 13967 14501
rect 16666 14492 16672 14504
rect 16724 14532 16730 14544
rect 16898 14535 16956 14541
rect 16898 14532 16910 14535
rect 16724 14504 16910 14532
rect 16724 14492 16730 14504
rect 16898 14501 16910 14504
rect 16944 14501 16956 14535
rect 16898 14495 16956 14501
rect 18230 14492 18236 14544
rect 18288 14532 18294 14544
rect 18325 14535 18383 14541
rect 18325 14532 18337 14535
rect 18288 14504 18337 14532
rect 18288 14492 18294 14504
rect 18325 14501 18337 14504
rect 18371 14501 18383 14535
rect 18325 14495 18383 14501
rect 18432 14476 18460 14572
rect 24118 14492 24124 14544
rect 24176 14532 24182 14544
rect 24213 14535 24271 14541
rect 24213 14532 24225 14535
rect 24176 14504 24225 14532
rect 24176 14492 24182 14504
rect 24213 14501 24225 14504
rect 24259 14501 24271 14535
rect 24213 14495 24271 14501
rect 24765 14535 24823 14541
rect 24765 14501 24777 14535
rect 24811 14532 24823 14535
rect 24854 14532 24860 14544
rect 24811 14504 24860 14532
rect 24811 14501 24823 14504
rect 24765 14495 24823 14501
rect 24854 14492 24860 14504
rect 24912 14492 24918 14544
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 4709 14467 4767 14473
rect 4709 14433 4721 14467
rect 4755 14464 4767 14467
rect 4982 14464 4988 14476
rect 4755 14436 4988 14464
rect 4755 14433 4767 14436
rect 4709 14427 4767 14433
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 5994 14464 6000 14476
rect 5955 14436 6000 14464
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6641 14467 6699 14473
rect 6641 14433 6653 14467
rect 6687 14464 6699 14467
rect 7650 14464 7656 14476
rect 6687 14436 7656 14464
rect 6687 14433 6699 14436
rect 6641 14427 6699 14433
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 13078 14424 13084 14476
rect 13136 14464 13142 14476
rect 13173 14467 13231 14473
rect 13173 14464 13185 14467
rect 13136 14436 13185 14464
rect 13136 14424 13142 14436
rect 13173 14433 13185 14436
rect 13219 14433 13231 14467
rect 13173 14427 13231 14433
rect 13725 14467 13783 14473
rect 13725 14433 13737 14467
rect 13771 14464 13783 14467
rect 13814 14464 13820 14476
rect 13771 14436 13820 14464
rect 13771 14433 13783 14436
rect 13725 14427 13783 14433
rect 13814 14424 13820 14436
rect 13872 14464 13878 14476
rect 14185 14467 14243 14473
rect 14185 14464 14197 14467
rect 13872 14436 14197 14464
rect 13872 14424 13878 14436
rect 14185 14433 14197 14436
rect 14231 14433 14243 14467
rect 18414 14464 18420 14476
rect 18327 14436 18420 14464
rect 14185 14427 14243 14433
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14396 7527 14399
rect 7834 14396 7840 14408
rect 7515 14368 7840 14396
rect 7515 14365 7527 14368
rect 7469 14359 7527 14365
rect 7834 14356 7840 14368
rect 7892 14356 7898 14408
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 9858 14396 9864 14408
rect 9723 14368 9864 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 11330 14356 11336 14408
rect 11388 14396 11394 14408
rect 11517 14399 11575 14405
rect 11517 14396 11529 14399
rect 11388 14368 11529 14396
rect 11388 14356 11394 14368
rect 11517 14365 11529 14368
rect 11563 14365 11575 14399
rect 11790 14396 11796 14408
rect 11751 14368 11796 14396
rect 11517 14359 11575 14365
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 16482 14356 16488 14408
rect 16540 14396 16546 14408
rect 16577 14399 16635 14405
rect 16577 14396 16589 14399
rect 16540 14368 16589 14396
rect 16540 14356 16546 14368
rect 16577 14365 16589 14368
rect 16623 14365 16635 14399
rect 16577 14359 16635 14365
rect 24121 14399 24179 14405
rect 24121 14365 24133 14399
rect 24167 14396 24179 14399
rect 24854 14396 24860 14408
rect 24167 14368 24860 14396
rect 24167 14365 24179 14368
rect 24121 14359 24179 14365
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 4338 14260 4344 14272
rect 4299 14232 4344 14260
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 8386 14220 8392 14272
rect 8444 14260 8450 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8444 14232 9045 14260
rect 8444 14220 8450 14232
rect 9033 14229 9045 14232
rect 9079 14260 9091 14263
rect 9490 14260 9496 14272
rect 9079 14232 9496 14260
rect 9079 14229 9091 14232
rect 9033 14223 9091 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 10594 14260 10600 14272
rect 10555 14232 10600 14260
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 15470 14260 15476 14272
rect 15431 14232 15476 14260
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 17494 14260 17500 14272
rect 17455 14232 17500 14260
rect 17494 14220 17500 14232
rect 17552 14220 17558 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 1673 14059 1731 14065
rect 1673 14056 1685 14059
rect 1452 14028 1685 14056
rect 1452 14016 1458 14028
rect 1673 14025 1685 14028
rect 1719 14056 1731 14059
rect 2915 14059 2973 14065
rect 2915 14056 2927 14059
rect 1719 14028 2927 14056
rect 1719 14025 1731 14028
rect 1673 14019 1731 14025
rect 2915 14025 2927 14028
rect 2961 14025 2973 14059
rect 5994 14056 6000 14068
rect 5955 14028 6000 14056
rect 2915 14019 2973 14025
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 8849 14059 8907 14065
rect 8849 14056 8861 14059
rect 8260 14028 8861 14056
rect 8260 14016 8266 14028
rect 8849 14025 8861 14028
rect 8895 14025 8907 14059
rect 10042 14056 10048 14068
rect 10003 14028 10048 14056
rect 8849 14019 8907 14025
rect 6641 13991 6699 13997
rect 6641 13957 6653 13991
rect 6687 13988 6699 13991
rect 7834 13988 7840 14000
rect 6687 13960 7840 13988
rect 6687 13957 6699 13960
rect 6641 13951 6699 13957
rect 7834 13948 7840 13960
rect 7892 13948 7898 14000
rect 8110 13988 8116 14000
rect 8071 13960 8116 13988
rect 8110 13948 8116 13960
rect 8168 13948 8174 14000
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 4430 13920 4436 13932
rect 2731 13892 4436 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 2827 13861 2855 13892
rect 4430 13880 4436 13892
rect 4488 13920 4494 13932
rect 4617 13923 4675 13929
rect 4617 13920 4629 13923
rect 4488 13892 4629 13920
rect 4488 13880 4494 13892
rect 4617 13889 4629 13892
rect 4663 13889 4675 13923
rect 4617 13883 4675 13889
rect 2812 13855 2870 13861
rect 2812 13852 2824 13855
rect 2790 13824 2824 13852
rect 2812 13821 2824 13824
rect 2858 13821 2870 13855
rect 8864 13852 8892 14019
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 11330 14016 11336 14068
rect 11388 14056 11394 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11388 14028 11989 14056
rect 11388 14016 11394 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 16666 14056 16672 14068
rect 16627 14028 16672 14056
rect 11977 14019 12035 14025
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 18414 14056 18420 14068
rect 18375 14028 18420 14056
rect 18414 14016 18420 14028
rect 18472 14016 18478 14068
rect 11333 13923 11391 13929
rect 11333 13889 11345 13923
rect 11379 13920 11391 13923
rect 11606 13920 11612 13932
rect 11379 13892 11612 13920
rect 11379 13889 11391 13892
rect 11333 13883 11391 13889
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 13170 13880 13176 13932
rect 13228 13920 13234 13932
rect 13814 13920 13820 13932
rect 13228 13892 13820 13920
rect 13228 13880 13234 13892
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 14277 13923 14335 13929
rect 14277 13889 14289 13923
rect 14323 13920 14335 13923
rect 16482 13920 16488 13932
rect 14323 13892 16488 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 16482 13880 16488 13892
rect 16540 13920 16546 13932
rect 16945 13923 17003 13929
rect 16945 13920 16957 13923
rect 16540 13892 16957 13920
rect 16540 13880 16546 13892
rect 16945 13889 16957 13892
rect 16991 13889 17003 13923
rect 16945 13883 17003 13889
rect 9033 13855 9091 13861
rect 9033 13852 9045 13855
rect 8864 13824 9045 13852
rect 2812 13815 2870 13821
rect 9033 13821 9045 13824
rect 9079 13852 9091 13855
rect 9306 13852 9312 13864
rect 9079 13824 9312 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 9548 13824 9597 13852
rect 9548 13812 9554 13824
rect 9585 13821 9597 13824
rect 9631 13821 9643 13855
rect 9585 13815 9643 13821
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 10594 13852 10600 13864
rect 10551 13824 10600 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 10594 13812 10600 13824
rect 10652 13852 10658 13864
rect 10689 13855 10747 13861
rect 10689 13852 10701 13855
rect 10652 13824 10701 13852
rect 10652 13812 10658 13824
rect 10689 13821 10701 13824
rect 10735 13821 10747 13855
rect 12434 13852 12440 13864
rect 12395 13824 12440 13852
rect 10689 13815 10747 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 13538 13852 13544 13864
rect 13451 13824 13544 13852
rect 13538 13812 13544 13824
rect 13596 13852 13602 13864
rect 13832 13852 13860 13880
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 13596 13824 13621 13852
rect 13832 13824 14013 13852
rect 13596 13812 13602 13824
rect 14001 13821 14013 13824
rect 14047 13821 14059 13855
rect 15105 13855 15163 13861
rect 15105 13852 15117 13855
rect 14001 13815 14059 13821
rect 14936 13824 15117 13852
rect 3421 13787 3479 13793
rect 3421 13753 3433 13787
rect 3467 13784 3479 13787
rect 4062 13784 4068 13796
rect 3467 13756 4068 13784
rect 3467 13753 3479 13756
rect 3421 13747 3479 13753
rect 4062 13744 4068 13756
rect 4120 13784 4126 13796
rect 4341 13787 4399 13793
rect 4341 13784 4353 13787
rect 4120 13756 4353 13784
rect 4120 13744 4126 13756
rect 4341 13753 4353 13756
rect 4387 13753 4399 13787
rect 4341 13747 4399 13753
rect 4433 13787 4491 13793
rect 4433 13753 4445 13787
rect 4479 13784 4491 13787
rect 4982 13784 4988 13796
rect 4479 13756 4988 13784
rect 4479 13753 4491 13756
rect 4433 13747 4491 13753
rect 3789 13719 3847 13725
rect 3789 13685 3801 13719
rect 3835 13716 3847 13719
rect 4157 13719 4215 13725
rect 4157 13716 4169 13719
rect 3835 13688 4169 13716
rect 3835 13685 3847 13688
rect 3789 13679 3847 13685
rect 4157 13685 4169 13688
rect 4203 13716 4215 13719
rect 4448 13716 4476 13747
rect 4982 13744 4988 13756
rect 5040 13744 5046 13796
rect 7285 13787 7343 13793
rect 7285 13784 7297 13787
rect 7024 13756 7297 13784
rect 4203 13688 4476 13716
rect 4203 13685 4215 13688
rect 4157 13679 4215 13685
rect 4614 13676 4620 13728
rect 4672 13716 4678 13728
rect 7024 13716 7052 13756
rect 7285 13753 7297 13756
rect 7331 13753 7343 13787
rect 7285 13747 7343 13753
rect 7374 13744 7380 13796
rect 7432 13784 7438 13796
rect 7561 13787 7619 13793
rect 7561 13784 7573 13787
rect 7432 13756 7573 13784
rect 7432 13744 7438 13756
rect 7561 13753 7573 13756
rect 7607 13753 7619 13787
rect 7561 13747 7619 13753
rect 4672 13688 7052 13716
rect 7576 13716 7604 13747
rect 7650 13744 7656 13796
rect 7708 13784 7714 13796
rect 9769 13787 9827 13793
rect 7708 13756 7753 13784
rect 7708 13744 7714 13756
rect 9769 13753 9781 13787
rect 9815 13784 9827 13787
rect 9858 13784 9864 13796
rect 9815 13756 9864 13784
rect 9815 13753 9827 13756
rect 9769 13747 9827 13753
rect 9858 13744 9864 13756
rect 9916 13744 9922 13796
rect 13556 13784 13584 13812
rect 14366 13784 14372 13796
rect 13556 13756 14372 13784
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 8481 13719 8539 13725
rect 8481 13716 8493 13719
rect 7576 13688 8493 13716
rect 4672 13676 4678 13688
rect 8481 13685 8493 13688
rect 8527 13685 8539 13719
rect 12618 13716 12624 13728
rect 12579 13688 12624 13716
rect 8481 13679 8539 13685
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 13078 13676 13084 13728
rect 13136 13716 13142 13728
rect 13173 13719 13231 13725
rect 13173 13716 13185 13719
rect 13136 13688 13185 13716
rect 13136 13676 13142 13688
rect 13173 13685 13185 13688
rect 13219 13716 13231 13719
rect 14826 13716 14832 13728
rect 13219 13688 14832 13716
rect 13219 13685 13231 13688
rect 13173 13679 13231 13685
rect 14826 13676 14832 13688
rect 14884 13716 14890 13728
rect 14936 13725 14964 13824
rect 15105 13821 15117 13824
rect 15151 13821 15163 13855
rect 15105 13815 15163 13821
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 15565 13855 15623 13861
rect 15565 13852 15577 13855
rect 15528 13824 15577 13852
rect 15528 13812 15534 13824
rect 15565 13821 15577 13824
rect 15611 13852 15623 13855
rect 15654 13852 15660 13864
rect 15611 13824 15660 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 15838 13852 15844 13864
rect 15799 13824 15844 13852
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 14921 13719 14979 13725
rect 14921 13716 14933 13719
rect 14884 13688 14933 13716
rect 14884 13676 14890 13688
rect 14921 13685 14933 13688
rect 14967 13685 14979 13719
rect 24026 13716 24032 13728
rect 23987 13688 24032 13716
rect 14921 13679 14979 13685
rect 24026 13676 24032 13688
rect 24084 13676 24090 13728
rect 24489 13719 24547 13725
rect 24489 13685 24501 13719
rect 24535 13716 24547 13719
rect 24854 13716 24860 13728
rect 24535 13688 24860 13716
rect 24535 13685 24547 13688
rect 24489 13679 24547 13685
rect 24854 13676 24860 13688
rect 24912 13676 24918 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 7561 13515 7619 13521
rect 7561 13481 7573 13515
rect 7607 13512 7619 13515
rect 7650 13512 7656 13524
rect 7607 13484 7656 13512
rect 7607 13481 7619 13484
rect 7561 13475 7619 13481
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 7834 13512 7840 13524
rect 7795 13484 7840 13512
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 9858 13512 9864 13524
rect 9819 13484 9864 13512
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 13538 13512 13544 13524
rect 9968 13484 13544 13512
rect 4249 13447 4307 13453
rect 4249 13413 4261 13447
rect 4295 13444 4307 13447
rect 4338 13444 4344 13456
rect 4295 13416 4344 13444
rect 4295 13413 4307 13416
rect 4249 13407 4307 13413
rect 4338 13404 4344 13416
rect 4396 13404 4402 13456
rect 7190 13444 7196 13456
rect 7103 13416 7196 13444
rect 7190 13404 7196 13416
rect 7248 13444 7254 13456
rect 9968 13444 9996 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 15562 13512 15568 13524
rect 15523 13484 15568 13512
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 7248 13416 9996 13444
rect 11149 13447 11207 13453
rect 7248 13404 7254 13416
rect 6270 13376 6276 13388
rect 6231 13348 6276 13376
rect 6270 13336 6276 13348
rect 6328 13336 6334 13388
rect 8036 13385 8064 13416
rect 11149 13413 11161 13447
rect 11195 13444 11207 13447
rect 11882 13444 11888 13456
rect 11195 13416 11888 13444
rect 11195 13413 11207 13416
rect 11149 13407 11207 13413
rect 11882 13404 11888 13416
rect 11940 13444 11946 13456
rect 12161 13447 12219 13453
rect 12161 13444 12173 13447
rect 11940 13416 12173 13444
rect 11940 13404 11946 13416
rect 12161 13413 12173 13416
rect 12207 13413 12219 13447
rect 12710 13444 12716 13456
rect 12671 13416 12716 13444
rect 12161 13407 12219 13413
rect 12710 13404 12716 13416
rect 12768 13404 12774 13456
rect 8021 13379 8079 13385
rect 8021 13376 8033 13379
rect 7999 13348 8033 13376
rect 8021 13345 8033 13348
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 8297 13379 8355 13385
rect 8297 13345 8309 13379
rect 8343 13376 8355 13379
rect 8386 13376 8392 13388
rect 8343 13348 8392 13376
rect 8343 13345 8355 13348
rect 8297 13339 8355 13345
rect 8386 13336 8392 13348
rect 8444 13336 8450 13388
rect 11054 13376 11060 13388
rect 11015 13348 11060 13376
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 13630 13376 13636 13388
rect 13591 13348 13636 13376
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 14366 13336 14372 13388
rect 14424 13376 14430 13388
rect 15286 13376 15292 13388
rect 14424 13348 15292 13376
rect 14424 13336 14430 13348
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15654 13336 15660 13388
rect 15712 13376 15718 13388
rect 15749 13379 15807 13385
rect 15749 13376 15761 13379
rect 15712 13348 15761 13376
rect 15712 13336 15718 13348
rect 15749 13345 15761 13348
rect 15795 13345 15807 13379
rect 15749 13339 15807 13345
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13308 3019 13311
rect 4154 13308 4160 13320
rect 3007 13280 4160 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 4154 13268 4160 13280
rect 4212 13308 4218 13320
rect 4430 13308 4436 13320
rect 4212 13280 4257 13308
rect 4391 13280 4436 13308
rect 4212 13268 4218 13280
rect 4430 13268 4436 13280
rect 4488 13268 4494 13320
rect 6730 13308 6736 13320
rect 6691 13280 6736 13308
rect 6730 13268 6736 13280
rect 6788 13268 6794 13320
rect 12066 13308 12072 13320
rect 12027 13280 12072 13308
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 9306 13200 9312 13252
rect 9364 13240 9370 13252
rect 13078 13240 13084 13252
rect 9364 13212 13084 13240
rect 9364 13200 9370 13212
rect 13078 13200 13084 13212
rect 13136 13200 13142 13252
rect 8849 13175 8907 13181
rect 8849 13141 8861 13175
rect 8895 13172 8907 13175
rect 8938 13172 8944 13184
rect 8895 13144 8944 13172
rect 8895 13141 8907 13144
rect 8849 13135 8907 13141
rect 8938 13132 8944 13144
rect 8996 13132 9002 13184
rect 11885 13175 11943 13181
rect 11885 13141 11897 13175
rect 11931 13172 11943 13175
rect 12250 13172 12256 13184
rect 11931 13144 12256 13172
rect 11931 13141 11943 13144
rect 11885 13135 11943 13141
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 13170 13172 13176 13184
rect 12492 13144 13176 13172
rect 12492 13132 12498 13144
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 13872 13144 13917 13172
rect 13872 13132 13878 13144
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 3605 12971 3663 12977
rect 3605 12937 3617 12971
rect 3651 12968 3663 12971
rect 4338 12968 4344 12980
rect 3651 12940 4344 12968
rect 3651 12937 3663 12940
rect 3605 12931 3663 12937
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 4982 12968 4988 12980
rect 4943 12940 4988 12968
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 6270 12968 6276 12980
rect 5951 12940 6276 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 8386 12968 8392 12980
rect 6687 12940 8392 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 8754 12928 8760 12980
rect 8812 12968 8818 12980
rect 8849 12971 8907 12977
rect 8849 12968 8861 12971
rect 8812 12940 8861 12968
rect 8812 12928 8818 12940
rect 8849 12937 8861 12940
rect 8895 12937 8907 12971
rect 8849 12931 8907 12937
rect 10134 12928 10140 12980
rect 10192 12968 10198 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10192 12940 10425 12968
rect 10192 12928 10198 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 4062 12860 4068 12912
rect 4120 12900 4126 12912
rect 4120 12872 7236 12900
rect 4120 12860 4126 12872
rect 1210 12792 1216 12844
rect 1268 12832 1274 12844
rect 1857 12835 1915 12841
rect 1857 12832 1869 12835
rect 1268 12804 1869 12832
rect 1268 12792 1274 12804
rect 1479 12773 1507 12804
rect 1857 12801 1869 12804
rect 1903 12801 1915 12835
rect 1857 12795 1915 12801
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12832 5595 12835
rect 6914 12832 6920 12844
rect 5583 12804 6920 12832
rect 5583 12801 5595 12804
rect 5537 12795 5595 12801
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7208 12841 7236 12872
rect 8202 12860 8208 12912
rect 8260 12900 8266 12912
rect 8665 12903 8723 12909
rect 8665 12900 8677 12903
rect 8260 12872 8677 12900
rect 8260 12860 8266 12872
rect 8665 12869 8677 12872
rect 8711 12869 8723 12903
rect 8665 12863 8723 12869
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12832 7251 12835
rect 7558 12832 7564 12844
rect 7239 12804 7564 12832
rect 7239 12801 7251 12804
rect 7193 12795 7251 12801
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 8754 12832 8760 12844
rect 8667 12804 8760 12832
rect 8754 12792 8760 12804
rect 8812 12832 8818 12844
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 8812 12804 9413 12832
rect 8812 12792 8818 12804
rect 9401 12801 9413 12804
rect 9447 12801 9459 12835
rect 10428 12832 10456 12931
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11940 12940 11989 12968
rect 11940 12928 11946 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 11977 12931 12035 12937
rect 13541 12971 13599 12977
rect 13541 12937 13553 12971
rect 13587 12968 13599 12971
rect 13630 12968 13636 12980
rect 13587 12940 13636 12968
rect 13587 12937 13599 12940
rect 13541 12931 13599 12937
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 15286 12968 15292 12980
rect 13872 12940 13917 12968
rect 15247 12940 15292 12968
rect 13872 12928 13878 12940
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 10428 12804 10961 12832
rect 9401 12795 9459 12801
rect 1464 12767 1522 12773
rect 1464 12733 1476 12767
rect 1510 12733 1522 12767
rect 1464 12727 1522 12733
rect 3237 12767 3295 12773
rect 3237 12733 3249 12767
rect 3283 12764 3295 12767
rect 4065 12767 4123 12773
rect 4065 12764 4077 12767
rect 3283 12736 4077 12764
rect 3283 12733 3295 12736
rect 3237 12727 3295 12733
rect 4065 12733 4077 12736
rect 4111 12764 4123 12767
rect 4706 12764 4712 12776
rect 4111 12736 4712 12764
rect 4111 12733 4123 12736
rect 4065 12727 4123 12733
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 8536 12767 8594 12773
rect 8536 12764 8548 12767
rect 7852 12736 8548 12764
rect 3973 12699 4031 12705
rect 3973 12665 3985 12699
rect 4019 12696 4031 12699
rect 4427 12699 4485 12705
rect 4427 12696 4439 12699
rect 4019 12668 4439 12696
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 4427 12665 4439 12668
rect 4473 12696 4485 12699
rect 4614 12696 4620 12708
rect 4473 12668 4620 12696
rect 4473 12665 4485 12668
rect 4427 12659 4485 12665
rect 4614 12656 4620 12668
rect 4672 12656 4678 12708
rect 6270 12656 6276 12708
rect 6328 12696 6334 12708
rect 7009 12699 7067 12705
rect 6328 12668 6776 12696
rect 6328 12656 6334 12668
rect 1535 12631 1593 12637
rect 1535 12597 1547 12631
rect 1581 12628 1593 12631
rect 3050 12628 3056 12640
rect 1581 12600 3056 12628
rect 1581 12597 1593 12600
rect 1535 12591 1593 12597
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 6748 12628 6776 12668
rect 7009 12665 7021 12699
rect 7055 12665 7067 12699
rect 7009 12659 7067 12665
rect 7024 12628 7052 12659
rect 6748 12600 7052 12628
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 7852 12637 7880 12736
rect 8536 12733 8548 12736
rect 8582 12733 8594 12767
rect 8536 12727 8594 12733
rect 10597 12767 10655 12773
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 10686 12764 10692 12776
rect 10643 12736 10692 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 8389 12699 8447 12705
rect 8389 12665 8401 12699
rect 8435 12696 8447 12699
rect 8938 12696 8944 12708
rect 8435 12668 8944 12696
rect 8435 12665 8447 12668
rect 8389 12659 8447 12665
rect 8938 12656 8944 12668
rect 8996 12656 9002 12708
rect 10933 12705 10961 12804
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12768 12804 12817 12832
rect 12768 12792 12774 12804
rect 12805 12801 12817 12804
rect 12851 12801 12863 12835
rect 14090 12832 14096 12844
rect 14051 12804 14096 12832
rect 12805 12795 12863 12801
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14366 12832 14372 12844
rect 14327 12804 14372 12832
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 10137 12699 10195 12705
rect 10137 12665 10149 12699
rect 10183 12696 10195 12699
rect 10918 12699 10976 12705
rect 10183 12668 10824 12696
rect 10183 12665 10195 12668
rect 10137 12659 10195 12665
rect 7837 12631 7895 12637
rect 7837 12628 7849 12631
rect 7340 12600 7849 12628
rect 7340 12588 7346 12600
rect 7837 12597 7849 12600
rect 7883 12597 7895 12631
rect 8202 12628 8208 12640
rect 8163 12600 8208 12628
rect 7837 12591 7895 12597
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 10796 12628 10824 12668
rect 10918 12665 10930 12699
rect 10964 12696 10976 12699
rect 12158 12696 12164 12708
rect 10964 12668 12164 12696
rect 10964 12665 10976 12668
rect 10918 12659 10976 12665
rect 12158 12656 12164 12668
rect 12216 12656 12222 12708
rect 12250 12656 12256 12708
rect 12308 12696 12314 12708
rect 12529 12699 12587 12705
rect 12529 12696 12541 12699
rect 12308 12668 12541 12696
rect 12308 12656 12314 12668
rect 12529 12665 12541 12668
rect 12575 12665 12587 12699
rect 12529 12659 12587 12665
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 14185 12699 14243 12705
rect 12676 12668 12721 12696
rect 12676 12656 12682 12668
rect 14185 12665 14197 12699
rect 14231 12665 14243 12699
rect 14185 12659 14243 12665
rect 11054 12628 11060 12640
rect 10796 12600 11060 12628
rect 11054 12588 11060 12600
rect 11112 12628 11118 12640
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 11112 12600 11529 12628
rect 11112 12588 11118 12600
rect 11517 12597 11529 12600
rect 11563 12628 11575 12631
rect 12636 12628 12664 12656
rect 11563 12600 12664 12628
rect 11563 12597 11575 12600
rect 11517 12591 11575 12597
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 14200 12628 14228 12659
rect 15654 12628 15660 12640
rect 13872 12600 14228 12628
rect 15615 12600 15660 12628
rect 13872 12588 13878 12600
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 4212 12396 4261 12424
rect 4212 12384 4218 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4249 12387 4307 12393
rect 6270 12384 6276 12436
rect 6328 12424 6334 12436
rect 6365 12427 6423 12433
rect 6365 12424 6377 12427
rect 6328 12396 6377 12424
rect 6328 12384 6334 12396
rect 6365 12393 6377 12396
rect 6411 12393 6423 12427
rect 6365 12387 6423 12393
rect 11793 12427 11851 12433
rect 11793 12393 11805 12427
rect 11839 12424 11851 12427
rect 12066 12424 12072 12436
rect 11839 12396 12072 12424
rect 11839 12393 11851 12396
rect 11793 12387 11851 12393
rect 12066 12384 12072 12396
rect 12124 12424 12130 12436
rect 12253 12427 12311 12433
rect 12253 12424 12265 12427
rect 12124 12396 12265 12424
rect 12124 12384 12130 12396
rect 12253 12393 12265 12396
rect 12299 12393 12311 12427
rect 12618 12424 12624 12436
rect 12579 12396 12624 12424
rect 12253 12387 12311 12393
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14553 12427 14611 12433
rect 14553 12424 14565 12427
rect 14148 12396 14565 12424
rect 14148 12384 14154 12396
rect 14553 12393 14565 12396
rect 14599 12393 14611 12427
rect 18138 12424 18144 12436
rect 18051 12396 18144 12424
rect 14553 12387 14611 12393
rect 18138 12384 18144 12396
rect 18196 12424 18202 12436
rect 19978 12424 19984 12436
rect 18196 12396 19984 12424
rect 18196 12384 18202 12396
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 4614 12316 4620 12368
rect 4672 12356 4678 12368
rect 5534 12356 5540 12368
rect 4672 12328 5540 12356
rect 4672 12316 4678 12328
rect 5534 12316 5540 12328
rect 5592 12356 5598 12368
rect 5766 12359 5824 12365
rect 5766 12356 5778 12359
rect 5592 12328 5778 12356
rect 5592 12316 5598 12328
rect 5766 12325 5778 12328
rect 5812 12325 5824 12359
rect 5766 12319 5824 12325
rect 6730 12316 6736 12368
rect 6788 12356 6794 12368
rect 7377 12359 7435 12365
rect 7377 12356 7389 12359
rect 6788 12328 7389 12356
rect 6788 12316 6794 12328
rect 7377 12325 7389 12328
rect 7423 12356 7435 12359
rect 7742 12356 7748 12368
rect 7423 12328 7748 12356
rect 7423 12325 7435 12328
rect 7377 12319 7435 12325
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 10413 12359 10471 12365
rect 10413 12325 10425 12359
rect 10459 12356 10471 12359
rect 10686 12356 10692 12368
rect 10459 12328 10692 12356
rect 10459 12325 10471 12328
rect 10413 12319 10471 12325
rect 10686 12316 10692 12328
rect 10744 12356 10750 12368
rect 11057 12359 11115 12365
rect 11057 12356 11069 12359
rect 10744 12328 11069 12356
rect 10744 12316 10750 12328
rect 11057 12325 11069 12328
rect 11103 12325 11115 12359
rect 11057 12319 11115 12325
rect 13081 12359 13139 12365
rect 13081 12325 13093 12359
rect 13127 12356 13139 12359
rect 13630 12356 13636 12368
rect 13127 12328 13636 12356
rect 13127 12325 13139 12328
rect 13081 12319 13139 12325
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 9674 12288 9680 12300
rect 9635 12260 9680 12288
rect 9674 12248 9680 12260
rect 9732 12288 9738 12300
rect 9950 12288 9956 12300
rect 9732 12260 9956 12288
rect 9732 12248 9738 12260
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12288 10287 12291
rect 10870 12288 10876 12300
rect 10275 12260 10876 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 15378 12288 15384 12300
rect 15339 12260 15384 12288
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 5442 12220 5448 12232
rect 5403 12192 5448 12220
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 6512 12192 7297 12220
rect 6512 12180 6518 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7558 12220 7564 12232
rect 7519 12192 7564 12220
rect 7285 12183 7343 12189
rect 7558 12180 7564 12192
rect 7616 12180 7622 12232
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 12986 12220 12992 12232
rect 12947 12192 12992 12220
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 9784 12152 9812 12180
rect 12894 12152 12900 12164
rect 9784 12124 12900 12152
rect 12894 12112 12900 12124
rect 12952 12112 12958 12164
rect 13541 12155 13599 12161
rect 13541 12121 13553 12155
rect 13587 12152 13599 12155
rect 13722 12152 13728 12164
rect 13587 12124 13728 12152
rect 13587 12121 13599 12124
rect 13541 12115 13599 12121
rect 13722 12112 13728 12124
rect 13780 12152 13786 12164
rect 14366 12152 14372 12164
rect 13780 12124 14372 12152
rect 13780 12112 13786 12124
rect 14366 12112 14372 12124
rect 14424 12112 14430 12164
rect 6917 12087 6975 12093
rect 6917 12053 6929 12087
rect 6963 12084 6975 12087
rect 7190 12084 7196 12096
rect 6963 12056 7196 12084
rect 6963 12053 6975 12056
rect 6917 12047 6975 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8389 12087 8447 12093
rect 8389 12084 8401 12087
rect 8260 12056 8401 12084
rect 8260 12044 8266 12056
rect 8389 12053 8401 12056
rect 8435 12053 8447 12087
rect 8389 12047 8447 12053
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 8757 12087 8815 12093
rect 8757 12084 8769 12087
rect 8628 12056 8769 12084
rect 8628 12044 8634 12056
rect 8757 12053 8769 12056
rect 8803 12084 8815 12087
rect 9766 12084 9772 12096
rect 8803 12056 9772 12084
rect 8803 12053 8815 12056
rect 8757 12047 8815 12053
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 10686 12084 10692 12096
rect 10647 12056 10692 12084
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 14274 12084 14280 12096
rect 14235 12056 14280 12084
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 15746 12084 15752 12096
rect 15707 12056 15752 12084
rect 15746 12044 15752 12056
rect 15804 12044 15810 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 5592 11852 5641 11880
rect 5592 11840 5598 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 5629 11843 5687 11849
rect 6178 11840 6184 11892
rect 6236 11880 6242 11892
rect 7285 11883 7343 11889
rect 7285 11880 7297 11883
rect 6236 11852 7297 11880
rect 6236 11840 6242 11852
rect 7285 11849 7297 11852
rect 7331 11849 7343 11883
rect 7285 11843 7343 11849
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 8570 11889 8576 11892
rect 7837 11883 7895 11889
rect 7837 11880 7849 11883
rect 7800 11852 7849 11880
rect 7800 11840 7806 11852
rect 7837 11849 7849 11852
rect 7883 11849 7895 11883
rect 8527 11883 8576 11889
rect 8527 11880 8539 11883
rect 7837 11843 7895 11849
rect 7925 11852 8539 11880
rect 6990 11815 7048 11821
rect 6990 11781 7002 11815
rect 7036 11812 7048 11815
rect 7098 11812 7104 11824
rect 7036 11784 7104 11812
rect 7036 11781 7048 11784
rect 6990 11775 7048 11781
rect 7098 11772 7104 11784
rect 7156 11812 7162 11824
rect 7925 11812 7953 11852
rect 8527 11849 8539 11852
rect 8573 11849 8576 11883
rect 8527 11843 8576 11849
rect 8570 11840 8576 11843
rect 8628 11840 8634 11892
rect 9030 11880 9036 11892
rect 8991 11852 9036 11880
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9674 11880 9680 11892
rect 9635 11852 9680 11880
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 10118 11883 10176 11889
rect 10118 11880 10130 11883
rect 9824 11852 10130 11880
rect 9824 11840 9830 11852
rect 10118 11849 10130 11852
rect 10164 11880 10176 11883
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 10164 11852 10977 11880
rect 10164 11849 10176 11852
rect 10118 11843 10176 11849
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 10965 11843 11023 11849
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 13357 11883 13415 11889
rect 13357 11849 13369 11883
rect 13403 11880 13415 11883
rect 13630 11880 13636 11892
rect 13403 11852 13636 11880
rect 13403 11849 13415 11852
rect 13357 11843 13415 11849
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 15105 11883 15163 11889
rect 15105 11849 15117 11883
rect 15151 11880 15163 11883
rect 15378 11880 15384 11892
rect 15151 11852 15384 11880
rect 15151 11849 15163 11852
rect 15105 11843 15163 11849
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 15746 11880 15752 11892
rect 15707 11852 15752 11880
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 7156 11784 7953 11812
rect 7156 11772 7162 11784
rect 8202 11772 8208 11824
rect 8260 11812 8266 11824
rect 8665 11815 8723 11821
rect 8665 11812 8677 11815
rect 8260 11784 8677 11812
rect 8260 11772 8266 11784
rect 8665 11781 8677 11784
rect 8711 11781 8723 11815
rect 8665 11775 8723 11781
rect 9585 11815 9643 11821
rect 9585 11781 9597 11815
rect 9631 11812 9643 11815
rect 10229 11815 10287 11821
rect 10229 11812 10241 11815
rect 9631 11784 10241 11812
rect 9631 11781 9643 11784
rect 9585 11775 9643 11781
rect 10229 11781 10241 11784
rect 10275 11812 10287 11815
rect 10686 11812 10692 11824
rect 10275 11784 10692 11812
rect 10275 11781 10287 11784
rect 10229 11775 10287 11781
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 6362 11744 6368 11756
rect 4571 11716 6368 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 4908 11685 4936 11716
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11744 6699 11747
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 6687 11716 7205 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 7193 11713 7205 11716
rect 7239 11744 7251 11747
rect 7834 11744 7840 11756
rect 7239 11716 7840 11744
rect 7239 11713 7251 11716
rect 7193 11707 7251 11713
rect 7834 11704 7840 11716
rect 7892 11744 7898 11756
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 7892 11716 8309 11744
rect 7892 11704 7898 11716
rect 8297 11713 8309 11716
rect 8343 11744 8355 11747
rect 8757 11747 8815 11753
rect 8757 11744 8769 11747
rect 8343 11716 8769 11744
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 8757 11713 8769 11716
rect 8803 11744 8815 11747
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 8803 11716 10333 11744
rect 8803 11713 8815 11716
rect 8757 11707 8815 11713
rect 10198 11688 10226 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 16022 11704 16028 11756
rect 16080 11744 16086 11756
rect 16301 11747 16359 11753
rect 16301 11744 16313 11747
rect 16080 11716 16313 11744
rect 16080 11704 16086 11716
rect 16301 11713 16313 11716
rect 16347 11713 16359 11747
rect 18138 11744 18144 11756
rect 18099 11716 18144 11744
rect 16301 11707 16359 11713
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 18414 11744 18420 11756
rect 18375 11716 18420 11744
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 1740 11679 1798 11685
rect 1740 11645 1752 11679
rect 1786 11676 1798 11679
rect 4893 11679 4951 11685
rect 1786 11648 2268 11676
rect 1786 11645 1798 11648
rect 1740 11639 1798 11645
rect 2240 11552 2268 11648
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 5169 11679 5227 11685
rect 5169 11645 5181 11679
rect 5215 11676 5227 11679
rect 5534 11676 5540 11688
rect 5215 11648 5540 11676
rect 5215 11645 5227 11648
rect 5169 11639 5227 11645
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 6273 11679 6331 11685
rect 6273 11645 6285 11679
rect 6319 11676 6331 11679
rect 7055 11679 7113 11685
rect 7055 11676 7067 11679
rect 6319 11648 7067 11676
rect 6319 11645 6331 11648
rect 6273 11639 6331 11645
rect 7055 11645 7067 11648
rect 7101 11676 7113 11679
rect 8570 11676 8576 11688
rect 7101 11648 8576 11676
rect 7101 11645 7113 11648
rect 7055 11639 7113 11645
rect 8570 11636 8576 11648
rect 8628 11676 8634 11688
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 8628 11648 9597 11676
rect 8628 11636 8634 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 10134 11636 10140 11688
rect 10192 11648 10226 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 11808 11648 12449 11676
rect 10192 11636 10198 11648
rect 6825 11611 6883 11617
rect 6825 11577 6837 11611
rect 6871 11608 6883 11611
rect 7190 11608 7196 11620
rect 6871 11580 7196 11608
rect 6871 11577 6883 11580
rect 6825 11571 6883 11577
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 8389 11611 8447 11617
rect 8389 11577 8401 11611
rect 8435 11608 8447 11611
rect 8938 11608 8944 11620
rect 8435 11580 8944 11608
rect 8435 11577 8447 11580
rect 8389 11571 8447 11577
rect 8938 11568 8944 11580
rect 8996 11608 9002 11620
rect 9953 11611 10011 11617
rect 9953 11608 9965 11611
rect 8996 11580 9965 11608
rect 8996 11568 9002 11580
rect 9953 11577 9965 11580
rect 9999 11577 10011 11611
rect 9953 11571 10011 11577
rect 10689 11611 10747 11617
rect 10689 11577 10701 11611
rect 10735 11608 10747 11611
rect 10870 11608 10876 11620
rect 10735 11580 10876 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 10870 11568 10876 11580
rect 10928 11608 10934 11620
rect 11333 11611 11391 11617
rect 11333 11608 11345 11611
rect 10928 11580 11345 11608
rect 10928 11568 10934 11580
rect 11333 11577 11345 11580
rect 11379 11577 11391 11611
rect 11333 11571 11391 11577
rect 1394 11500 1400 11552
rect 1452 11540 1458 11552
rect 1811 11543 1869 11549
rect 1811 11540 1823 11543
rect 1452 11512 1823 11540
rect 1452 11500 1458 11512
rect 1811 11509 1823 11512
rect 1857 11509 1869 11543
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 1811 11503 1869 11509
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 4706 11540 4712 11552
rect 4667 11512 4712 11540
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 11514 11500 11520 11552
rect 11572 11540 11578 11552
rect 11808 11549 11836 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 14274 11676 14280 11688
rect 14231 11648 14280 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12758 11611 12816 11617
rect 12758 11608 12770 11611
rect 12216 11580 12770 11608
rect 12216 11568 12222 11580
rect 12758 11577 12770 11580
rect 12804 11608 12816 11611
rect 16025 11611 16083 11617
rect 16025 11608 16037 11611
rect 12804 11580 13814 11608
rect 12804 11577 12816 11580
rect 12758 11571 12816 11577
rect 13786 11552 13814 11580
rect 15396 11580 16037 11608
rect 15396 11552 15424 11580
rect 16025 11577 16037 11580
rect 16071 11577 16083 11611
rect 16025 11571 16083 11577
rect 16117 11611 16175 11617
rect 16117 11577 16129 11611
rect 16163 11577 16175 11611
rect 16117 11571 16175 11577
rect 18233 11611 18291 11617
rect 18233 11577 18245 11611
rect 18279 11577 18291 11611
rect 18233 11571 18291 11577
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11572 11512 11805 11540
rect 11572 11500 11578 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 13786 11512 13820 11552
rect 11793 11503 11851 11509
rect 13814 11500 13820 11512
rect 13872 11540 13878 11552
rect 14093 11543 14151 11549
rect 14093 11540 14105 11543
rect 13872 11512 14105 11540
rect 13872 11500 13878 11512
rect 14093 11509 14105 11512
rect 14139 11540 14151 11543
rect 14550 11540 14556 11552
rect 14139 11512 14556 11540
rect 14139 11509 14151 11512
rect 14093 11503 14151 11509
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 15378 11540 15384 11552
rect 15339 11512 15384 11540
rect 15378 11500 15384 11512
rect 15436 11500 15442 11552
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 16132 11540 16160 11571
rect 17770 11540 17776 11552
rect 15804 11512 16160 11540
rect 17731 11512 17776 11540
rect 15804 11500 15810 11512
rect 17770 11500 17776 11512
rect 17828 11540 17834 11552
rect 18248 11540 18276 11571
rect 17828 11512 18276 11540
rect 17828 11500 17834 11512
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 5353 11339 5411 11345
rect 5353 11305 5365 11339
rect 5399 11336 5411 11339
rect 5442 11336 5448 11348
rect 5399 11308 5448 11336
rect 5399 11305 5411 11308
rect 5353 11299 5411 11305
rect 5442 11296 5448 11308
rect 5500 11336 5506 11348
rect 6089 11339 6147 11345
rect 6089 11336 6101 11339
rect 5500 11308 6101 11336
rect 5500 11296 5506 11308
rect 6089 11305 6101 11308
rect 6135 11305 6147 11339
rect 6089 11299 6147 11305
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 6604 11308 7389 11336
rect 6604 11296 6610 11308
rect 7377 11305 7389 11308
rect 7423 11336 7435 11339
rect 8754 11336 8760 11348
rect 7423 11308 8760 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9953 11339 10011 11345
rect 9953 11336 9965 11339
rect 9364 11308 9965 11336
rect 9364 11296 9370 11308
rect 9953 11305 9965 11308
rect 9999 11305 10011 11339
rect 9953 11299 10011 11305
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10229 11339 10287 11345
rect 10229 11336 10241 11339
rect 10192 11308 10241 11336
rect 10192 11296 10198 11308
rect 10229 11305 10241 11308
rect 10275 11305 10287 11339
rect 10229 11299 10287 11305
rect 12529 11339 12587 11345
rect 12529 11305 12541 11339
rect 12575 11305 12587 11339
rect 12986 11336 12992 11348
rect 12947 11308 12992 11336
rect 12529 11299 12587 11305
rect 7190 11228 7196 11280
rect 7248 11268 7254 11280
rect 7469 11271 7527 11277
rect 7469 11268 7481 11271
rect 7248 11240 7481 11268
rect 7248 11228 7254 11240
rect 7469 11237 7481 11240
rect 7515 11268 7527 11271
rect 8294 11268 8300 11280
rect 7515 11240 8300 11268
rect 7515 11237 7527 11240
rect 7469 11231 7527 11237
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 9674 11228 9680 11280
rect 9732 11268 9738 11280
rect 10962 11268 10968 11280
rect 9732 11240 10968 11268
rect 9732 11228 9738 11240
rect 10962 11228 10968 11240
rect 11020 11268 11026 11280
rect 12544 11268 12572 11299
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 14185 11339 14243 11345
rect 14185 11305 14197 11339
rect 14231 11336 14243 11339
rect 15378 11336 15384 11348
rect 14231 11308 15384 11336
rect 14231 11305 14243 11308
rect 14185 11299 14243 11305
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 17770 11336 17776 11348
rect 15528 11308 15573 11336
rect 17731 11308 17776 11336
rect 15528 11296 15534 11308
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 11020 11240 12572 11268
rect 11020 11228 11026 11240
rect 14550 11228 14556 11280
rect 14608 11268 14614 11280
rect 16111 11271 16169 11277
rect 16111 11268 16123 11271
rect 14608 11240 16123 11268
rect 14608 11228 14614 11240
rect 16111 11237 16123 11240
rect 16157 11268 16169 11271
rect 16298 11268 16304 11280
rect 16157 11240 16304 11268
rect 16157 11237 16169 11240
rect 16111 11231 16169 11237
rect 16298 11228 16304 11240
rect 16356 11228 16362 11280
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 5166 11200 5172 11212
rect 5127 11172 5172 11200
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 5592 11172 5641 11200
rect 5592 11160 5598 11172
rect 5629 11169 5641 11172
rect 5675 11200 5687 11203
rect 5675 11172 6224 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 5552 11132 5580 11160
rect 4755 11104 5580 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 1578 11064 1584 11076
rect 1539 11036 1584 11064
rect 1578 11024 1584 11036
rect 1636 11024 1642 11076
rect 6196 11064 6224 11172
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 9769 11203 9827 11209
rect 9769 11200 9781 11203
rect 9640 11172 9781 11200
rect 9640 11160 9646 11172
rect 9769 11169 9781 11172
rect 9815 11200 9827 11203
rect 10781 11203 10839 11209
rect 10781 11200 10793 11203
rect 9815 11172 10793 11200
rect 9815 11169 9827 11172
rect 9769 11163 9827 11169
rect 10781 11169 10793 11172
rect 10827 11169 10839 11203
rect 10781 11163 10839 11169
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11200 11483 11203
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 11471 11172 12357 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 12345 11169 12357 11172
rect 12391 11200 12403 11203
rect 12710 11200 12716 11212
rect 12391 11172 12716 11200
rect 12391 11169 12403 11172
rect 12345 11163 12403 11169
rect 7834 11132 7840 11144
rect 7795 11104 7840 11132
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 10796 11132 10824 11163
rect 12710 11160 12716 11172
rect 12768 11160 12774 11212
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11200 16727 11203
rect 17586 11200 17592 11212
rect 16715 11172 17592 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 24581 11203 24639 11209
rect 24581 11169 24593 11203
rect 24627 11200 24639 11203
rect 24670 11200 24676 11212
rect 24627 11172 24676 11200
rect 24627 11169 24639 11172
rect 24581 11163 24639 11169
rect 24670 11160 24676 11172
rect 24728 11160 24734 11212
rect 11238 11132 11244 11144
rect 10796 11104 11244 11132
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 15746 11132 15752 11144
rect 15707 11104 15752 11132
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 7929 11067 7987 11073
rect 7929 11064 7941 11067
rect 6196 11036 7941 11064
rect 7929 11033 7941 11036
rect 7975 11033 7987 11067
rect 8938 11064 8944 11076
rect 8851 11036 8944 11064
rect 7929 11027 7987 11033
rect 8938 11024 8944 11036
rect 8996 11064 9002 11076
rect 9766 11064 9772 11076
rect 8996 11036 9772 11064
rect 8996 11024 9002 11036
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 10134 11024 10140 11076
rect 10192 11064 10198 11076
rect 11422 11064 11428 11076
rect 10192 11036 11428 11064
rect 10192 11024 10198 11036
rect 11422 11024 11428 11036
rect 11480 11024 11486 11076
rect 11882 11024 11888 11076
rect 11940 11064 11946 11076
rect 13357 11067 13415 11073
rect 13357 11064 13369 11067
rect 11940 11036 13369 11064
rect 11940 11024 11946 11036
rect 13357 11033 13369 11036
rect 13403 11064 13415 11067
rect 14090 11064 14096 11076
rect 13403 11036 14096 11064
rect 13403 11033 13415 11036
rect 13357 11027 13415 11033
rect 14090 11024 14096 11036
rect 14148 11024 14154 11076
rect 6454 10996 6460 11008
rect 6415 10968 6460 10996
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 6917 10999 6975 11005
rect 6917 10965 6929 10999
rect 6963 10996 6975 10999
rect 7282 10996 7288 11008
rect 6963 10968 7288 10996
rect 6963 10965 6975 10968
rect 6917 10959 6975 10965
rect 7282 10956 7288 10968
rect 7340 10996 7346 11008
rect 7607 10999 7665 11005
rect 7607 10996 7619 10999
rect 7340 10968 7619 10996
rect 7340 10956 7346 10968
rect 7607 10965 7619 10968
rect 7653 10965 7665 10999
rect 7607 10959 7665 10965
rect 7745 10999 7803 11005
rect 7745 10965 7757 10999
rect 7791 10996 7803 10999
rect 8202 10996 8208 11008
rect 7791 10968 8208 10996
rect 7791 10965 7803 10968
rect 7745 10959 7803 10965
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 8478 10996 8484 11008
rect 8439 10968 8484 10996
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 8570 10956 8576 11008
rect 8628 10996 8634 11008
rect 9217 10999 9275 11005
rect 9217 10996 9229 10999
rect 8628 10968 9229 10996
rect 8628 10956 8634 10968
rect 9217 10965 9229 10968
rect 9263 10965 9275 10999
rect 9784 10996 9812 11024
rect 10597 10999 10655 11005
rect 10597 10996 10609 10999
rect 9784 10968 10609 10996
rect 9217 10959 9275 10965
rect 10597 10965 10609 10968
rect 10643 10965 10655 10999
rect 13630 10996 13636 11008
rect 13591 10968 13636 10996
rect 10597 10959 10655 10965
rect 13630 10956 13636 10968
rect 13688 10956 13694 11008
rect 23934 10956 23940 11008
rect 23992 10996 23998 11008
rect 24719 10999 24777 11005
rect 24719 10996 24731 10999
rect 23992 10968 24731 10996
rect 23992 10956 23998 10968
rect 24719 10965 24731 10968
rect 24765 10965 24777 10999
rect 24719 10959 24777 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1394 10752 1400 10804
rect 1452 10792 1458 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1452 10764 1593 10792
rect 1452 10752 1458 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 5166 10792 5172 10804
rect 5127 10764 5172 10792
rect 1581 10755 1639 10761
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5534 10792 5540 10804
rect 5495 10764 5540 10792
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 7834 10792 7840 10804
rect 7795 10764 7840 10792
rect 7834 10752 7840 10764
rect 7892 10752 7898 10804
rect 8570 10792 8576 10804
rect 8531 10764 8576 10792
rect 8570 10752 8576 10764
rect 8628 10752 8634 10804
rect 9582 10752 9588 10804
rect 9640 10792 9646 10804
rect 9769 10795 9827 10801
rect 9769 10792 9781 10795
rect 9640 10764 9781 10792
rect 9640 10752 9646 10764
rect 9769 10761 9781 10764
rect 9815 10761 9827 10795
rect 11882 10792 11888 10804
rect 11843 10764 11888 10792
rect 9769 10755 9827 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 14369 10795 14427 10801
rect 14369 10761 14381 10795
rect 14415 10792 14427 10795
rect 15197 10795 15255 10801
rect 15197 10792 15209 10795
rect 14415 10764 15209 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 15197 10761 15209 10764
rect 15243 10792 15255 10795
rect 15746 10792 15752 10804
rect 15243 10764 15752 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 17586 10792 17592 10804
rect 17547 10764 17592 10792
rect 17586 10752 17592 10764
rect 17644 10752 17650 10804
rect 24670 10792 24676 10804
rect 24631 10764 24676 10792
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 6641 10727 6699 10733
rect 6641 10693 6653 10727
rect 6687 10724 6699 10727
rect 7190 10724 7196 10736
rect 6687 10696 7196 10724
rect 6687 10693 6699 10696
rect 6641 10687 6699 10693
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 8754 10656 8760 10668
rect 8711 10628 8760 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10656 9091 10659
rect 11790 10656 11796 10668
rect 9079 10628 11796 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10656 15439 10659
rect 16761 10659 16819 10665
rect 16761 10656 16773 10659
rect 15427 10628 16773 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 16761 10625 16773 10628
rect 16807 10656 16819 10659
rect 18414 10656 18420 10668
rect 16807 10628 18420 10656
rect 16807 10625 16819 10628
rect 16761 10619 16819 10625
rect 18414 10616 18420 10628
rect 18472 10616 18478 10668
rect 8478 10597 8484 10600
rect 7285 10591 7343 10597
rect 7285 10588 7297 10591
rect 7116 10560 7297 10588
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7116 10461 7144 10560
rect 7285 10557 7297 10560
rect 7331 10588 7343 10591
rect 8444 10591 8484 10597
rect 8444 10588 8456 10591
rect 7331 10560 8456 10588
rect 7331 10557 7343 10560
rect 7285 10551 7343 10557
rect 8444 10557 8456 10560
rect 8444 10551 8484 10557
rect 8478 10548 8484 10551
rect 8536 10548 8542 10600
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10557 10471 10591
rect 10413 10551 10471 10557
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10588 11115 10591
rect 11146 10588 11152 10600
rect 11103 10560 11152 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 8294 10520 8300 10532
rect 8207 10492 8300 10520
rect 8294 10480 8300 10492
rect 8352 10480 8358 10532
rect 7101 10455 7159 10461
rect 7101 10452 7113 10455
rect 6972 10424 7113 10452
rect 6972 10412 6978 10424
rect 7101 10421 7113 10424
rect 7147 10421 7159 10455
rect 7101 10415 7159 10421
rect 7282 10412 7288 10464
rect 7340 10452 7346 10464
rect 7469 10455 7527 10461
rect 7469 10452 7481 10455
rect 7340 10424 7481 10452
rect 7340 10412 7346 10424
rect 7469 10421 7481 10424
rect 7515 10421 7527 10455
rect 8202 10452 8208 10464
rect 8163 10424 8208 10452
rect 7469 10415 7527 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8312 10452 8340 10480
rect 9398 10452 9404 10464
rect 8312 10424 9404 10452
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 9824 10424 10241 10452
rect 9824 10412 9830 10424
rect 10229 10421 10241 10424
rect 10275 10452 10287 10455
rect 10428 10452 10456 10551
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10588 11299 10591
rect 11422 10588 11428 10600
rect 11287 10560 11428 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 11422 10548 11428 10560
rect 11480 10588 11486 10600
rect 11882 10588 11888 10600
rect 11480 10560 11888 10588
rect 11480 10548 11486 10560
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 13173 10591 13231 10597
rect 13173 10557 13185 10591
rect 13219 10588 13231 10591
rect 13446 10588 13452 10600
rect 13219 10560 13452 10588
rect 13219 10557 13231 10560
rect 13173 10551 13231 10557
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 13725 10591 13783 10597
rect 13725 10557 13737 10591
rect 13771 10557 13783 10591
rect 14090 10588 14096 10600
rect 14051 10560 14096 10588
rect 13725 10551 13783 10557
rect 11164 10520 11192 10548
rect 12161 10523 12219 10529
rect 12161 10520 12173 10523
rect 11164 10492 12173 10520
rect 12161 10489 12173 10492
rect 12207 10520 12219 10523
rect 13630 10520 13636 10532
rect 12207 10492 13636 10520
rect 12207 10489 12219 10492
rect 12161 10483 12219 10489
rect 13630 10480 13636 10492
rect 13688 10520 13694 10532
rect 13740 10520 13768 10551
rect 14090 10548 14096 10560
rect 14148 10548 14154 10600
rect 16022 10548 16028 10600
rect 16080 10588 16086 10600
rect 16080 10560 16125 10588
rect 16080 10548 16086 10560
rect 13688 10492 13768 10520
rect 13688 10480 13694 10492
rect 15470 10480 15476 10532
rect 15528 10520 15534 10532
rect 15528 10492 15573 10520
rect 15528 10480 15534 10492
rect 10275 10424 10456 10452
rect 10689 10455 10747 10461
rect 10275 10421 10287 10424
rect 10229 10415 10287 10421
rect 10689 10421 10701 10455
rect 10735 10452 10747 10455
rect 10778 10452 10784 10464
rect 10735 10424 10784 10452
rect 10735 10421 10747 10424
rect 10689 10415 10747 10421
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 12710 10452 12716 10464
rect 12671 10424 12716 10452
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 14829 10455 14887 10461
rect 14829 10421 14841 10455
rect 14875 10452 14887 10455
rect 15488 10452 15516 10480
rect 16298 10452 16304 10464
rect 14875 10424 15516 10452
rect 16259 10424 16304 10452
rect 14875 10421 14887 10424
rect 14829 10415 14887 10421
rect 16298 10412 16304 10424
rect 16356 10412 16362 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 6822 10248 6828 10260
rect 6783 10220 6828 10248
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7653 10251 7711 10257
rect 7653 10217 7665 10251
rect 7699 10248 7711 10251
rect 8570 10248 8576 10260
rect 7699 10220 8576 10248
rect 7699 10217 7711 10220
rect 7653 10211 7711 10217
rect 8570 10208 8576 10220
rect 8628 10248 8634 10260
rect 9122 10248 9128 10260
rect 8628 10220 9128 10248
rect 8628 10208 8634 10220
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 12526 10248 12532 10260
rect 12487 10220 12532 10248
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 14274 10248 14280 10260
rect 14235 10220 14280 10248
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 23382 10208 23388 10260
rect 23440 10248 23446 10260
rect 23934 10248 23940 10260
rect 23440 10220 23940 10248
rect 23440 10208 23446 10220
rect 23934 10208 23940 10220
rect 23992 10208 23998 10260
rect 6181 10183 6239 10189
rect 6181 10149 6193 10183
rect 6227 10180 6239 10183
rect 7190 10180 7196 10192
rect 6227 10152 7196 10180
rect 6227 10149 6239 10152
rect 6181 10143 6239 10149
rect 7190 10140 7196 10152
rect 7248 10140 7254 10192
rect 8481 10183 8539 10189
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 8846 10180 8852 10192
rect 8527 10152 8852 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 8846 10140 8852 10152
rect 8904 10140 8910 10192
rect 9398 10140 9404 10192
rect 9456 10180 9462 10192
rect 17313 10183 17371 10189
rect 9456 10152 11376 10180
rect 9456 10140 9462 10152
rect 6328 10115 6386 10121
rect 6328 10081 6340 10115
rect 6374 10112 6386 10115
rect 6638 10112 6644 10124
rect 6374 10084 6644 10112
rect 6374 10081 6386 10084
rect 6328 10075 6386 10081
rect 6638 10072 6644 10084
rect 6696 10112 6702 10124
rect 7282 10112 7288 10124
rect 6696 10084 7288 10112
rect 6696 10072 6702 10084
rect 7282 10072 7288 10084
rect 7340 10112 7346 10124
rect 7469 10115 7527 10121
rect 7469 10112 7481 10115
rect 7340 10084 7481 10112
rect 7340 10072 7346 10084
rect 7469 10081 7481 10084
rect 7515 10081 7527 10115
rect 7469 10075 7527 10081
rect 7745 10115 7803 10121
rect 7745 10081 7757 10115
rect 7791 10081 7803 10115
rect 8202 10112 8208 10124
rect 7745 10075 7803 10081
rect 7944 10084 8208 10112
rect 6546 10044 6552 10056
rect 6507 10016 6552 10044
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 7098 10004 7104 10056
rect 7156 10044 7162 10056
rect 7760 10044 7788 10075
rect 7944 10044 7972 10084
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 9674 10112 9680 10124
rect 9635 10084 9680 10112
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10112 10287 10115
rect 10870 10112 10876 10124
rect 10275 10084 10876 10112
rect 10275 10081 10287 10084
rect 10229 10075 10287 10081
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 11238 10112 11244 10124
rect 11199 10084 11244 10112
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11348 10112 11376 10152
rect 17313 10149 17325 10183
rect 17359 10180 17371 10183
rect 17586 10180 17592 10192
rect 17359 10152 17592 10180
rect 17359 10149 17371 10152
rect 17313 10143 17371 10149
rect 17586 10140 17592 10152
rect 17644 10140 17650 10192
rect 17865 10183 17923 10189
rect 17865 10149 17877 10183
rect 17911 10180 17923 10183
rect 18414 10180 18420 10192
rect 17911 10152 18420 10180
rect 17911 10149 17923 10152
rect 17865 10143 17923 10149
rect 18414 10140 18420 10152
rect 18472 10140 18478 10192
rect 13446 10112 13452 10124
rect 11348 10084 13452 10112
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 13630 10112 13636 10124
rect 13591 10084 13636 10112
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 13998 10112 14004 10124
rect 13786 10084 14004 10112
rect 8110 10044 8116 10056
rect 7156 10016 7788 10044
rect 7852 10016 7972 10044
rect 8071 10016 8116 10044
rect 7156 10004 7162 10016
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 6457 9979 6515 9985
rect 6457 9976 6469 9979
rect 6328 9948 6469 9976
rect 6328 9936 6334 9948
rect 6457 9945 6469 9948
rect 6503 9976 6515 9979
rect 7852 9976 7880 10016
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9916 10016 10149 10044
rect 9916 10004 9922 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 11606 10044 11612 10056
rect 10137 10007 10195 10013
rect 11440 10016 11612 10044
rect 11440 9985 11468 10016
rect 11606 10004 11612 10016
rect 11664 10044 11670 10056
rect 13786 10044 13814 10084
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 14826 10072 14832 10124
rect 14884 10112 14890 10124
rect 15381 10115 15439 10121
rect 15381 10112 15393 10115
rect 14884 10084 15393 10112
rect 14884 10072 14890 10084
rect 15381 10081 15393 10084
rect 15427 10112 15439 10115
rect 15654 10112 15660 10124
rect 15427 10084 15660 10112
rect 15427 10081 15439 10084
rect 15381 10075 15439 10081
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 15838 10112 15844 10124
rect 15799 10084 15844 10112
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 16114 10044 16120 10056
rect 11664 10016 13814 10044
rect 16075 10016 16120 10044
rect 11664 10004 11670 10016
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 16960 10016 17233 10044
rect 6503 9948 7880 9976
rect 7910 9979 7968 9985
rect 6503 9945 6515 9948
rect 6457 9939 6515 9945
rect 7910 9945 7922 9979
rect 7956 9976 7968 9979
rect 11425 9979 11483 9985
rect 7956 9948 8156 9976
rect 7956 9945 7968 9948
rect 7910 9939 7968 9945
rect 8128 9920 8156 9948
rect 11425 9945 11437 9979
rect 11471 9945 11483 9979
rect 11425 9939 11483 9945
rect 16960 9920 16988 10016
rect 17221 10013 17233 10016
rect 17267 10013 17279 10047
rect 17221 10007 17279 10013
rect 7653 9911 7711 9917
rect 7653 9877 7665 9911
rect 7699 9908 7711 9911
rect 8021 9911 8079 9917
rect 8021 9908 8033 9911
rect 7699 9880 8033 9908
rect 7699 9877 7711 9880
rect 7653 9871 7711 9877
rect 8021 9877 8033 9880
rect 8067 9877 8079 9911
rect 8021 9871 8079 9877
rect 8110 9868 8116 9920
rect 8168 9868 8174 9920
rect 8754 9908 8760 9920
rect 8715 9880 8760 9908
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 10873 9911 10931 9917
rect 10873 9877 10885 9911
rect 10919 9908 10931 9911
rect 12710 9908 12716 9920
rect 10919 9880 12716 9908
rect 10919 9877 10931 9880
rect 10873 9871 10931 9877
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 16942 9908 16948 9920
rect 16903 9880 16948 9908
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 6178 9664 6184 9716
rect 6236 9704 6242 9716
rect 7469 9707 7527 9713
rect 7469 9704 7481 9707
rect 6236 9676 7481 9704
rect 6236 9664 6242 9676
rect 7469 9673 7481 9676
rect 7515 9704 7527 9707
rect 7834 9704 7840 9716
rect 7515 9676 7840 9704
rect 7515 9673 7527 9676
rect 7469 9667 7527 9673
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 8386 9704 8392 9716
rect 8347 9676 8392 9704
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 8478 9664 8484 9716
rect 8536 9704 8542 9716
rect 9309 9707 9367 9713
rect 9309 9704 9321 9707
rect 8536 9676 9321 9704
rect 8536 9664 8542 9676
rect 9309 9673 9321 9676
rect 9355 9704 9367 9707
rect 9631 9707 9689 9713
rect 9631 9704 9643 9707
rect 9355 9676 9643 9704
rect 9355 9673 9367 9676
rect 9309 9667 9367 9673
rect 9631 9673 9643 9676
rect 9677 9673 9689 9707
rect 10870 9704 10876 9716
rect 10831 9676 10876 9704
rect 9631 9667 9689 9673
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11296 9676 11805 9704
rect 11296 9664 11302 9676
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 13446 9704 13452 9716
rect 13407 9676 13452 9704
rect 11793 9667 11851 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 13909 9707 13967 9713
rect 13909 9673 13921 9707
rect 13955 9704 13967 9707
rect 13998 9704 14004 9716
rect 13955 9676 14004 9704
rect 13955 9673 13967 9676
rect 13909 9667 13967 9673
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 14458 9704 14464 9716
rect 14419 9676 14464 9704
rect 14458 9664 14464 9676
rect 14516 9664 14522 9716
rect 15654 9704 15660 9716
rect 15615 9676 15660 9704
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 17497 9707 17555 9713
rect 17497 9673 17509 9707
rect 17543 9704 17555 9707
rect 17586 9704 17592 9716
rect 17543 9676 17592 9704
rect 17543 9673 17555 9676
rect 17497 9667 17555 9673
rect 17586 9664 17592 9676
rect 17644 9664 17650 9716
rect 6270 9636 6276 9648
rect 6231 9608 6276 9636
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 6638 9636 6644 9648
rect 6599 9608 6644 9636
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 7101 9639 7159 9645
rect 7101 9605 7113 9639
rect 7147 9636 7159 9639
rect 7190 9636 7196 9648
rect 7147 9608 7196 9636
rect 7147 9605 7159 9608
rect 7101 9599 7159 9605
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 7116 9568 7144 9599
rect 7190 9596 7196 9608
rect 7248 9596 7254 9648
rect 5951 9540 7144 9568
rect 7852 9568 7880 9664
rect 8110 9645 8116 9648
rect 8094 9639 8116 9645
rect 8094 9605 8106 9639
rect 8094 9599 8116 9605
rect 8110 9596 8116 9599
rect 8168 9596 8174 9648
rect 8202 9596 8208 9648
rect 8260 9636 8266 9648
rect 8941 9639 8999 9645
rect 8941 9636 8953 9639
rect 8260 9608 8953 9636
rect 8260 9596 8266 9608
rect 8941 9605 8953 9608
rect 8987 9605 8999 9639
rect 8941 9599 8999 9605
rect 9122 9596 9128 9648
rect 9180 9636 9186 9648
rect 9769 9639 9827 9645
rect 9769 9636 9781 9639
rect 9180 9608 9781 9636
rect 9180 9596 9186 9608
rect 9769 9605 9781 9608
rect 9815 9636 9827 9639
rect 10042 9636 10048 9648
rect 9815 9608 10048 9636
rect 9815 9605 9827 9608
rect 9769 9599 9827 9605
rect 10042 9596 10048 9608
rect 10100 9596 10106 9648
rect 10137 9639 10195 9645
rect 10137 9605 10149 9639
rect 10183 9636 10195 9639
rect 15746 9636 15752 9648
rect 10183 9608 15752 9636
rect 10183 9605 10195 9608
rect 10137 9599 10195 9605
rect 15746 9596 15752 9608
rect 15804 9596 15810 9648
rect 8297 9571 8355 9577
rect 8297 9568 8309 9571
rect 7852 9540 8309 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 8297 9537 8309 9540
rect 8343 9537 8355 9571
rect 8297 9531 8355 9537
rect 8846 9528 8852 9580
rect 8904 9568 8910 9580
rect 9398 9568 9404 9580
rect 8904 9540 9404 9568
rect 8904 9528 8910 9540
rect 9398 9528 9404 9540
rect 9456 9568 9462 9580
rect 9861 9571 9919 9577
rect 9861 9568 9873 9571
rect 9456 9540 9873 9568
rect 9456 9528 9462 9540
rect 9861 9537 9873 9540
rect 9907 9537 9919 9571
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 9861 9531 9919 9537
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12802 9568 12808 9580
rect 12763 9540 12808 9568
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 16114 9528 16120 9580
rect 16172 9568 16178 9580
rect 16209 9571 16267 9577
rect 16209 9568 16221 9571
rect 16172 9540 16221 9568
rect 16172 9528 16178 9540
rect 16209 9537 16221 9540
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 23382 9528 23388 9580
rect 23440 9568 23446 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 23440 9540 23949 9568
rect 23440 9528 23446 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 6546 9500 6552 9512
rect 5583 9472 6552 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 6546 9460 6552 9472
rect 6604 9460 6610 9512
rect 6917 9503 6975 9509
rect 6917 9469 6929 9503
rect 6963 9500 6975 9503
rect 7098 9500 7104 9512
rect 6963 9472 7104 9500
rect 6963 9469 6975 9472
rect 6917 9463 6975 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9500 7987 9503
rect 8018 9500 8024 9512
rect 7975 9472 8024 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 8018 9460 8024 9472
rect 8076 9500 8082 9512
rect 8754 9500 8760 9512
rect 8076 9472 8760 9500
rect 8076 9460 8082 9472
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 9732 9472 10517 9500
rect 9732 9460 9738 9472
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 10505 9463 10563 9469
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 14645 9503 14703 9509
rect 14645 9500 14657 9503
rect 14516 9472 14657 9500
rect 14516 9460 14522 9472
rect 14645 9469 14657 9472
rect 14691 9469 14703 9503
rect 15102 9500 15108 9512
rect 15063 9472 15108 9500
rect 14645 9463 14703 9469
rect 15102 9460 15108 9472
rect 15160 9500 15166 9512
rect 15838 9500 15844 9512
rect 15160 9472 15844 9500
rect 15160 9460 15166 9472
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9500 17187 9503
rect 17865 9503 17923 9509
rect 17865 9500 17877 9503
rect 17175 9472 17877 9500
rect 17175 9469 17187 9472
rect 17129 9463 17187 9469
rect 17865 9469 17877 9472
rect 17911 9500 17923 9503
rect 18693 9503 18751 9509
rect 18693 9500 18705 9503
rect 17911 9472 18705 9500
rect 17911 9469 17923 9472
rect 17865 9463 17923 9469
rect 18693 9469 18705 9472
rect 18739 9500 18751 9503
rect 19058 9500 19064 9512
rect 18739 9472 19064 9500
rect 18739 9469 18751 9472
rect 18693 9463 18751 9469
rect 19058 9460 19064 9472
rect 19116 9460 19122 9512
rect 7190 9392 7196 9444
rect 7248 9432 7254 9444
rect 9493 9435 9551 9441
rect 9493 9432 9505 9435
rect 7248 9404 9505 9432
rect 7248 9392 7254 9404
rect 9493 9401 9505 9404
rect 9539 9432 9551 9435
rect 9766 9432 9772 9444
rect 9539 9404 9772 9432
rect 9539 9401 9551 9404
rect 9493 9395 9551 9401
rect 9766 9392 9772 9404
rect 9824 9392 9830 9444
rect 12253 9435 12311 9441
rect 12253 9401 12265 9435
rect 12299 9432 12311 9435
rect 12618 9432 12624 9444
rect 12299 9404 12624 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 12618 9392 12624 9404
rect 12676 9392 12682 9444
rect 15381 9435 15439 9441
rect 15381 9401 15393 9435
rect 15427 9432 15439 9435
rect 16206 9432 16212 9444
rect 15427 9404 16212 9432
rect 15427 9401 15439 9404
rect 15381 9395 15439 9401
rect 16206 9392 16212 9404
rect 16264 9392 16270 9444
rect 16298 9392 16304 9444
rect 16356 9432 16362 9444
rect 16571 9435 16629 9441
rect 16571 9432 16583 9435
rect 16356 9404 16583 9432
rect 16356 9392 16362 9404
rect 16571 9401 16583 9404
rect 16617 9432 16629 9435
rect 17402 9432 17408 9444
rect 16617 9404 17408 9432
rect 16617 9401 16629 9404
rect 16571 9395 16629 9401
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 18046 9432 18052 9444
rect 18007 9404 18052 9432
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 24029 9435 24087 9441
rect 24029 9401 24041 9435
rect 24075 9401 24087 9435
rect 24578 9432 24584 9444
rect 24539 9404 24584 9432
rect 24029 9395 24087 9401
rect 7837 9367 7895 9373
rect 7837 9333 7849 9367
rect 7883 9364 7895 9367
rect 7926 9364 7932 9376
rect 7883 9336 7932 9364
rect 7883 9333 7895 9336
rect 7837 9327 7895 9333
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 11330 9364 11336 9376
rect 11291 9336 11336 9364
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 16117 9367 16175 9373
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 16316 9364 16344 9392
rect 23382 9364 23388 9376
rect 16163 9336 16344 9364
rect 23343 9336 23388 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 23382 9324 23388 9336
rect 23440 9364 23446 9376
rect 24044 9364 24072 9395
rect 24578 9392 24584 9404
rect 24636 9392 24642 9444
rect 23440 9336 24072 9364
rect 23440 9324 23446 9336
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 6178 9160 6184 9172
rect 6139 9132 6184 9160
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 7190 9160 7196 9172
rect 7151 9132 7196 9160
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 9398 9160 9404 9172
rect 9359 9132 9404 9160
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 9861 9163 9919 9169
rect 9861 9160 9873 9163
rect 9824 9132 9873 9160
rect 9824 9120 9830 9132
rect 9861 9129 9873 9132
rect 9907 9129 9919 9163
rect 9861 9123 9919 9129
rect 8018 9092 8024 9104
rect 7024 9064 8024 9092
rect 7024 9036 7052 9064
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1670 9024 1676 9036
rect 1443 8996 1676 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 2501 9027 2559 9033
rect 2501 8993 2513 9027
rect 2547 9024 2559 9027
rect 2590 9024 2596 9036
rect 2547 8996 2596 9024
rect 2547 8993 2559 8996
rect 2501 8987 2559 8993
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 5997 9027 6055 9033
rect 5997 8993 6009 9027
rect 6043 9024 6055 9027
rect 6086 9024 6092 9036
rect 6043 8996 6092 9024
rect 6043 8993 6055 8996
rect 5997 8987 6055 8993
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 7006 9024 7012 9036
rect 6919 8996 7012 9024
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7837 9027 7895 9033
rect 7837 8993 7849 9027
rect 7883 9024 7895 9027
rect 8202 9024 8208 9036
rect 7883 8996 8208 9024
rect 7883 8993 7895 8996
rect 7837 8987 7895 8993
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8956 6975 8959
rect 7098 8956 7104 8968
rect 6963 8928 7104 8956
rect 6963 8925 6975 8928
rect 6917 8919 6975 8925
rect 7098 8916 7104 8928
rect 7156 8956 7162 8968
rect 7852 8956 7880 8987
rect 8202 8984 8208 8996
rect 8260 9024 8266 9036
rect 9033 9027 9091 9033
rect 9033 9024 9045 9027
rect 8260 8996 9045 9024
rect 8260 8984 8266 8996
rect 9033 8993 9045 8996
rect 9079 8993 9091 9027
rect 9876 9024 9904 9123
rect 10042 9120 10048 9172
rect 10100 9160 10106 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 10100 9132 10241 9160
rect 10100 9120 10106 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 12434 9160 12440 9172
rect 10229 9123 10287 9129
rect 11348 9132 12440 9160
rect 10594 9024 10600 9036
rect 9876 8996 10600 9024
rect 9033 8987 9091 8993
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 11146 9024 11152 9036
rect 11107 8996 11152 9024
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 7156 8928 7880 8956
rect 7156 8916 7162 8928
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 8076 8928 8401 8956
rect 8076 8916 8082 8928
rect 8389 8925 8401 8928
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 11348 8956 11376 9132
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 13814 9160 13820 9172
rect 13556 9132 13820 9160
rect 11882 9052 11888 9104
rect 11940 9092 11946 9104
rect 12850 9095 12908 9101
rect 12850 9092 12862 9095
rect 11940 9064 12862 9092
rect 11940 9052 11946 9064
rect 12850 9061 12862 9064
rect 12896 9092 12908 9095
rect 13556 9092 13584 9132
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 16114 9120 16120 9172
rect 16172 9160 16178 9172
rect 16301 9163 16359 9169
rect 16301 9160 16313 9163
rect 16172 9132 16313 9160
rect 16172 9120 16178 9132
rect 16301 9129 16313 9132
rect 16347 9129 16359 9163
rect 19518 9160 19524 9172
rect 16301 9123 16359 9129
rect 18708 9132 19524 9160
rect 12896 9064 13584 9092
rect 12896 9061 12908 9064
rect 12850 9055 12908 9061
rect 13630 9052 13636 9104
rect 13688 9092 13694 9104
rect 13725 9095 13783 9101
rect 13725 9092 13737 9095
rect 13688 9064 13737 9092
rect 13688 9052 13694 9064
rect 13725 9061 13737 9064
rect 13771 9061 13783 9095
rect 13725 9055 13783 9061
rect 17215 9095 17273 9101
rect 17215 9061 17227 9095
rect 17261 9092 17273 9095
rect 17402 9092 17408 9104
rect 17261 9064 17408 9092
rect 17261 9061 17273 9064
rect 17215 9055 17273 9061
rect 17402 9052 17408 9064
rect 17460 9052 17466 9104
rect 18708 9101 18736 9132
rect 19518 9120 19524 9132
rect 19576 9160 19582 9172
rect 24486 9160 24492 9172
rect 19576 9132 24492 9160
rect 19576 9120 19582 9132
rect 24486 9120 24492 9132
rect 24544 9120 24550 9172
rect 24854 9120 24860 9172
rect 24912 9160 24918 9172
rect 25547 9163 25605 9169
rect 25547 9160 25559 9163
rect 24912 9132 25559 9160
rect 24912 9120 24918 9132
rect 25547 9129 25559 9132
rect 25593 9129 25605 9163
rect 25547 9123 25605 9129
rect 18693 9095 18751 9101
rect 18693 9061 18705 9095
rect 18739 9061 18751 9095
rect 18693 9055 18751 9061
rect 18785 9095 18843 9101
rect 18785 9061 18797 9095
rect 18831 9092 18843 9095
rect 19058 9092 19064 9104
rect 18831 9064 19064 9092
rect 18831 9061 18843 9064
rect 18785 9055 18843 9061
rect 19058 9052 19064 9064
rect 19116 9052 19122 9104
rect 24026 9092 24032 9104
rect 23987 9064 24032 9092
rect 24026 9052 24032 9064
rect 24084 9052 24090 9104
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 9024 11483 9027
rect 11606 9024 11612 9036
rect 11471 8996 11612 9024
rect 11471 8993 11483 8996
rect 11425 8987 11483 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 14458 8984 14464 9036
rect 14516 9024 14522 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 14516 8996 15301 9024
rect 14516 8984 14522 8996
rect 15289 8993 15301 8996
rect 15335 9024 15347 9027
rect 15470 9024 15476 9036
rect 15335 8996 15476 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 15746 9024 15752 9036
rect 15707 8996 15752 9024
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 16758 9024 16764 9036
rect 16264 8996 16764 9024
rect 16264 8984 16270 8996
rect 16758 8984 16764 8996
rect 16816 9024 16822 9036
rect 16853 9027 16911 9033
rect 16853 9024 16865 9027
rect 16816 8996 16865 9024
rect 16816 8984 16822 8996
rect 16853 8993 16865 8996
rect 16899 8993 16911 9027
rect 16853 8987 16911 8993
rect 22741 9027 22799 9033
rect 22741 8993 22753 9027
rect 22787 9024 22799 9027
rect 22922 9024 22928 9036
rect 22787 8996 22928 9024
rect 22787 8993 22799 8996
rect 22741 8987 22799 8993
rect 22922 8984 22928 8996
rect 22980 8984 22986 9036
rect 24578 8984 24584 9036
rect 24636 9024 24642 9036
rect 25498 9033 25504 9036
rect 25476 9027 25504 9033
rect 25476 9024 25488 9027
rect 24636 8996 24681 9024
rect 25411 8996 25488 9024
rect 24636 8984 24642 8996
rect 25476 8993 25488 8996
rect 25556 9024 25562 9036
rect 27614 9024 27620 9036
rect 25556 8996 27620 9024
rect 25476 8987 25504 8993
rect 25498 8984 25504 8987
rect 25556 8984 25562 8996
rect 27614 8984 27620 8996
rect 27672 8984 27678 9036
rect 8803 8928 11376 8956
rect 11701 8959 11759 8965
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 11701 8925 11713 8959
rect 11747 8956 11759 8959
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 11747 8928 12541 8956
rect 11747 8925 11759 8928
rect 11701 8919 11759 8925
rect 12529 8925 12541 8928
rect 12575 8956 12587 8959
rect 13446 8956 13452 8968
rect 12575 8928 13452 8956
rect 12575 8925 12587 8928
rect 12529 8919 12587 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 16022 8956 16028 8968
rect 15983 8928 16028 8956
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 18782 8916 18788 8968
rect 18840 8956 18846 8968
rect 18969 8959 19027 8965
rect 18969 8956 18981 8959
rect 18840 8928 18981 8956
rect 18840 8916 18846 8928
rect 18969 8925 18981 8928
rect 19015 8925 19027 8959
rect 23934 8956 23940 8968
rect 23895 8928 23940 8956
rect 18969 8919 19027 8925
rect 23934 8916 23940 8928
rect 23992 8916 23998 8968
rect 1578 8888 1584 8900
rect 1539 8860 1584 8888
rect 1578 8848 1584 8860
rect 1636 8848 1642 8900
rect 7558 8848 7564 8900
rect 7616 8888 7622 8900
rect 8297 8891 8355 8897
rect 8297 8888 8309 8891
rect 7616 8860 8309 8888
rect 7616 8848 7622 8860
rect 8297 8857 8309 8860
rect 8343 8888 8355 8891
rect 9122 8888 9128 8900
rect 8343 8860 9128 8888
rect 8343 8857 8355 8860
rect 8297 8851 8355 8857
rect 9122 8848 9128 8860
rect 9180 8848 9186 8900
rect 15102 8848 15108 8900
rect 15160 8848 15166 8900
rect 17773 8891 17831 8897
rect 17773 8857 17785 8891
rect 17819 8888 17831 8891
rect 23382 8888 23388 8900
rect 17819 8860 23388 8888
rect 17819 8857 17831 8860
rect 17773 8851 17831 8857
rect 23382 8848 23388 8860
rect 23440 8848 23446 8900
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 2639 8823 2697 8829
rect 2639 8820 2651 8823
rect 1728 8792 2651 8820
rect 1728 8780 1734 8792
rect 2639 8789 2651 8792
rect 2685 8789 2697 8823
rect 6546 8820 6552 8832
rect 6507 8792 6552 8820
rect 2639 8783 2697 8789
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 8110 8780 8116 8832
rect 8168 8829 8174 8832
rect 8168 8823 8217 8829
rect 8168 8789 8171 8823
rect 8205 8789 8217 8823
rect 8168 8783 8217 8789
rect 8168 8780 8174 8783
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 13449 8823 13507 8829
rect 13449 8820 13461 8823
rect 12676 8792 13461 8820
rect 12676 8780 12682 8792
rect 13449 8789 13461 8792
rect 13495 8789 13507 8823
rect 14642 8820 14648 8832
rect 14603 8792 14648 8820
rect 13449 8783 13507 8789
rect 14642 8780 14648 8792
rect 14700 8820 14706 8832
rect 15013 8823 15071 8829
rect 15013 8820 15025 8823
rect 14700 8792 15025 8820
rect 14700 8780 14706 8792
rect 15013 8789 15025 8792
rect 15059 8820 15071 8823
rect 15120 8820 15148 8848
rect 18138 8820 18144 8832
rect 15059 8792 15148 8820
rect 18099 8792 18144 8820
rect 15059 8789 15071 8792
rect 15013 8783 15071 8789
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 22830 8780 22836 8832
rect 22888 8820 22894 8832
rect 22971 8823 23029 8829
rect 22971 8820 22983 8823
rect 22888 8792 22983 8820
rect 22888 8780 22894 8792
rect 22971 8789 22983 8792
rect 23017 8789 23029 8823
rect 22971 8783 23029 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 7006 8616 7012 8628
rect 6967 8588 7012 8616
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 7377 8619 7435 8625
rect 7377 8585 7389 8619
rect 7423 8616 7435 8619
rect 7558 8616 7564 8628
rect 7423 8588 7564 8616
rect 7423 8585 7435 8588
rect 7377 8579 7435 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 7834 8616 7840 8628
rect 7791 8588 7840 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 8352 8588 8493 8616
rect 8352 8576 8358 8588
rect 8481 8585 8493 8588
rect 8527 8616 8539 8619
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 8527 8588 9229 8616
rect 8527 8585 8539 8588
rect 8481 8579 8539 8585
rect 9217 8585 9229 8588
rect 9263 8616 9275 8619
rect 9953 8619 10011 8625
rect 9953 8616 9965 8619
rect 9263 8588 9965 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9953 8585 9965 8588
rect 9999 8585 10011 8619
rect 10594 8616 10600 8628
rect 10555 8588 10600 8616
rect 9953 8579 10011 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 14458 8616 14464 8628
rect 14415 8588 14464 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15654 8616 15660 8628
rect 15243 8588 15660 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 7852 8480 7880 8576
rect 11422 8548 11428 8560
rect 10888 8520 11428 8548
rect 8573 8483 8631 8489
rect 8573 8480 8585 8483
rect 7852 8452 8585 8480
rect 8573 8449 8585 8452
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9585 8483 9643 8489
rect 9585 8480 9597 8483
rect 9180 8452 9597 8480
rect 9180 8440 9186 8452
rect 9585 8449 9597 8452
rect 9631 8449 9643 8483
rect 9585 8443 9643 8449
rect 10888 8424 10916 8520
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 11514 8480 11520 8492
rect 11475 8452 11520 8480
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 7190 8412 7196 8424
rect 7151 8384 7196 8412
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 8110 8412 8116 8424
rect 7576 8384 8116 8412
rect 7576 8356 7604 8384
rect 8110 8372 8116 8384
rect 8168 8412 8174 8424
rect 8352 8415 8410 8421
rect 8352 8412 8364 8415
rect 8168 8384 8364 8412
rect 8168 8372 8174 8384
rect 8352 8381 8364 8384
rect 8398 8381 8410 8415
rect 8352 8375 8410 8381
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 9769 8415 9827 8421
rect 9769 8412 9781 8415
rect 8536 8384 9781 8412
rect 8536 8372 8542 8384
rect 9769 8381 9781 8384
rect 9815 8412 9827 8415
rect 10229 8415 10287 8421
rect 10229 8412 10241 8415
rect 9815 8384 10241 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 10229 8381 10241 8384
rect 10275 8381 10287 8415
rect 10870 8412 10876 8424
rect 10831 8384 10876 8412
rect 10229 8375 10287 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 11333 8415 11391 8421
rect 11333 8412 11345 8415
rect 11296 8384 11345 8412
rect 11296 8372 11302 8384
rect 11333 8381 11345 8384
rect 11379 8412 11391 8415
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 11379 8384 11805 8412
rect 11379 8381 11391 8384
rect 11333 8375 11391 8381
rect 11793 8381 11805 8384
rect 11839 8381 11851 8415
rect 12618 8412 12624 8424
rect 12579 8384 12624 8412
rect 11793 8375 11851 8381
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 15304 8421 15332 8588
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 16758 8616 16764 8628
rect 16719 8588 16764 8616
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 17402 8616 17408 8628
rect 17363 8588 17408 8616
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8616 17923 8619
rect 18046 8616 18052 8628
rect 17911 8588 18052 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 19058 8616 19064 8628
rect 19019 8588 19064 8616
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 19518 8616 19524 8628
rect 19479 8588 19524 8616
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 22922 8616 22928 8628
rect 22883 8588 22928 8616
rect 22922 8576 22928 8588
rect 22980 8576 22986 8628
rect 23382 8616 23388 8628
rect 23343 8588 23388 8616
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 25498 8616 25504 8628
rect 25459 8588 25504 8616
rect 25498 8576 25504 8588
rect 25556 8576 25562 8628
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8480 17003 8483
rect 18138 8480 18144 8492
rect 16991 8452 18144 8480
rect 16991 8449 17003 8452
rect 16945 8443 17003 8449
rect 18138 8440 18144 8452
rect 18196 8440 18202 8492
rect 18782 8480 18788 8492
rect 18743 8452 18788 8480
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 24026 8440 24032 8492
rect 24084 8480 24090 8492
rect 24397 8483 24455 8489
rect 24397 8480 24409 8483
rect 24084 8452 24409 8480
rect 24084 8440 24090 8452
rect 24397 8449 24409 8452
rect 24443 8480 24455 8483
rect 24673 8483 24731 8489
rect 24673 8480 24685 8483
rect 24443 8452 24685 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 24673 8449 24685 8452
rect 24719 8449 24731 8483
rect 24673 8443 24731 8449
rect 14185 8415 14243 8421
rect 14185 8412 14197 8415
rect 13786 8384 14197 8412
rect 6546 8304 6552 8356
rect 6604 8344 6610 8356
rect 6641 8347 6699 8353
rect 6641 8344 6653 8347
rect 6604 8316 6653 8344
rect 6604 8304 6610 8316
rect 6641 8313 6653 8316
rect 6687 8344 6699 8347
rect 7558 8344 7564 8356
rect 6687 8316 7564 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 8202 8344 8208 8356
rect 8163 8316 8208 8344
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8938 8344 8944 8356
rect 8899 8316 8944 8344
rect 8938 8304 8944 8316
rect 8996 8304 9002 8356
rect 11974 8304 11980 8356
rect 12032 8344 12038 8356
rect 12437 8347 12495 8353
rect 12437 8344 12449 8347
rect 12032 8316 12449 8344
rect 12032 8304 12038 8316
rect 12437 8313 12449 8316
rect 12483 8313 12495 8347
rect 12437 8307 12495 8313
rect 2590 8276 2596 8288
rect 2551 8248 2596 8276
rect 2590 8236 2596 8248
rect 2648 8236 2654 8288
rect 6086 8276 6092 8288
rect 6047 8248 6092 8276
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 8018 8276 8024 8288
rect 7979 8248 8024 8276
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 11882 8236 11888 8288
rect 11940 8276 11946 8288
rect 12161 8279 12219 8285
rect 12161 8276 12173 8279
rect 11940 8248 12173 8276
rect 11940 8236 11946 8248
rect 12161 8245 12173 8248
rect 12207 8245 12219 8279
rect 12161 8239 12219 8245
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 13630 8276 13636 8288
rect 12768 8248 13636 8276
rect 12768 8236 12774 8248
rect 13630 8236 13636 8248
rect 13688 8276 13694 8288
rect 13786 8276 13814 8384
rect 14185 8381 14197 8384
rect 14231 8412 14243 8415
rect 14645 8415 14703 8421
rect 14645 8412 14657 8415
rect 14231 8384 14657 8412
rect 14231 8381 14243 8384
rect 14185 8375 14243 8381
rect 14645 8381 14657 8384
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 15289 8415 15347 8421
rect 15289 8381 15301 8415
rect 15335 8381 15347 8415
rect 15746 8412 15752 8424
rect 15707 8384 15752 8412
rect 15289 8375 15347 8381
rect 15746 8372 15752 8384
rect 15804 8412 15810 8424
rect 16301 8415 16359 8421
rect 16301 8412 16313 8415
rect 15804 8384 16313 8412
rect 15804 8372 15810 8384
rect 16301 8381 16313 8384
rect 16347 8381 16359 8415
rect 16301 8375 16359 8381
rect 23382 8372 23388 8424
rect 23440 8412 23446 8424
rect 23753 8415 23811 8421
rect 23753 8412 23765 8415
rect 23440 8384 23765 8412
rect 23440 8372 23446 8384
rect 23753 8381 23765 8384
rect 23799 8381 23811 8415
rect 23753 8375 23811 8381
rect 16025 8347 16083 8353
rect 16025 8313 16037 8347
rect 16071 8344 16083 8347
rect 16666 8344 16672 8356
rect 16071 8316 16672 8344
rect 16071 8313 16083 8316
rect 16025 8307 16083 8313
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 18138 8304 18144 8356
rect 18196 8344 18202 8356
rect 18233 8347 18291 8353
rect 18233 8344 18245 8347
rect 18196 8316 18245 8344
rect 18196 8304 18202 8316
rect 18233 8313 18245 8316
rect 18279 8313 18291 8347
rect 18233 8307 18291 8313
rect 23934 8304 23940 8356
rect 23992 8344 23998 8356
rect 25041 8347 25099 8353
rect 25041 8344 25053 8347
rect 23992 8316 25053 8344
rect 23992 8304 23998 8316
rect 25041 8313 25053 8316
rect 25087 8313 25099 8347
rect 25041 8307 25099 8313
rect 13688 8248 13814 8276
rect 13688 8236 13694 8248
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 7190 8072 7196 8084
rect 7151 8044 7196 8072
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 8754 8072 8760 8084
rect 8715 8044 8760 8072
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 11146 8072 11152 8084
rect 9907 8044 11152 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 11146 8032 11152 8044
rect 11204 8072 11210 8084
rect 11333 8075 11391 8081
rect 11333 8072 11345 8075
rect 11204 8044 11345 8072
rect 11204 8032 11210 8044
rect 11333 8041 11345 8044
rect 11379 8041 11391 8075
rect 11333 8035 11391 8041
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12805 8075 12863 8081
rect 12805 8072 12817 8075
rect 12676 8044 12817 8072
rect 12676 8032 12682 8044
rect 12805 8041 12817 8044
rect 12851 8041 12863 8075
rect 12805 8035 12863 8041
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 15746 8072 15752 8084
rect 15611 8044 15752 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 23934 8032 23940 8084
rect 23992 8072 23998 8084
rect 24259 8075 24317 8081
rect 24259 8072 24271 8075
rect 23992 8044 24271 8072
rect 23992 8032 23998 8044
rect 24259 8041 24271 8044
rect 24305 8041 24317 8075
rect 24259 8035 24317 8041
rect 11974 8004 11980 8016
rect 11935 7976 11980 8004
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 15470 7964 15476 8016
rect 15528 8004 15534 8016
rect 15841 8007 15899 8013
rect 15841 8004 15853 8007
rect 15528 7976 15853 8004
rect 15528 7964 15534 7976
rect 15841 7973 15853 7976
rect 15887 7973 15899 8007
rect 15841 7967 15899 7973
rect 16390 7964 16396 8016
rect 16448 8004 16454 8016
rect 16622 8007 16680 8013
rect 16622 8004 16634 8007
rect 16448 7976 16634 8004
rect 16448 7964 16454 7976
rect 16622 7973 16634 7976
rect 16668 7973 16680 8007
rect 16622 7967 16680 7973
rect 6181 7939 6239 7945
rect 6181 7905 6193 7939
rect 6227 7936 6239 7939
rect 6270 7936 6276 7948
rect 6227 7908 6276 7936
rect 6227 7905 6239 7908
rect 6181 7899 6239 7905
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8018 7936 8024 7948
rect 7883 7908 8024 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 6546 7868 6552 7880
rect 6144 7840 6552 7868
rect 6144 7828 6150 7840
rect 6546 7828 6552 7840
rect 6604 7868 6610 7880
rect 7852 7868 7880 7899
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 10686 7936 10692 7948
rect 10599 7908 10692 7936
rect 10686 7896 10692 7908
rect 10744 7936 10750 7948
rect 11606 7936 11612 7948
rect 10744 7908 11612 7936
rect 10744 7896 10750 7908
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 12526 7896 12532 7948
rect 12584 7936 12590 7948
rect 12802 7936 12808 7948
rect 12584 7908 12808 7936
rect 12584 7896 12590 7908
rect 12802 7896 12808 7908
rect 12860 7896 12866 7948
rect 13446 7936 13452 7948
rect 13407 7908 13452 7936
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 16022 7896 16028 7948
rect 16080 7936 16086 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 16080 7908 16313 7936
rect 16080 7896 16086 7908
rect 16301 7905 16313 7908
rect 16347 7905 16359 7939
rect 16301 7899 16359 7905
rect 17221 7939 17279 7945
rect 17221 7905 17233 7939
rect 17267 7936 17279 7939
rect 18230 7936 18236 7948
rect 17267 7908 18236 7936
rect 17267 7905 17279 7908
rect 17221 7899 17279 7905
rect 18230 7896 18236 7908
rect 18288 7896 18294 7948
rect 24188 7939 24246 7945
rect 24188 7905 24200 7939
rect 24234 7936 24246 7939
rect 24762 7936 24768 7948
rect 24234 7908 24768 7936
rect 24234 7905 24246 7908
rect 24188 7899 24246 7905
rect 24762 7896 24768 7908
rect 24820 7896 24826 7948
rect 8478 7868 8484 7880
rect 6604 7840 7880 7868
rect 8439 7840 8484 7868
rect 6604 7828 6610 7840
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 11885 7871 11943 7877
rect 11885 7868 11897 7871
rect 11388 7840 11897 7868
rect 11388 7828 11394 7840
rect 11885 7837 11897 7840
rect 11931 7868 11943 7871
rect 12158 7868 12164 7880
rect 11931 7840 12164 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 13354 7868 13360 7880
rect 13315 7840 13360 7868
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 6346 7803 6404 7809
rect 6346 7769 6358 7803
rect 6392 7800 6404 7803
rect 7006 7800 7012 7812
rect 6392 7772 7012 7800
rect 6392 7769 6404 7772
rect 6346 7763 6404 7769
rect 7006 7760 7012 7772
rect 7064 7760 7070 7812
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 22278 7800 22284 7812
rect 17828 7772 22284 7800
rect 17828 7760 17834 7772
rect 22278 7760 22284 7772
rect 22336 7760 22342 7812
rect 6457 7735 6515 7741
rect 6457 7701 6469 7735
rect 6503 7732 6515 7735
rect 6638 7732 6644 7744
rect 6503 7704 6644 7732
rect 6503 7701 6515 7704
rect 6457 7695 6515 7701
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 6822 7732 6828 7744
rect 6783 7704 6828 7732
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7732 7622 7744
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 7616 7704 9137 7732
rect 7616 7692 7622 7704
rect 9125 7701 9137 7704
rect 9171 7701 9183 7735
rect 9125 7695 9183 7701
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 10965 7735 11023 7741
rect 10965 7732 10977 7735
rect 10928 7704 10977 7732
rect 10928 7692 10934 7704
rect 10965 7701 10977 7704
rect 11011 7701 11023 7735
rect 18322 7732 18328 7744
rect 18283 7704 18328 7732
rect 10965 7695 11023 7701
rect 18322 7692 18328 7704
rect 18380 7692 18386 7744
rect 23750 7732 23756 7744
rect 23711 7704 23756 7732
rect 23750 7692 23756 7704
rect 23808 7692 23814 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 9309 7531 9367 7537
rect 9309 7528 9321 7531
rect 6880 7500 9321 7528
rect 6880 7488 6886 7500
rect 9309 7497 9321 7500
rect 9355 7528 9367 7531
rect 9674 7528 9680 7540
rect 9355 7500 9680 7528
rect 9355 7497 9367 7500
rect 9309 7491 9367 7497
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 10686 7528 10692 7540
rect 10647 7500 10692 7528
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 11974 7528 11980 7540
rect 11931 7500 11980 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 12158 7528 12164 7540
rect 12119 7500 12164 7528
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 13446 7528 13452 7540
rect 13407 7500 13452 7528
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 16022 7488 16028 7540
rect 16080 7528 16086 7540
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 16080 7500 16681 7528
rect 16080 7488 16086 7500
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 16669 7491 16727 7497
rect 17402 7488 17408 7500
rect 17460 7528 17466 7540
rect 17460 7500 18184 7528
rect 17460 7488 17466 7500
rect 6273 7463 6331 7469
rect 6273 7429 6285 7463
rect 6319 7460 6331 7463
rect 6638 7460 6644 7472
rect 6319 7432 6644 7460
rect 6319 7429 6331 7432
rect 6273 7423 6331 7429
rect 6638 7420 6644 7432
rect 6696 7460 6702 7472
rect 7561 7463 7619 7469
rect 7561 7460 7573 7463
rect 6696 7432 7573 7460
rect 6696 7420 6702 7432
rect 7561 7429 7573 7432
rect 7607 7429 7619 7463
rect 7561 7423 7619 7429
rect 1535 7395 1593 7401
rect 1535 7361 1547 7395
rect 1581 7392 1593 7395
rect 8938 7392 8944 7404
rect 1581 7364 8944 7392
rect 1581 7361 1593 7364
rect 1535 7355 1593 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13722 7392 13728 7404
rect 13679 7364 13728 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 14090 7392 14096 7404
rect 14051 7364 14096 7392
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 18156 7401 18184 7500
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7361 18199 7395
rect 18506 7392 18512 7404
rect 18467 7364 18512 7392
rect 18141 7355 18199 7361
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 23750 7392 23756 7404
rect 23446 7364 23756 7392
rect 106 7284 112 7336
rect 164 7324 170 7336
rect 1432 7327 1490 7333
rect 1432 7324 1444 7327
rect 164 7296 1444 7324
rect 164 7284 170 7296
rect 1432 7293 1444 7296
rect 1478 7324 1490 7327
rect 1857 7327 1915 7333
rect 1857 7324 1869 7327
rect 1478 7296 1869 7324
rect 1478 7293 1490 7296
rect 1432 7287 1490 7293
rect 1857 7293 1869 7296
rect 1903 7293 1915 7327
rect 1857 7287 1915 7293
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 6546 7324 6552 7336
rect 5132 7296 6552 7324
rect 5132 7284 5138 7296
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 7190 7284 7196 7336
rect 7248 7324 7254 7336
rect 7926 7324 7932 7336
rect 7248 7296 7932 7324
rect 7248 7284 7254 7296
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 8386 7324 8392 7336
rect 8347 7296 8392 7324
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 8478 7284 8484 7336
rect 8536 7324 8542 7336
rect 9493 7327 9551 7333
rect 9493 7324 9505 7327
rect 8536 7296 9505 7324
rect 8536 7284 8542 7296
rect 9493 7293 9505 7296
rect 9539 7324 9551 7327
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9539 7296 9965 7324
rect 9539 7293 9551 7296
rect 9493 7287 9551 7293
rect 9953 7293 9965 7296
rect 9999 7324 10011 7327
rect 10042 7324 10048 7336
rect 9999 7296 10048 7324
rect 9999 7293 10011 7296
rect 9953 7287 10011 7293
rect 10042 7284 10048 7296
rect 10100 7284 10106 7336
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 10744 7296 10793 7324
rect 10744 7284 10750 7296
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 11238 7324 11244 7336
rect 11199 7296 11244 7324
rect 10781 7287 10839 7293
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14884 7296 15117 7324
rect 14884 7284 14890 7296
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7293 15623 7327
rect 15565 7287 15623 7293
rect 5905 7259 5963 7265
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 6270 7256 6276 7268
rect 5951 7228 6276 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 6270 7216 6276 7228
rect 6328 7216 6334 7268
rect 6564 7256 6592 7284
rect 7377 7259 7435 7265
rect 7377 7256 7389 7259
rect 6564 7228 7389 7256
rect 7377 7225 7389 7228
rect 7423 7225 7435 7259
rect 7377 7219 7435 7225
rect 7561 7259 7619 7265
rect 7561 7225 7573 7259
rect 7607 7256 7619 7259
rect 7837 7259 7895 7265
rect 7837 7256 7849 7259
rect 7607 7228 7849 7256
rect 7607 7225 7619 7228
rect 7561 7219 7619 7225
rect 7837 7225 7849 7228
rect 7883 7256 7895 7259
rect 8404 7256 8432 7284
rect 11514 7256 11520 7268
rect 7883 7228 8432 7256
rect 11475 7228 11520 7256
rect 7883 7225 7895 7228
rect 7837 7219 7895 7225
rect 11514 7216 11520 7228
rect 11572 7216 11578 7268
rect 13725 7259 13783 7265
rect 13725 7225 13737 7259
rect 13771 7225 13783 7259
rect 14642 7256 14648 7268
rect 14555 7228 14648 7256
rect 13725 7219 13783 7225
rect 7006 7188 7012 7200
rect 6967 7160 7012 7188
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 9398 7148 9404 7200
rect 9456 7188 9462 7200
rect 9677 7191 9735 7197
rect 9677 7188 9689 7191
rect 9456 7160 9689 7188
rect 9456 7148 9462 7160
rect 9677 7157 9689 7160
rect 9723 7157 9735 7191
rect 9677 7151 9735 7157
rect 13081 7191 13139 7197
rect 13081 7157 13093 7191
rect 13127 7188 13139 7191
rect 13446 7188 13452 7200
rect 13127 7160 13452 7188
rect 13127 7157 13139 7160
rect 13081 7151 13139 7157
rect 13446 7148 13452 7160
rect 13504 7188 13510 7200
rect 13740 7188 13768 7219
rect 14642 7216 14648 7228
rect 14700 7256 14706 7268
rect 15580 7256 15608 7287
rect 14700 7228 15608 7256
rect 14700 7216 14706 7228
rect 18230 7216 18236 7268
rect 18288 7256 18294 7268
rect 18288 7228 18333 7256
rect 18288 7216 18294 7228
rect 22094 7216 22100 7268
rect 22152 7256 22158 7268
rect 23446 7256 23474 7364
rect 23750 7352 23756 7364
rect 23808 7352 23814 7404
rect 23934 7352 23940 7404
rect 23992 7392 23998 7404
rect 24029 7395 24087 7401
rect 24029 7392 24041 7395
rect 23992 7364 24041 7392
rect 23992 7352 23998 7364
rect 24029 7361 24041 7364
rect 24075 7361 24087 7395
rect 24029 7355 24087 7361
rect 23842 7256 23848 7268
rect 22152 7228 23474 7256
rect 23803 7228 23848 7256
rect 22152 7216 22158 7228
rect 23842 7216 23848 7228
rect 23900 7216 23906 7268
rect 13504 7160 13768 7188
rect 13504 7148 13510 7160
rect 14826 7148 14832 7200
rect 14884 7188 14890 7200
rect 14921 7191 14979 7197
rect 14921 7188 14933 7191
rect 14884 7160 14933 7188
rect 14884 7148 14890 7160
rect 14921 7157 14933 7160
rect 14967 7157 14979 7191
rect 15378 7188 15384 7200
rect 15339 7160 15384 7188
rect 14921 7151 14979 7157
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 16298 7188 16304 7200
rect 16259 7160 16304 7188
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 17865 7191 17923 7197
rect 17865 7157 17877 7191
rect 17911 7188 17923 7191
rect 18248 7188 18276 7216
rect 17911 7160 18276 7188
rect 23477 7191 23535 7197
rect 17911 7157 17923 7160
rect 17865 7151 17923 7157
rect 23477 7157 23489 7191
rect 23523 7188 23535 7191
rect 23860 7188 23888 7216
rect 24762 7188 24768 7200
rect 23523 7160 23888 7188
rect 24675 7160 24768 7188
rect 23523 7157 23535 7160
rect 23477 7151 23535 7157
rect 24762 7148 24768 7160
rect 24820 7188 24826 7200
rect 25498 7188 25504 7200
rect 24820 7160 25504 7188
rect 24820 7148 24826 7160
rect 25498 7148 25504 7160
rect 25556 7148 25562 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 7926 6944 7932 6996
rect 7984 6984 7990 6996
rect 8386 6984 8392 6996
rect 7984 6956 8392 6984
rect 7984 6944 7990 6956
rect 8386 6944 8392 6956
rect 8444 6984 8450 6996
rect 8665 6987 8723 6993
rect 8665 6984 8677 6987
rect 8444 6956 8677 6984
rect 8444 6944 8450 6956
rect 8665 6953 8677 6956
rect 8711 6953 8723 6987
rect 8665 6947 8723 6953
rect 10321 6987 10379 6993
rect 10321 6953 10333 6987
rect 10367 6984 10379 6987
rect 11238 6984 11244 6996
rect 10367 6956 11244 6984
rect 10367 6953 10379 6956
rect 10321 6947 10379 6953
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 13173 6987 13231 6993
rect 13173 6953 13185 6987
rect 13219 6984 13231 6987
rect 13446 6984 13452 6996
rect 13219 6956 13452 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 13633 6987 13691 6993
rect 13633 6953 13645 6987
rect 13679 6984 13691 6987
rect 13722 6984 13728 6996
rect 13679 6956 13728 6984
rect 13679 6953 13691 6956
rect 13633 6947 13691 6953
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 15378 6944 15384 6996
rect 15436 6984 15442 6996
rect 15565 6987 15623 6993
rect 15565 6984 15577 6987
rect 15436 6956 15577 6984
rect 15436 6944 15442 6956
rect 15565 6953 15577 6956
rect 15611 6953 15623 6987
rect 15565 6947 15623 6953
rect 18141 6987 18199 6993
rect 18141 6953 18153 6987
rect 18187 6984 18199 6987
rect 18230 6984 18236 6996
rect 18187 6956 18236 6984
rect 18187 6953 18199 6956
rect 18141 6947 18199 6953
rect 18230 6944 18236 6956
rect 18288 6944 18294 6996
rect 18340 6956 18644 6984
rect 7006 6876 7012 6928
rect 7064 6916 7070 6928
rect 7064 6888 8248 6916
rect 7064 6876 7070 6888
rect 6178 6848 6184 6860
rect 6139 6820 6184 6848
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6270 6808 6276 6860
rect 6328 6848 6334 6860
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 6328 6820 6837 6848
rect 6328 6808 6334 6820
rect 6825 6817 6837 6820
rect 6871 6848 6883 6851
rect 7650 6848 7656 6860
rect 6871 6820 7656 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 8220 6857 8248 6888
rect 11882 6876 11888 6928
rect 11940 6916 11946 6928
rect 12574 6919 12632 6925
rect 12574 6916 12586 6919
rect 11940 6888 12586 6916
rect 11940 6876 11946 6888
rect 12574 6885 12586 6888
rect 12620 6885 12632 6919
rect 12574 6879 12632 6885
rect 16298 6876 16304 6928
rect 16356 6916 16362 6928
rect 16990 6919 17048 6925
rect 16990 6916 17002 6919
rect 16356 6888 17002 6916
rect 16356 6876 16362 6888
rect 16990 6885 17002 6888
rect 17036 6885 17048 6919
rect 18340 6916 18368 6956
rect 18506 6916 18512 6928
rect 16990 6879 17048 6885
rect 18248 6888 18368 6916
rect 18467 6888 18512 6916
rect 18248 6860 18276 6888
rect 18506 6876 18512 6888
rect 18564 6876 18570 6928
rect 18616 6925 18644 6956
rect 22830 6944 22836 6996
rect 22888 6984 22894 6996
rect 22888 6956 22968 6984
rect 22888 6944 22894 6956
rect 18601 6919 18659 6925
rect 18601 6885 18613 6919
rect 18647 6916 18659 6919
rect 19610 6916 19616 6928
rect 18647 6888 19616 6916
rect 18647 6885 18659 6888
rect 18601 6879 18659 6885
rect 19610 6876 19616 6888
rect 19668 6876 19674 6928
rect 22940 6925 22968 6956
rect 22925 6919 22983 6925
rect 22925 6885 22937 6919
rect 22971 6885 22983 6919
rect 22925 6879 22983 6885
rect 23014 6876 23020 6928
rect 23072 6916 23078 6928
rect 23072 6888 23117 6916
rect 23072 6876 23078 6888
rect 23842 6876 23848 6928
rect 23900 6916 23906 6928
rect 24397 6919 24455 6925
rect 24397 6916 24409 6919
rect 23900 6888 24409 6916
rect 23900 6876 23906 6888
rect 24397 6885 24409 6888
rect 24443 6885 24455 6919
rect 24397 6879 24455 6885
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6817 8263 6851
rect 9674 6848 9680 6860
rect 9635 6820 9680 6848
rect 8205 6811 8263 6817
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 16666 6848 16672 6860
rect 16627 6820 16672 6848
rect 16666 6808 16672 6820
rect 16724 6808 16730 6860
rect 17589 6851 17647 6857
rect 17589 6817 17601 6851
rect 17635 6848 17647 6851
rect 18230 6848 18236 6860
rect 17635 6820 18236 6848
rect 17635 6817 17647 6820
rect 17589 6811 17647 6817
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 24670 6848 24676 6860
rect 24631 6820 24676 6848
rect 24670 6808 24676 6820
rect 24728 6808 24734 6860
rect 7098 6740 7104 6792
rect 7156 6780 7162 6792
rect 7193 6783 7251 6789
rect 7193 6780 7205 6783
rect 7156 6752 7205 6780
rect 7156 6740 7162 6752
rect 7193 6749 7205 6752
rect 7239 6780 7251 6783
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7239 6752 7573 6780
rect 7239 6749 7251 6752
rect 7193 6743 7251 6749
rect 7561 6749 7573 6752
rect 7607 6780 7619 6783
rect 8018 6780 8024 6792
rect 7607 6752 8024 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 10042 6780 10048 6792
rect 10003 6752 10048 6780
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 11514 6740 11520 6792
rect 11572 6780 11578 6792
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 11572 6752 12265 6780
rect 11572 6740 11578 6752
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 13998 6780 14004 6792
rect 13959 6752 14004 6780
rect 12253 6743 12311 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 19150 6780 19156 6792
rect 19111 6752 19156 6780
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6780 23627 6783
rect 24026 6780 24032 6792
rect 23615 6752 24032 6780
rect 23615 6749 23627 6752
rect 23569 6743 23627 6749
rect 24026 6740 24032 6752
rect 24084 6740 24090 6792
rect 8386 6672 8392 6724
rect 8444 6712 8450 6724
rect 9950 6712 9956 6724
rect 8444 6684 9956 6712
rect 8444 6672 8450 6684
rect 9950 6672 9956 6684
rect 10008 6672 10014 6724
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 9815 6647 9873 6653
rect 9815 6644 9827 6647
rect 9548 6616 9827 6644
rect 9548 6604 9554 6616
rect 9815 6613 9827 6616
rect 9861 6613 9873 6647
rect 10870 6644 10876 6656
rect 10831 6616 10876 6644
rect 9815 6607 9873 6613
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 23842 6644 23848 6656
rect 23803 6616 23848 6644
rect 23842 6604 23848 6616
rect 23900 6604 23906 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8278 6443 8336 6449
rect 8278 6440 8290 6443
rect 8076 6412 8290 6440
rect 8076 6400 8082 6412
rect 8278 6409 8290 6412
rect 8324 6440 8336 6443
rect 9490 6440 9496 6452
rect 8324 6412 9496 6440
rect 8324 6409 8336 6412
rect 8278 6403 8336 6409
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10100 6412 10425 6440
rect 10100 6400 10106 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 10413 6403 10471 6409
rect 11514 6400 11520 6452
rect 11572 6440 11578 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11572 6412 11805 6440
rect 11572 6400 11578 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 13354 6440 13360 6452
rect 13315 6412 13360 6440
rect 11793 6403 11851 6409
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 14826 6440 14832 6452
rect 13648 6412 14832 6440
rect 8386 6372 8392 6384
rect 8347 6344 8392 6372
rect 8386 6332 8392 6344
rect 8444 6332 8450 6384
rect 10870 6372 10876 6384
rect 10783 6344 10876 6372
rect 8478 6304 8484 6316
rect 8439 6276 8484 6304
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 9950 6264 9956 6316
rect 10008 6304 10014 6316
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 10008 6276 10057 6304
rect 10008 6264 10014 6276
rect 10045 6273 10057 6276
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 7098 6236 7104 6248
rect 7059 6208 7104 6236
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 8018 6196 8024 6248
rect 8076 6236 8082 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 8076 6208 8125 6236
rect 8076 6196 8082 6208
rect 8113 6205 8125 6208
rect 8159 6236 8171 6239
rect 8754 6236 8760 6248
rect 8159 6208 8760 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8754 6196 8760 6208
rect 8812 6236 8818 6248
rect 10796 6245 10824 6344
rect 10870 6332 10876 6344
rect 10928 6372 10934 6384
rect 12621 6375 12679 6381
rect 12621 6372 12633 6375
rect 10928 6344 12633 6372
rect 10928 6332 10934 6344
rect 12621 6341 12633 6344
rect 12667 6372 12679 6375
rect 13648 6372 13676 6412
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 16666 6400 16672 6452
rect 16724 6440 16730 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 16724 6412 17141 6440
rect 16724 6400 16730 6412
rect 17129 6409 17141 6412
rect 17175 6409 17187 6443
rect 19610 6440 19616 6452
rect 17129 6403 17187 6409
rect 18800 6412 19472 6440
rect 19571 6412 19616 6440
rect 14090 6372 14096 6384
rect 12667 6344 13676 6372
rect 14051 6344 14096 6372
rect 12667 6341 12679 6344
rect 12621 6335 12679 6341
rect 14090 6332 14096 6344
rect 14148 6372 14154 6384
rect 16485 6375 16543 6381
rect 14148 6344 16436 6372
rect 14148 6332 14154 6344
rect 13538 6264 13544 6316
rect 13596 6304 13602 6316
rect 13998 6304 14004 6316
rect 13596 6276 14004 6304
rect 13596 6264 13602 6276
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 15378 6264 15384 6316
rect 15436 6304 15442 6316
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 15436 6276 15577 6304
rect 15436 6264 15442 6276
rect 15565 6273 15577 6276
rect 15611 6273 15623 6307
rect 16408 6304 16436 6344
rect 16485 6341 16497 6375
rect 16531 6372 16543 6375
rect 18800 6372 18828 6412
rect 16531 6344 18828 6372
rect 16531 6341 16543 6344
rect 16485 6335 16543 6341
rect 19150 6332 19156 6384
rect 19208 6372 19214 6384
rect 19245 6375 19303 6381
rect 19245 6372 19257 6375
rect 19208 6344 19257 6372
rect 19208 6332 19214 6344
rect 19245 6341 19257 6344
rect 19291 6341 19303 6375
rect 19444 6372 19472 6412
rect 19610 6400 19616 6412
rect 19668 6400 19674 6452
rect 24670 6440 24676 6452
rect 23446 6412 24676 6440
rect 23446 6384 23474 6412
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 25409 6443 25467 6449
rect 25409 6409 25421 6443
rect 25455 6440 25467 6443
rect 25590 6440 25596 6452
rect 25455 6412 25596 6440
rect 25455 6409 25467 6412
rect 25409 6403 25467 6409
rect 25590 6400 25596 6412
rect 25648 6400 25654 6452
rect 21821 6375 21879 6381
rect 21821 6372 21833 6375
rect 19444 6344 21833 6372
rect 19245 6335 19303 6341
rect 21821 6341 21833 6344
rect 21867 6341 21879 6375
rect 21821 6335 21879 6341
rect 17586 6304 17592 6316
rect 16408 6276 17592 6304
rect 15565 6267 15623 6273
rect 17586 6264 17592 6276
rect 17644 6264 17650 6316
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 17911 6276 18705 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 18693 6273 18705 6276
rect 18739 6304 18751 6307
rect 20165 6307 20223 6313
rect 20165 6304 20177 6307
rect 18739 6276 20177 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 20165 6273 20177 6276
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8812 6208 9137 6236
rect 8812 6196 8818 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 10781 6239 10839 6245
rect 10781 6205 10793 6239
rect 10827 6205 10839 6239
rect 10781 6199 10839 6205
rect 10962 6196 10968 6248
rect 11020 6236 11026 6248
rect 11241 6239 11299 6245
rect 11241 6236 11253 6239
rect 11020 6208 11253 6236
rect 11020 6196 11026 6208
rect 11241 6205 11253 6208
rect 11287 6205 11299 6239
rect 11241 6199 11299 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 21836 6236 21864 6335
rect 23382 6332 23388 6384
rect 23440 6344 23474 6384
rect 23440 6332 23446 6344
rect 22741 6307 22799 6313
rect 22741 6273 22753 6307
rect 22787 6304 22799 6307
rect 23477 6307 23535 6313
rect 23477 6304 23489 6307
rect 22787 6276 23489 6304
rect 22787 6273 22799 6276
rect 22741 6267 22799 6273
rect 23477 6273 23489 6276
rect 23523 6273 23535 6307
rect 23477 6267 23535 6273
rect 23753 6307 23811 6313
rect 23753 6273 23765 6307
rect 23799 6304 23811 6307
rect 23842 6304 23848 6316
rect 23799 6276 23848 6304
rect 23799 6273 23811 6276
rect 23753 6267 23811 6273
rect 22097 6239 22155 6245
rect 22097 6236 22109 6239
rect 12483 6208 13032 6236
rect 21836 6208 22109 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 6638 6128 6644 6180
rect 6696 6168 6702 6180
rect 7006 6168 7012 6180
rect 6696 6140 7012 6168
rect 6696 6128 6702 6140
rect 7006 6128 7012 6140
rect 7064 6168 7070 6180
rect 7653 6171 7711 6177
rect 7653 6168 7665 6171
rect 7064 6140 7665 6168
rect 7064 6128 7070 6140
rect 7653 6137 7665 6140
rect 7699 6137 7711 6171
rect 7653 6131 7711 6137
rect 8849 6171 8907 6177
rect 8849 6137 8861 6171
rect 8895 6168 8907 6171
rect 12710 6168 12716 6180
rect 8895 6140 12716 6168
rect 8895 6137 8907 6140
rect 8849 6131 8907 6137
rect 12710 6128 12716 6140
rect 12768 6128 12774 6180
rect 13004 6112 13032 6208
rect 22097 6205 22109 6208
rect 22143 6236 22155 6239
rect 23014 6236 23020 6248
rect 22143 6208 23020 6236
rect 22143 6205 22155 6208
rect 22097 6199 22155 6205
rect 23014 6196 23020 6208
rect 23072 6196 23078 6248
rect 13538 6168 13544 6180
rect 13499 6140 13544 6168
rect 13538 6128 13544 6140
rect 13596 6128 13602 6180
rect 13633 6171 13691 6177
rect 13633 6137 13645 6171
rect 13679 6137 13691 6171
rect 15886 6171 15944 6177
rect 15886 6168 15898 6171
rect 13633 6131 13691 6137
rect 15488 6140 15898 6168
rect 6178 6100 6184 6112
rect 6139 6072 6184 6100
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 7285 6103 7343 6109
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 7558 6100 7564 6112
rect 7331 6072 7564 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 7558 6060 7564 6072
rect 7616 6100 7622 6112
rect 8110 6100 8116 6112
rect 7616 6072 8116 6100
rect 7616 6060 7622 6072
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8386 6100 8392 6112
rect 8260 6072 8392 6100
rect 8260 6060 8266 6072
rect 8386 6060 8392 6072
rect 8444 6100 8450 6112
rect 9674 6100 9680 6112
rect 8444 6072 9680 6100
rect 8444 6060 8450 6072
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 11054 6100 11060 6112
rect 11015 6072 11060 6100
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 11940 6072 12173 6100
rect 11940 6060 11946 6072
rect 12161 6069 12173 6072
rect 12207 6069 12219 6103
rect 12986 6100 12992 6112
rect 12947 6072 12992 6100
rect 12161 6063 12219 6069
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 13354 6060 13360 6112
rect 13412 6100 13418 6112
rect 13648 6100 13676 6131
rect 15488 6112 15516 6140
rect 15886 6137 15898 6140
rect 15932 6168 15944 6171
rect 16298 6168 16304 6180
rect 15932 6140 16304 6168
rect 15932 6137 15944 6140
rect 15886 6131 15944 6137
rect 16298 6128 16304 6140
rect 16356 6168 16362 6180
rect 16761 6171 16819 6177
rect 16761 6168 16773 6171
rect 16356 6140 16773 6168
rect 16356 6128 16362 6140
rect 16761 6137 16773 6140
rect 16807 6137 16819 6171
rect 16761 6131 16819 6137
rect 18785 6171 18843 6177
rect 18785 6137 18797 6171
rect 18831 6137 18843 6171
rect 23492 6168 23520 6267
rect 23842 6264 23848 6276
rect 23900 6264 23906 6316
rect 24026 6304 24032 6316
rect 23987 6276 24032 6304
rect 24026 6264 24032 6276
rect 24084 6264 24090 6316
rect 25222 6236 25228 6248
rect 25135 6208 25228 6236
rect 25222 6196 25228 6208
rect 25280 6236 25286 6248
rect 25777 6239 25835 6245
rect 25777 6236 25789 6239
rect 25280 6208 25789 6236
rect 25280 6196 25286 6208
rect 25777 6205 25789 6208
rect 25823 6205 25835 6239
rect 25777 6199 25835 6205
rect 23845 6171 23903 6177
rect 23845 6168 23857 6171
rect 23492 6140 23857 6168
rect 18785 6131 18843 6137
rect 23845 6137 23857 6140
rect 23891 6137 23903 6171
rect 23845 6131 23903 6137
rect 15470 6100 15476 6112
rect 13412 6072 13676 6100
rect 15431 6072 15476 6100
rect 13412 6060 13418 6072
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 18414 6100 18420 6112
rect 18375 6072 18420 6100
rect 18414 6060 18420 6072
rect 18472 6100 18478 6112
rect 18800 6100 18828 6131
rect 18472 6072 18828 6100
rect 18472 6060 18478 6072
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 6825 5899 6883 5905
rect 6825 5865 6837 5899
rect 6871 5896 6883 5899
rect 6914 5896 6920 5908
rect 6871 5868 6920 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7561 5899 7619 5905
rect 7561 5865 7573 5899
rect 7607 5896 7619 5899
rect 7650 5896 7656 5908
rect 7607 5868 7656 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 7929 5899 7987 5905
rect 7929 5865 7941 5899
rect 7975 5896 7987 5899
rect 8478 5896 8484 5908
rect 7975 5868 8484 5896
rect 7975 5865 7987 5868
rect 7929 5859 7987 5865
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 9490 5896 9496 5908
rect 9451 5868 9496 5896
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 13538 5896 13544 5908
rect 11664 5868 12388 5896
rect 13499 5868 13544 5896
rect 11664 5856 11670 5868
rect 8018 5828 8024 5840
rect 7979 5800 8024 5828
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 9950 5788 9956 5840
rect 10008 5828 10014 5840
rect 10182 5831 10240 5837
rect 10182 5828 10194 5831
rect 10008 5800 10194 5828
rect 10008 5788 10014 5800
rect 10182 5797 10194 5800
rect 10228 5797 10240 5831
rect 11790 5828 11796 5840
rect 11751 5800 11796 5828
rect 10182 5791 10240 5797
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 6236 5732 6561 5760
rect 6236 5720 6242 5732
rect 6549 5729 6561 5732
rect 6595 5729 6607 5763
rect 6549 5723 6607 5729
rect 6638 5720 6644 5772
rect 6696 5760 6702 5772
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6696 5732 6745 5760
rect 6696 5720 6702 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 9398 5760 9404 5772
rect 6733 5723 6791 5729
rect 8404 5732 9404 5760
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 8404 5701 8432 5732
rect 9398 5720 9404 5732
rect 9456 5720 9462 5772
rect 9858 5760 9864 5772
rect 9819 5732 9864 5760
rect 9858 5720 9864 5732
rect 9916 5720 9922 5772
rect 12360 5760 12388 5868
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 16577 5899 16635 5905
rect 16577 5865 16589 5899
rect 16623 5896 16635 5899
rect 22094 5896 22100 5908
rect 16623 5868 19748 5896
rect 22055 5868 22100 5896
rect 16623 5865 16635 5868
rect 16577 5859 16635 5865
rect 12986 5788 12992 5840
rect 13044 5828 13050 5840
rect 13722 5828 13728 5840
rect 13044 5800 13728 5828
rect 13044 5788 13050 5800
rect 13722 5788 13728 5800
rect 13780 5788 13786 5840
rect 15470 5788 15476 5840
rect 15528 5828 15534 5840
rect 15978 5831 16036 5837
rect 15978 5828 15990 5831
rect 15528 5800 15990 5828
rect 15528 5788 15534 5800
rect 15978 5797 15990 5800
rect 16024 5797 16036 5831
rect 15978 5791 16036 5797
rect 18322 5788 18328 5840
rect 18380 5828 18386 5840
rect 18417 5831 18475 5837
rect 18417 5828 18429 5831
rect 18380 5800 18429 5828
rect 18380 5788 18386 5800
rect 18417 5797 18429 5800
rect 18463 5797 18475 5831
rect 19720 5828 19748 5868
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 22830 5896 22836 5908
rect 22791 5868 22836 5896
rect 22830 5856 22836 5868
rect 22888 5856 22894 5908
rect 24811 5899 24869 5905
rect 24811 5865 24823 5899
rect 24857 5896 24869 5899
rect 25222 5896 25228 5908
rect 24857 5868 25228 5896
rect 24857 5865 24869 5868
rect 24811 5859 24869 5865
rect 25222 5856 25228 5868
rect 25280 5856 25286 5908
rect 23293 5831 23351 5837
rect 23293 5828 23305 5831
rect 19720 5800 23305 5828
rect 18417 5791 18475 5797
rect 23293 5797 23305 5800
rect 23339 5828 23351 5831
rect 23382 5828 23388 5840
rect 23339 5800 23388 5828
rect 23339 5797 23351 5800
rect 23293 5791 23351 5797
rect 23382 5788 23388 5800
rect 23440 5788 23446 5840
rect 23845 5831 23903 5837
rect 23845 5797 23857 5831
rect 23891 5828 23903 5831
rect 23934 5828 23940 5840
rect 23891 5800 23940 5828
rect 23891 5797 23903 5800
rect 23845 5791 23903 5797
rect 23934 5788 23940 5800
rect 23992 5788 23998 5840
rect 13078 5760 13084 5772
rect 12360 5732 13084 5760
rect 13078 5720 13084 5732
rect 13136 5760 13142 5772
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 13136 5732 13645 5760
rect 13136 5720 13142 5732
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 14185 5763 14243 5769
rect 14185 5729 14197 5763
rect 14231 5760 14243 5763
rect 14642 5760 14648 5772
rect 14231 5732 14648 5760
rect 14231 5729 14243 5732
rect 14185 5723 14243 5729
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 7800 5664 8401 5692
rect 7800 5652 7806 5664
rect 8389 5661 8401 5664
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5692 8815 5695
rect 9766 5692 9772 5704
rect 8803 5664 9772 5692
rect 8803 5661 8815 5664
rect 8757 5655 8815 5661
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5692 11759 5695
rect 12066 5692 12072 5704
rect 11747 5664 12072 5692
rect 11747 5661 11759 5664
rect 11701 5655 11759 5661
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 12158 5652 12164 5704
rect 12216 5692 12222 5704
rect 12216 5664 12261 5692
rect 12216 5652 12222 5664
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 14200 5692 14228 5723
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 23952 5760 23980 5788
rect 24708 5763 24766 5769
rect 24708 5760 24720 5763
rect 23952 5732 24720 5760
rect 24708 5729 24720 5732
rect 24754 5760 24766 5763
rect 25406 5760 25412 5772
rect 24754 5732 25412 5760
rect 24754 5729 24766 5732
rect 24708 5723 24766 5729
rect 25406 5720 25412 5732
rect 25464 5720 25470 5772
rect 12768 5664 14228 5692
rect 14369 5695 14427 5701
rect 12768 5652 12774 5664
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 15657 5695 15715 5701
rect 15657 5692 15669 5695
rect 14415 5664 15669 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 15657 5661 15669 5664
rect 15703 5692 15715 5695
rect 16574 5692 16580 5704
rect 15703 5664 16580 5692
rect 15703 5661 15715 5664
rect 15657 5655 15715 5661
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 8110 5584 8116 5636
rect 8168 5633 8174 5636
rect 8168 5627 8217 5633
rect 8168 5593 8171 5627
rect 8205 5593 8217 5627
rect 8294 5624 8300 5636
rect 8255 5596 8300 5624
rect 8168 5587 8217 5593
rect 8168 5584 8174 5587
rect 8294 5584 8300 5596
rect 8352 5584 8358 5636
rect 18340 5624 18368 5655
rect 18506 5652 18512 5704
rect 18564 5692 18570 5704
rect 18601 5695 18659 5701
rect 18601 5692 18613 5695
rect 18564 5664 18613 5692
rect 18564 5652 18570 5664
rect 18601 5661 18613 5664
rect 18647 5692 18659 5695
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 18647 5664 19257 5692
rect 18647 5661 18659 5664
rect 18601 5655 18659 5661
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 23201 5695 23259 5701
rect 23201 5661 23213 5695
rect 23247 5692 23259 5695
rect 24026 5692 24032 5704
rect 23247 5664 24032 5692
rect 23247 5661 23259 5664
rect 23201 5655 23259 5661
rect 24026 5652 24032 5664
rect 24084 5652 24090 5704
rect 18340 5596 18644 5624
rect 18616 5568 18644 5596
rect 9030 5556 9036 5568
rect 8991 5528 9036 5556
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 10781 5559 10839 5565
rect 10781 5556 10793 5559
rect 10744 5528 10793 5556
rect 10744 5516 10750 5528
rect 10781 5525 10793 5528
rect 10827 5525 10839 5559
rect 10781 5519 10839 5525
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 11020 5528 11069 5556
rect 11020 5516 11026 5528
rect 11057 5525 11069 5528
rect 11103 5525 11115 5559
rect 11057 5519 11115 5525
rect 18598 5516 18604 5568
rect 18656 5516 18662 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 8294 5352 8300 5364
rect 8255 5324 8300 5352
rect 8294 5312 8300 5324
rect 8352 5352 8358 5364
rect 8665 5355 8723 5361
rect 8665 5352 8677 5355
rect 8352 5324 8677 5352
rect 8352 5312 8358 5324
rect 8665 5321 8677 5324
rect 8711 5321 8723 5355
rect 9398 5352 9404 5364
rect 9359 5324 9404 5352
rect 8665 5315 8723 5321
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 11149 5355 11207 5361
rect 11149 5352 11161 5355
rect 9916 5324 11161 5352
rect 9916 5312 9922 5324
rect 11149 5321 11161 5324
rect 11195 5321 11207 5355
rect 12710 5352 12716 5364
rect 12671 5324 12716 5352
rect 11149 5315 11207 5321
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 13078 5352 13084 5364
rect 13039 5324 13084 5352
rect 13078 5312 13084 5324
rect 13136 5352 13142 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 13136 5324 13461 5352
rect 13136 5312 13142 5324
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 13449 5315 13507 5321
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 8018 5216 8024 5228
rect 7423 5188 8024 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9416 5216 9444 5312
rect 10781 5287 10839 5293
rect 10781 5253 10793 5287
rect 10827 5284 10839 5287
rect 12158 5284 12164 5296
rect 10827 5256 12164 5284
rect 10827 5253 10839 5256
rect 10781 5247 10839 5253
rect 12158 5244 12164 5256
rect 12216 5244 12222 5296
rect 8803 5188 9444 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 11609 5219 11667 5225
rect 11609 5216 11621 5219
rect 10744 5188 11621 5216
rect 10744 5176 10750 5188
rect 11609 5185 11621 5188
rect 11655 5216 11667 5219
rect 11790 5216 11796 5228
rect 11655 5188 11796 5216
rect 11655 5185 11667 5188
rect 11609 5179 11667 5185
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 12066 5216 12072 5228
rect 12027 5188 12072 5216
rect 12066 5176 12072 5188
rect 12124 5176 12130 5228
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 7009 5151 7067 5157
rect 7009 5148 7021 5151
rect 6788 5120 7021 5148
rect 6788 5108 6794 5120
rect 7009 5117 7021 5120
rect 7055 5148 7067 5151
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 7055 5120 7665 5148
rect 7055 5117 7067 5120
rect 7009 5111 7067 5117
rect 7653 5117 7665 5120
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 8110 5108 8116 5160
rect 8168 5148 8174 5160
rect 8536 5151 8594 5157
rect 8536 5148 8548 5151
rect 8168 5120 8548 5148
rect 8168 5108 8174 5120
rect 8536 5117 8548 5120
rect 8582 5148 8594 5151
rect 9030 5148 9036 5160
rect 8582 5120 9036 5148
rect 8582 5117 8594 5120
rect 8536 5111 8594 5117
rect 9030 5108 9036 5120
rect 9088 5108 9094 5160
rect 13464 5148 13492 5315
rect 15470 5312 15476 5364
rect 15528 5352 15534 5364
rect 16209 5355 16267 5361
rect 16209 5352 16221 5355
rect 15528 5324 16221 5352
rect 15528 5312 15534 5324
rect 16209 5321 16221 5324
rect 16255 5321 16267 5355
rect 16574 5352 16580 5364
rect 16535 5324 16580 5352
rect 16209 5315 16267 5321
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 18414 5352 18420 5364
rect 18375 5324 18420 5352
rect 18414 5312 18420 5324
rect 18472 5312 18478 5364
rect 22695 5355 22753 5361
rect 22695 5321 22707 5355
rect 22741 5352 22753 5355
rect 23842 5352 23848 5364
rect 22741 5324 23848 5352
rect 22741 5321 22753 5324
rect 22695 5315 22753 5321
rect 23842 5312 23848 5324
rect 23900 5312 23906 5364
rect 23937 5355 23995 5361
rect 23937 5321 23949 5355
rect 23983 5352 23995 5355
rect 24026 5352 24032 5364
rect 23983 5324 24032 5352
rect 23983 5321 23995 5324
rect 23937 5315 23995 5321
rect 24026 5312 24032 5324
rect 24084 5312 24090 5364
rect 25406 5352 25412 5364
rect 25367 5324 25412 5352
rect 25406 5312 25412 5324
rect 25464 5312 25470 5364
rect 14737 5287 14795 5293
rect 14737 5253 14749 5287
rect 14783 5284 14795 5287
rect 14826 5284 14832 5296
rect 14783 5256 14832 5284
rect 14783 5253 14795 5256
rect 14737 5247 14795 5253
rect 14826 5244 14832 5256
rect 14884 5284 14890 5296
rect 17865 5287 17923 5293
rect 14884 5256 15240 5284
rect 14884 5244 14890 5256
rect 13633 5151 13691 5157
rect 13633 5148 13645 5151
rect 13464 5120 13645 5148
rect 13633 5117 13645 5120
rect 13679 5117 13691 5151
rect 14090 5148 14096 5160
rect 14051 5120 14096 5148
rect 13633 5111 13691 5117
rect 14090 5108 14096 5120
rect 14148 5148 14154 5160
rect 15212 5157 15240 5256
rect 17865 5253 17877 5287
rect 17911 5284 17923 5287
rect 18322 5284 18328 5296
rect 17911 5256 18328 5284
rect 17911 5253 17923 5256
rect 17865 5247 17923 5253
rect 18322 5244 18328 5256
rect 18380 5244 18386 5296
rect 23382 5284 23388 5296
rect 23343 5256 23388 5284
rect 23382 5244 23388 5256
rect 23440 5244 23446 5296
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14148 5120 15025 5148
rect 14148 5108 14154 5120
rect 15013 5117 15025 5120
rect 15059 5117 15071 5151
rect 15013 5111 15071 5117
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5117 15255 5151
rect 15197 5111 15255 5117
rect 15657 5151 15715 5157
rect 15657 5117 15669 5151
rect 15703 5117 15715 5151
rect 18230 5148 18236 5160
rect 18191 5120 18236 5148
rect 15657 5111 15715 5117
rect 6822 5080 6828 5092
rect 6783 5052 6828 5080
rect 6822 5040 6828 5052
rect 6880 5040 6886 5092
rect 8386 5080 8392 5092
rect 8347 5052 8392 5080
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 9122 5080 9128 5092
rect 9083 5052 9128 5080
rect 9122 5040 9128 5052
rect 9180 5040 9186 5092
rect 10226 5080 10232 5092
rect 10187 5052 10232 5080
rect 10226 5040 10232 5052
rect 10284 5040 10290 5092
rect 10321 5083 10379 5089
rect 10321 5049 10333 5083
rect 10367 5049 10379 5083
rect 14366 5080 14372 5092
rect 14327 5052 14372 5080
rect 10321 5043 10379 5049
rect 6178 5012 6184 5024
rect 6139 4984 6184 5012
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 9858 5012 9864 5024
rect 9819 4984 9864 5012
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 9950 4972 9956 5024
rect 10008 5012 10014 5024
rect 10336 5012 10364 5043
rect 14366 5040 14372 5052
rect 14424 5040 14430 5092
rect 15028 5080 15056 5111
rect 15672 5080 15700 5111
rect 18230 5108 18236 5120
rect 18288 5108 18294 5160
rect 19150 5108 19156 5160
rect 19208 5148 19214 5160
rect 19740 5151 19798 5157
rect 19740 5148 19752 5151
rect 19208 5120 19752 5148
rect 19208 5108 19214 5120
rect 19740 5117 19752 5120
rect 19786 5148 19798 5151
rect 20165 5151 20223 5157
rect 20165 5148 20177 5151
rect 19786 5120 20177 5148
rect 19786 5117 19798 5120
rect 19740 5111 19798 5117
rect 20165 5117 20177 5120
rect 20211 5117 20223 5151
rect 20165 5111 20223 5117
rect 22624 5151 22682 5157
rect 22624 5117 22636 5151
rect 22670 5148 22682 5151
rect 24648 5151 24706 5157
rect 22670 5120 23152 5148
rect 22670 5117 22682 5120
rect 22624 5111 22682 5117
rect 23124 5089 23152 5120
rect 24648 5117 24660 5151
rect 24694 5148 24706 5151
rect 24694 5120 25176 5148
rect 24694 5117 24706 5120
rect 24648 5111 24706 5117
rect 15028 5052 15700 5080
rect 23109 5083 23167 5089
rect 23109 5049 23121 5083
rect 23155 5080 23167 5083
rect 24118 5080 24124 5092
rect 23155 5052 24124 5080
rect 23155 5049 23167 5052
rect 23109 5043 23167 5049
rect 24118 5040 24124 5052
rect 24176 5040 24182 5092
rect 25148 5089 25176 5120
rect 25133 5083 25191 5089
rect 25133 5049 25145 5083
rect 25179 5080 25191 5083
rect 27614 5080 27620 5092
rect 25179 5052 27620 5080
rect 25179 5049 25191 5052
rect 25133 5043 25191 5049
rect 27614 5040 27620 5052
rect 27672 5040 27678 5092
rect 15286 5012 15292 5024
rect 10008 4984 10364 5012
rect 15247 4984 15292 5012
rect 10008 4972 10014 4984
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 19843 5015 19901 5021
rect 19843 4981 19855 5015
rect 19889 5012 19901 5015
rect 19978 5012 19984 5024
rect 19889 4984 19984 5012
rect 19889 4981 19901 4984
rect 19843 4975 19901 4981
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 24026 4972 24032 5024
rect 24084 5012 24090 5024
rect 24719 5015 24777 5021
rect 24719 5012 24731 5015
rect 24084 4984 24731 5012
rect 24084 4972 24090 4984
rect 24719 4981 24731 4984
rect 24765 4981 24777 5015
rect 24719 4975 24777 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 6880 4780 7297 4808
rect 6880 4768 6886 4780
rect 7285 4777 7297 4780
rect 7331 4777 7343 4811
rect 7742 4808 7748 4820
rect 7703 4780 7748 4808
rect 7285 4771 7343 4777
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 8076 4780 8401 4808
rect 8076 4768 8082 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 8389 4771 8447 4777
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 10781 4811 10839 4817
rect 10781 4808 10793 4811
rect 9180 4780 10793 4808
rect 9180 4768 9186 4780
rect 10781 4777 10793 4780
rect 10827 4808 10839 4811
rect 10962 4808 10968 4820
rect 10827 4780 10968 4808
rect 10827 4777 10839 4780
rect 10781 4771 10839 4777
rect 10962 4768 10968 4780
rect 11020 4808 11026 4820
rect 11238 4808 11244 4820
rect 11020 4780 11244 4808
rect 11020 4768 11026 4780
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 13909 4811 13967 4817
rect 13909 4777 13921 4811
rect 13955 4808 13967 4811
rect 14090 4808 14096 4820
rect 13955 4780 14096 4808
rect 13955 4777 13967 4780
rect 13909 4771 13967 4777
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 18230 4808 18236 4820
rect 18191 4780 18236 4808
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 8113 4743 8171 4749
rect 8113 4709 8125 4743
rect 8159 4740 8171 4743
rect 8294 4740 8300 4752
rect 8159 4712 8300 4740
rect 8159 4709 8171 4712
rect 8113 4703 8171 4709
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 9858 4700 9864 4752
rect 9916 4740 9922 4752
rect 11419 4743 11477 4749
rect 11419 4740 11431 4743
rect 9916 4712 11431 4740
rect 9916 4700 9922 4712
rect 11419 4709 11431 4712
rect 11465 4740 11477 4743
rect 11790 4740 11796 4752
rect 11465 4712 11796 4740
rect 11465 4709 11477 4712
rect 11419 4703 11477 4709
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 15470 4700 15476 4752
rect 15528 4740 15534 4752
rect 15610 4743 15668 4749
rect 15610 4740 15622 4743
rect 15528 4712 15622 4740
rect 15528 4700 15534 4712
rect 15610 4709 15622 4712
rect 15656 4709 15668 4743
rect 17218 4740 17224 4752
rect 17179 4712 17224 4740
rect 15610 4703 15668 4709
rect 17218 4700 17224 4712
rect 17276 4700 17282 4752
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 1578 4672 1584 4684
rect 1510 4644 1584 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 1578 4632 1584 4644
rect 1636 4632 1642 4684
rect 6270 4672 6276 4684
rect 6231 4644 6276 4672
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 6730 4632 6736 4684
rect 6788 4672 6794 4684
rect 6825 4675 6883 4681
rect 6825 4672 6837 4675
rect 6788 4644 6837 4672
rect 6788 4632 6794 4644
rect 6825 4641 6837 4644
rect 6871 4641 6883 4675
rect 11054 4672 11060 4684
rect 11015 4644 11060 4672
rect 6825 4635 6883 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 13262 4672 13268 4684
rect 13223 4644 13268 4672
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 15286 4672 15292 4684
rect 15247 4644 15292 4672
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 18598 4672 18604 4684
rect 18559 4644 18604 4672
rect 18598 4632 18604 4644
rect 18656 4632 18662 4684
rect 19705 4675 19763 4681
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 19978 4672 19984 4684
rect 19751 4644 19984 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4604 6699 4607
rect 8386 4604 8392 4616
rect 6687 4576 8392 4604
rect 6687 4573 6699 4576
rect 6641 4567 6699 4573
rect 8386 4564 8392 4576
rect 8444 4604 8450 4616
rect 8757 4607 8815 4613
rect 8757 4604 8769 4607
rect 8444 4576 8769 4604
rect 8444 4564 8450 4576
rect 8757 4573 8769 4576
rect 8803 4573 8815 4607
rect 8757 4567 8815 4573
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4604 17187 4607
rect 17770 4604 17776 4616
rect 17175 4576 17776 4604
rect 17175 4573 17187 4576
rect 17129 4567 17187 4573
rect 17770 4564 17776 4576
rect 17828 4564 17834 4616
rect 1535 4539 1593 4545
rect 1535 4505 1547 4539
rect 1581 4536 1593 4539
rect 10226 4536 10232 4548
rect 1581 4508 10232 4536
rect 1581 4505 1593 4508
rect 1535 4499 1593 4505
rect 10226 4496 10232 4508
rect 10284 4496 10290 4548
rect 13449 4539 13507 4545
rect 13449 4505 13461 4539
rect 13495 4536 13507 4539
rect 14550 4536 14556 4548
rect 13495 4508 14556 4536
rect 13495 4505 13507 4508
rect 13449 4499 13507 4505
rect 14550 4496 14556 4508
rect 14608 4496 14614 4548
rect 17678 4536 17684 4548
rect 17639 4508 17684 4536
rect 17678 4496 17684 4508
rect 17736 4496 17742 4548
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 10008 4440 10149 4468
rect 10008 4428 10014 4440
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 11974 4468 11980 4480
rect 11935 4440 11980 4468
rect 10137 4431 10195 4437
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 16209 4471 16267 4477
rect 16209 4437 16221 4471
rect 16255 4468 16267 4471
rect 16482 4468 16488 4480
rect 16255 4440 16488 4468
rect 16255 4437 16267 4440
rect 16209 4431 16267 4437
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 19889 4471 19947 4477
rect 19889 4437 19901 4471
rect 19935 4468 19947 4471
rect 21358 4468 21364 4480
rect 19935 4440 21364 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 21358 4428 21364 4440
rect 21416 4428 21422 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1578 4264 1584 4276
rect 1539 4236 1584 4264
rect 1578 4224 1584 4236
rect 1636 4224 1642 4276
rect 6822 4224 6828 4276
rect 6880 4264 6886 4276
rect 7101 4267 7159 4273
rect 7101 4264 7113 4267
rect 6880 4236 7113 4264
rect 6880 4224 6886 4236
rect 7101 4233 7113 4236
rect 7147 4233 7159 4267
rect 8110 4264 8116 4276
rect 8071 4236 8116 4264
rect 7101 4227 7159 4233
rect 8110 4224 8116 4236
rect 8168 4224 8174 4276
rect 10226 4264 10232 4276
rect 10187 4236 10232 4264
rect 10226 4224 10232 4236
rect 10284 4224 10290 4276
rect 10689 4267 10747 4273
rect 10689 4233 10701 4267
rect 10735 4264 10747 4267
rect 11606 4264 11612 4276
rect 10735 4236 11612 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 3786 4156 3792 4208
rect 3844 4196 3850 4208
rect 6273 4199 6331 4205
rect 6273 4196 6285 4199
rect 3844 4168 6285 4196
rect 3844 4156 3850 4168
rect 6273 4165 6285 4168
rect 6319 4196 6331 4199
rect 6730 4196 6736 4208
rect 6319 4168 6736 4196
rect 6319 4165 6331 4168
rect 6273 4159 6331 4165
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 10134 4196 10140 4208
rect 8352 4168 10140 4196
rect 8352 4156 8358 4168
rect 10134 4156 10140 4168
rect 10192 4156 10198 4208
rect 9950 4128 9956 4140
rect 9911 4100 9956 4128
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6822 4060 6828 4072
rect 6328 4032 6828 4060
rect 6328 4020 6334 4032
rect 6822 4020 6828 4032
rect 6880 4060 6886 4072
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6880 4032 6929 4060
rect 6880 4020 6886 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4060 9183 4063
rect 9861 4063 9919 4069
rect 9861 4060 9873 4063
rect 9171 4032 9873 4060
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 9861 4029 9873 4032
rect 9907 4060 9919 4063
rect 10686 4060 10692 4072
rect 9907 4032 10692 4060
rect 9907 4029 9919 4032
rect 9861 4023 9919 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 10796 4069 10824 4236
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 18187 4267 18245 4273
rect 18187 4264 18199 4267
rect 13786 4236 18199 4264
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 13786 4196 13814 4236
rect 18187 4233 18199 4236
rect 18233 4233 18245 4267
rect 18187 4227 18245 4233
rect 18601 4267 18659 4273
rect 18601 4233 18613 4267
rect 18647 4264 18659 4267
rect 18782 4264 18788 4276
rect 18647 4236 18788 4264
rect 18647 4233 18659 4236
rect 18601 4227 18659 4233
rect 17770 4196 17776 4208
rect 10928 4168 13814 4196
rect 17731 4168 17776 4196
rect 10928 4156 10934 4168
rect 17770 4156 17776 4168
rect 17828 4156 17834 4208
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 14277 4131 14335 4137
rect 14277 4128 14289 4131
rect 11848 4100 14289 4128
rect 11848 4088 11854 4100
rect 14277 4097 14289 4100
rect 14323 4097 14335 4131
rect 14277 4091 14335 4097
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4029 10839 4063
rect 11238 4060 11244 4072
rect 11199 4032 11244 4060
rect 10781 4023 10839 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12253 4063 12311 4069
rect 12253 4060 12265 4063
rect 12032 4032 12265 4060
rect 12032 4020 12038 4032
rect 12253 4029 12265 4032
rect 12299 4060 12311 4063
rect 13081 4063 13139 4069
rect 13081 4060 13093 4063
rect 12299 4032 13093 4060
rect 12299 4029 12311 4032
rect 12253 4023 12311 4029
rect 13081 4029 13093 4032
rect 13127 4060 13139 4063
rect 13446 4060 13452 4072
rect 13127 4032 13452 4060
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 11422 3952 11428 4004
rect 11480 3992 11486 4004
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 11480 3964 11529 3992
rect 11480 3952 11486 3964
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 12434 3992 12440 4004
rect 12395 3964 12440 3992
rect 11517 3955 11575 3961
rect 12434 3952 12440 3964
rect 12492 3952 12498 4004
rect 14292 3992 14320 4091
rect 14458 4060 14464 4072
rect 14419 4032 14464 4060
rect 14458 4020 14464 4032
rect 14516 4020 14522 4072
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4060 16267 4063
rect 16482 4060 16488 4072
rect 16255 4032 16488 4060
rect 16255 4029 16267 4032
rect 16209 4023 16267 4029
rect 16482 4020 16488 4032
rect 16540 4020 16546 4072
rect 18116 4063 18174 4069
rect 18116 4029 18128 4063
rect 18162 4060 18174 4063
rect 18616 4060 18644 4227
rect 18782 4224 18788 4236
rect 18840 4224 18846 4276
rect 19797 4267 19855 4273
rect 19797 4233 19809 4267
rect 19843 4264 19855 4267
rect 19978 4264 19984 4276
rect 19843 4236 19984 4264
rect 19843 4233 19855 4236
rect 19797 4227 19855 4233
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 24854 4264 24860 4276
rect 24815 4236 24860 4264
rect 24854 4224 24860 4236
rect 24912 4224 24918 4276
rect 18162 4032 18644 4060
rect 24648 4063 24706 4069
rect 18162 4029 18174 4032
rect 18116 4023 18174 4029
rect 24648 4029 24660 4063
rect 24694 4060 24706 4063
rect 24694 4032 25176 4060
rect 24694 4029 24706 4032
rect 24648 4023 24706 4029
rect 14782 3995 14840 4001
rect 14782 3992 14794 3995
rect 14292 3964 14794 3992
rect 14782 3961 14794 3964
rect 14828 3992 14840 3995
rect 15470 3992 15476 4004
rect 14828 3964 15476 3992
rect 14828 3961 14840 3964
rect 14782 3955 14840 3961
rect 15470 3952 15476 3964
rect 15528 3992 15534 4004
rect 15657 3995 15715 4001
rect 15657 3992 15669 3995
rect 15528 3964 15669 3992
rect 15528 3952 15534 3964
rect 15657 3961 15669 3964
rect 15703 3961 15715 3995
rect 15657 3955 15715 3961
rect 17037 3995 17095 4001
rect 17037 3961 17049 3995
rect 17083 3992 17095 3995
rect 17218 3992 17224 4004
rect 17083 3964 17224 3992
rect 17083 3961 17095 3964
rect 17037 3955 17095 3961
rect 17218 3952 17224 3964
rect 17276 3992 17282 4004
rect 17313 3995 17371 4001
rect 17313 3992 17325 3995
rect 17276 3964 17325 3992
rect 17276 3952 17282 3964
rect 17313 3961 17325 3964
rect 17359 3961 17371 3995
rect 17313 3955 17371 3961
rect 566 3884 572 3936
rect 624 3924 630 3936
rect 5905 3927 5963 3933
rect 5905 3924 5917 3927
rect 624 3896 5917 3924
rect 624 3884 630 3896
rect 5905 3893 5917 3896
rect 5951 3924 5963 3927
rect 6270 3924 6276 3936
rect 5951 3896 6276 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 11790 3924 11796 3936
rect 11751 3896 11796 3924
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 13262 3924 13268 3936
rect 12216 3896 13268 3924
rect 12216 3884 12222 3896
rect 13262 3884 13268 3896
rect 13320 3924 13326 3936
rect 13449 3927 13507 3933
rect 13449 3924 13461 3927
rect 13320 3896 13461 3924
rect 13320 3884 13326 3896
rect 13449 3893 13461 3896
rect 13495 3893 13507 3927
rect 15378 3924 15384 3936
rect 15339 3896 15384 3924
rect 13449 3887 13507 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 25148 3933 25176 4032
rect 25133 3927 25191 3933
rect 25133 3893 25145 3927
rect 25179 3924 25191 3927
rect 26878 3924 26884 3936
rect 25179 3896 26884 3924
rect 25179 3893 25191 3896
rect 25133 3887 25191 3893
rect 26878 3884 26884 3896
rect 26936 3884 26942 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 6822 3720 6828 3732
rect 6783 3692 6828 3720
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 11054 3720 11060 3732
rect 11015 3692 11060 3720
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 11790 3720 11796 3732
rect 11751 3692 11796 3720
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 14458 3720 14464 3732
rect 14419 3692 14464 3720
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15749 3723 15807 3729
rect 15749 3720 15761 3723
rect 15344 3692 15761 3720
rect 15344 3680 15350 3692
rect 15749 3689 15761 3692
rect 15795 3689 15807 3723
rect 15749 3683 15807 3689
rect 13078 3612 13084 3664
rect 13136 3652 13142 3664
rect 13262 3652 13268 3664
rect 13136 3624 13268 3652
rect 13136 3612 13142 3624
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 13357 3655 13415 3661
rect 13357 3621 13369 3655
rect 13403 3652 13415 3655
rect 13446 3652 13452 3664
rect 13403 3624 13452 3652
rect 13403 3621 13415 3624
rect 13357 3615 13415 3621
rect 13446 3612 13452 3624
rect 13504 3612 13510 3664
rect 16482 3652 16488 3664
rect 16443 3624 16488 3652
rect 16482 3612 16488 3624
rect 16540 3612 16546 3664
rect 16666 3612 16672 3664
rect 16724 3652 16730 3664
rect 17037 3655 17095 3661
rect 17037 3652 17049 3655
rect 16724 3624 17049 3652
rect 16724 3612 16730 3624
rect 17037 3621 17049 3624
rect 17083 3652 17095 3655
rect 17678 3652 17684 3664
rect 17083 3624 17684 3652
rect 17083 3621 17095 3624
rect 17037 3615 17095 3621
rect 17678 3612 17684 3624
rect 17736 3612 17742 3664
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 5994 3593 6000 3596
rect 5940 3587 6000 3593
rect 5940 3584 5952 3587
rect 5316 3556 5952 3584
rect 5316 3544 5322 3556
rect 5940 3553 5952 3556
rect 5986 3553 6000 3587
rect 5940 3547 6000 3553
rect 5994 3544 6000 3547
rect 6052 3544 6058 3596
rect 18506 3584 18512 3596
rect 18467 3556 18512 3584
rect 18506 3544 18512 3556
rect 18564 3544 18570 3596
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3516 10471 3519
rect 10686 3516 10692 3528
rect 10459 3488 10692 3516
rect 10459 3485 10471 3488
rect 10413 3479 10471 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 11422 3516 11428 3528
rect 11383 3488 11428 3516
rect 11422 3476 11428 3488
rect 11480 3476 11486 3528
rect 13538 3516 13544 3528
rect 13499 3488 13544 3516
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 16390 3516 16396 3528
rect 16351 3488 16396 3516
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 17865 3519 17923 3525
rect 17865 3516 17877 3519
rect 16632 3488 17877 3516
rect 16632 3476 16638 3488
rect 17865 3485 17877 3488
rect 17911 3485 17923 3519
rect 17865 3479 17923 3485
rect 6043 3383 6101 3389
rect 6043 3349 6055 3383
rect 6089 3380 6101 3383
rect 10962 3380 10968 3392
rect 6089 3352 10968 3380
rect 6089 3349 6101 3352
rect 6043 3343 6101 3349
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 12342 3380 12348 3392
rect 12303 3352 12348 3380
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 12526 3340 12532 3392
rect 12584 3380 12590 3392
rect 12621 3383 12679 3389
rect 12621 3380 12633 3383
rect 12584 3352 12633 3380
rect 12584 3340 12590 3352
rect 12621 3349 12633 3352
rect 12667 3349 12679 3383
rect 12621 3343 12679 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 5994 3176 6000 3188
rect 5955 3148 6000 3176
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 7147 3179 7205 3185
rect 7147 3176 7159 3179
rect 6512 3148 7159 3176
rect 6512 3136 6518 3148
rect 7147 3145 7159 3148
rect 7193 3145 7205 3179
rect 7147 3139 7205 3145
rect 8895 3179 8953 3185
rect 8895 3145 8907 3179
rect 8941 3176 8953 3179
rect 9950 3176 9956 3188
rect 8941 3148 9956 3176
rect 8941 3145 8953 3148
rect 8895 3139 8953 3145
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 10045 3179 10103 3185
rect 10045 3145 10057 3179
rect 10091 3176 10103 3179
rect 12158 3176 12164 3188
rect 10091 3148 12164 3176
rect 10091 3145 10103 3148
rect 10045 3139 10103 3145
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12434 3176 12440 3188
rect 12299 3148 12440 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 16482 3176 16488 3188
rect 16443 3148 16488 3176
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 18506 3176 18512 3188
rect 18467 3148 18512 3176
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 13078 3068 13084 3120
rect 13136 3108 13142 3120
rect 14185 3111 14243 3117
rect 14185 3108 14197 3111
rect 13136 3080 14197 3108
rect 13136 3068 13142 3080
rect 14185 3077 14197 3080
rect 14231 3077 14243 3111
rect 14185 3071 14243 3077
rect 14645 3111 14703 3117
rect 14645 3077 14657 3111
rect 14691 3108 14703 3111
rect 18187 3111 18245 3117
rect 18187 3108 18199 3111
rect 14691 3080 18199 3108
rect 14691 3077 14703 3080
rect 14645 3071 14703 3077
rect 18187 3077 18199 3080
rect 18233 3077 18245 3111
rect 18187 3071 18245 3077
rect 198 3000 204 3052
rect 256 3040 262 3052
rect 13173 3043 13231 3049
rect 256 3012 8846 3040
rect 256 3000 262 3012
rect 8818 2981 8846 3012
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13538 3040 13544 3052
rect 13219 3012 13544 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 7076 2975 7134 2981
rect 7076 2941 7088 2975
rect 7122 2972 7134 2975
rect 8803 2975 8861 2981
rect 7122 2944 7604 2972
rect 7122 2941 7134 2944
rect 7076 2935 7134 2941
rect 7576 2845 7604 2944
rect 8803 2941 8815 2975
rect 8849 2972 8861 2975
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 8849 2944 9229 2972
rect 8849 2941 8861 2944
rect 8803 2935 8861 2941
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9217 2935 9275 2941
rect 9836 2975 9894 2981
rect 9836 2941 9848 2975
rect 9882 2972 9894 2975
rect 10689 2975 10747 2981
rect 9882 2944 10364 2972
rect 9882 2941 9894 2944
rect 9836 2935 9894 2941
rect 7561 2839 7619 2845
rect 7561 2805 7573 2839
rect 7607 2836 7619 2839
rect 8662 2836 8668 2848
rect 7607 2808 8668 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 10336 2845 10364 2944
rect 10689 2941 10701 2975
rect 10735 2972 10747 2975
rect 10873 2975 10931 2981
rect 10873 2972 10885 2975
rect 10735 2944 10885 2972
rect 10735 2941 10747 2944
rect 10689 2935 10747 2941
rect 10873 2941 10885 2944
rect 10919 2972 10931 2975
rect 12342 2972 12348 2984
rect 10919 2944 12348 2972
rect 10919 2941 10931 2944
rect 10873 2935 10931 2941
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 13262 2932 13268 2984
rect 13320 2972 13326 2984
rect 13817 2975 13875 2981
rect 13817 2972 13829 2975
rect 13320 2944 13829 2972
rect 13320 2932 13326 2944
rect 13817 2941 13829 2944
rect 13863 2941 13875 2975
rect 13817 2935 13875 2941
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2972 14059 2975
rect 14660 2972 14688 3071
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 15059 3012 15577 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 15565 3009 15577 3012
rect 15611 3040 15623 3043
rect 16666 3040 16672 3052
rect 15611 3012 16672 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 17586 3000 17592 3052
rect 17644 3040 17650 3052
rect 17644 3012 19334 3040
rect 17644 3000 17650 3012
rect 14047 2944 14688 2972
rect 14047 2941 14059 2944
rect 14001 2935 14059 2941
rect 16206 2932 16212 2984
rect 16264 2972 16270 2984
rect 19076 2981 19104 3012
rect 18116 2975 18174 2981
rect 18116 2972 18128 2975
rect 16264 2944 18128 2972
rect 16264 2932 16270 2944
rect 18116 2941 18128 2944
rect 18162 2972 18174 2975
rect 18877 2975 18935 2981
rect 18877 2972 18889 2975
rect 18162 2944 18889 2972
rect 18162 2941 18174 2944
rect 18116 2935 18174 2941
rect 18877 2941 18889 2944
rect 18923 2941 18935 2975
rect 19076 2975 19154 2981
rect 19076 2944 19108 2975
rect 18877 2935 18935 2941
rect 19096 2941 19108 2944
rect 19142 2941 19154 2975
rect 19306 2972 19334 3012
rect 19521 2975 19579 2981
rect 19521 2972 19533 2975
rect 19306 2944 19533 2972
rect 19096 2935 19154 2941
rect 19521 2941 19533 2944
rect 19567 2941 19579 2975
rect 19521 2935 19579 2941
rect 10778 2904 10784 2916
rect 10739 2876 10784 2904
rect 10778 2864 10784 2876
rect 10836 2864 10842 2916
rect 12526 2904 12532 2916
rect 12487 2876 12532 2904
rect 12526 2864 12532 2876
rect 12584 2864 12590 2916
rect 12621 2907 12679 2913
rect 12621 2873 12633 2907
rect 12667 2873 12679 2907
rect 12621 2867 12679 2873
rect 15657 2907 15715 2913
rect 15657 2873 15669 2907
rect 15703 2904 15715 2907
rect 18506 2904 18512 2916
rect 15703 2876 18512 2904
rect 15703 2873 15715 2876
rect 15657 2867 15715 2873
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 11606 2836 11612 2848
rect 10367 2808 11612 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 11790 2836 11796 2848
rect 11751 2808 11796 2836
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12636 2836 12664 2867
rect 15378 2836 15384 2848
rect 12492 2808 12664 2836
rect 15291 2808 15384 2836
rect 12492 2796 12498 2808
rect 15378 2796 15384 2808
rect 15436 2836 15442 2848
rect 15672 2836 15700 2867
rect 18506 2864 18512 2876
rect 18564 2864 18570 2916
rect 15436 2808 15700 2836
rect 15436 2796 15442 2808
rect 16390 2796 16396 2848
rect 16448 2836 16454 2848
rect 16945 2839 17003 2845
rect 16945 2836 16957 2839
rect 16448 2808 16957 2836
rect 16448 2796 16454 2808
rect 16945 2805 16957 2808
rect 16991 2836 17003 2839
rect 17494 2836 17500 2848
rect 16991 2808 17500 2836
rect 16991 2805 17003 2808
rect 16945 2799 17003 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 17586 2796 17592 2848
rect 17644 2836 17650 2848
rect 19199 2839 19257 2845
rect 19199 2836 19211 2839
rect 17644 2808 19211 2836
rect 17644 2796 17650 2808
rect 19199 2805 19211 2808
rect 19245 2805 19257 2839
rect 19199 2799 19257 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7193 2635 7251 2641
rect 7193 2632 7205 2635
rect 7156 2604 7205 2632
rect 7156 2592 7162 2604
rect 7193 2601 7205 2604
rect 7239 2601 7251 2635
rect 7193 2595 7251 2601
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 8803 2635 8861 2641
rect 8803 2632 8815 2635
rect 7524 2604 8815 2632
rect 7524 2592 7530 2604
rect 8803 2601 8815 2604
rect 8849 2601 8861 2635
rect 10778 2632 10784 2644
rect 10739 2604 10784 2632
rect 8803 2595 8861 2601
rect 10778 2592 10784 2604
rect 10836 2632 10842 2644
rect 10836 2604 11192 2632
rect 10836 2592 10842 2604
rect 10505 2567 10563 2573
rect 10505 2533 10517 2567
rect 10551 2564 10563 2567
rect 10686 2564 10692 2576
rect 10551 2536 10692 2564
rect 10551 2533 10563 2536
rect 10505 2527 10563 2533
rect 10686 2524 10692 2536
rect 10744 2564 10750 2576
rect 11164 2573 11192 2604
rect 11422 2592 11428 2644
rect 11480 2632 11486 2644
rect 11977 2635 12035 2641
rect 11977 2632 11989 2635
rect 11480 2604 11989 2632
rect 11480 2592 11486 2604
rect 11977 2601 11989 2604
rect 12023 2601 12035 2635
rect 12342 2632 12348 2644
rect 12303 2604 12348 2632
rect 11977 2595 12035 2601
rect 12342 2592 12348 2604
rect 12400 2632 12406 2644
rect 12618 2632 12624 2644
rect 12400 2604 12624 2632
rect 12400 2592 12406 2604
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 12768 2604 12848 2632
rect 12768 2592 12774 2604
rect 12820 2573 12848 2604
rect 12894 2592 12900 2644
rect 12952 2632 12958 2644
rect 13538 2632 13544 2644
rect 12952 2604 13544 2632
rect 12952 2592 12958 2604
rect 13538 2592 13544 2604
rect 13596 2632 13602 2644
rect 13633 2635 13691 2641
rect 13633 2632 13645 2635
rect 13596 2604 13645 2632
rect 13596 2592 13602 2604
rect 13633 2601 13645 2604
rect 13679 2601 13691 2635
rect 13633 2595 13691 2601
rect 15197 2635 15255 2641
rect 15197 2601 15209 2635
rect 15243 2632 15255 2635
rect 16574 2632 16580 2644
rect 15243 2604 16580 2632
rect 15243 2601 15255 2604
rect 15197 2595 15255 2601
rect 11057 2567 11115 2573
rect 11057 2564 11069 2567
rect 10744 2536 11069 2564
rect 10744 2524 10750 2536
rect 11057 2533 11069 2536
rect 11103 2533 11115 2567
rect 11057 2527 11115 2533
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2533 11207 2567
rect 11149 2527 11207 2533
rect 12805 2567 12863 2573
rect 12805 2533 12817 2567
rect 12851 2533 12863 2567
rect 12805 2527 12863 2533
rect 14921 2567 14979 2573
rect 14921 2533 14933 2567
rect 14967 2564 14979 2567
rect 15286 2564 15292 2576
rect 14967 2536 15292 2564
rect 14967 2533 14979 2536
rect 14921 2527 14979 2533
rect 15286 2524 15292 2536
rect 15344 2564 15350 2576
rect 15672 2573 15700 2604
rect 16574 2592 16580 2604
rect 16632 2592 16638 2644
rect 16942 2592 16948 2644
rect 17000 2632 17006 2644
rect 17359 2635 17417 2641
rect 17359 2632 17371 2635
rect 17000 2604 17371 2632
rect 17000 2592 17006 2604
rect 17359 2601 17371 2604
rect 17405 2601 17417 2635
rect 17359 2595 17417 2601
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 19567 2635 19625 2641
rect 19567 2632 19579 2635
rect 17552 2604 19579 2632
rect 17552 2592 17558 2604
rect 19567 2601 19579 2604
rect 19613 2601 19625 2635
rect 19567 2595 19625 2601
rect 15565 2567 15623 2573
rect 15565 2564 15577 2567
rect 15344 2536 15577 2564
rect 15344 2524 15350 2536
rect 15565 2533 15577 2536
rect 15611 2533 15623 2567
rect 15565 2527 15623 2533
rect 15657 2567 15715 2573
rect 15657 2533 15669 2567
rect 15703 2533 15715 2567
rect 16206 2564 16212 2576
rect 16167 2536 16212 2564
rect 15657 2527 15715 2533
rect 16206 2524 16212 2536
rect 16264 2524 16270 2576
rect 17770 2524 17776 2576
rect 17828 2564 17834 2576
rect 17828 2536 19539 2564
rect 17828 2524 17834 2536
rect 6984 2499 7042 2505
rect 6984 2465 6996 2499
rect 7030 2496 7042 2499
rect 7466 2496 7472 2508
rect 7030 2468 7472 2496
rect 7030 2465 7042 2468
rect 6984 2459 7042 2465
rect 7466 2456 7472 2468
rect 7524 2456 7530 2508
rect 8732 2499 8790 2505
rect 8732 2465 8744 2499
rect 8778 2496 8790 2499
rect 9585 2499 9643 2505
rect 8778 2468 9260 2496
rect 8778 2465 8790 2468
rect 8732 2459 8790 2465
rect 9232 2437 9260 2468
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 9861 2499 9919 2505
rect 9861 2496 9873 2499
rect 9631 2468 9873 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 9861 2465 9873 2468
rect 9907 2496 9919 2499
rect 10870 2496 10876 2508
rect 9907 2468 10876 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 17288 2499 17346 2505
rect 17288 2465 17300 2499
rect 17334 2496 17346 2499
rect 18322 2496 18328 2508
rect 17334 2468 17816 2496
rect 18283 2468 18328 2496
rect 17334 2465 17346 2468
rect 17288 2459 17346 2465
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 10134 2428 10140 2440
rect 9263 2400 10140 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 12710 2388 12716 2440
rect 12768 2428 12774 2440
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12768 2400 12813 2428
rect 12912 2400 13001 2428
rect 12768 2388 12774 2400
rect 10045 2363 10103 2369
rect 10045 2329 10057 2363
rect 10091 2360 10103 2363
rect 11514 2360 11520 2372
rect 10091 2332 11520 2360
rect 10091 2329 10103 2332
rect 10045 2323 10103 2329
rect 11514 2320 11520 2332
rect 11572 2320 11578 2372
rect 11606 2320 11612 2372
rect 11664 2360 11670 2372
rect 12912 2360 12940 2400
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 14185 2431 14243 2437
rect 14185 2397 14197 2431
rect 14231 2428 14243 2431
rect 14292 2428 14320 2459
rect 17586 2428 17592 2440
rect 14231 2400 17592 2428
rect 14231 2397 14243 2400
rect 14185 2391 14243 2397
rect 17586 2388 17592 2400
rect 17644 2388 17650 2440
rect 11664 2332 12940 2360
rect 14461 2363 14519 2369
rect 11664 2320 11670 2332
rect 14461 2329 14473 2363
rect 14507 2360 14519 2363
rect 15654 2360 15660 2372
rect 14507 2332 15660 2360
rect 14507 2329 14519 2332
rect 14461 2323 14519 2329
rect 15654 2320 15660 2332
rect 15712 2320 15718 2372
rect 7466 2292 7472 2304
rect 7427 2264 7472 2292
rect 7466 2252 7472 2264
rect 7524 2252 7530 2304
rect 17788 2301 17816 2468
rect 18322 2456 18328 2468
rect 18380 2496 18386 2508
rect 19511 2505 19539 2536
rect 18877 2499 18935 2505
rect 18877 2496 18889 2499
rect 18380 2468 18889 2496
rect 18380 2456 18386 2468
rect 18877 2465 18889 2468
rect 18923 2465 18935 2499
rect 18877 2459 18935 2465
rect 19496 2499 19554 2505
rect 19496 2465 19508 2499
rect 19542 2496 19554 2499
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19542 2468 19901 2496
rect 19542 2465 19554 2468
rect 19496 2459 19554 2465
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 21244 2499 21302 2505
rect 21244 2465 21256 2499
rect 21290 2496 21302 2499
rect 21290 2468 21772 2496
rect 21290 2465 21302 2468
rect 21244 2459 21302 2465
rect 18509 2363 18567 2369
rect 18509 2329 18521 2363
rect 18555 2360 18567 2363
rect 19978 2360 19984 2372
rect 18555 2332 19984 2360
rect 18555 2329 18567 2332
rect 18509 2323 18567 2329
rect 19978 2320 19984 2332
rect 20036 2320 20042 2372
rect 17773 2295 17831 2301
rect 17773 2261 17785 2295
rect 17819 2292 17831 2295
rect 18414 2292 18420 2304
rect 17819 2264 18420 2292
rect 17819 2261 17831 2264
rect 17773 2255 17831 2261
rect 18414 2252 18420 2264
rect 18472 2252 18478 2304
rect 19702 2252 19708 2304
rect 19760 2292 19766 2304
rect 21744 2301 21772 2468
rect 21315 2295 21373 2301
rect 21315 2292 21327 2295
rect 19760 2264 21327 2292
rect 19760 2252 19766 2264
rect 21315 2261 21327 2264
rect 21361 2261 21373 2295
rect 21315 2255 21373 2261
rect 21729 2295 21787 2301
rect 21729 2261 21741 2295
rect 21775 2292 21787 2295
rect 22646 2292 22652 2304
rect 21775 2264 22652 2292
rect 21775 2261 21787 2264
rect 21729 2255 21787 2261
rect 22646 2252 22652 2264
rect 22704 2252 22710 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 23756 27480 23808 27532
rect 25136 27480 25188 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 6276 24216 6328 24268
rect 7564 24216 7616 24268
rect 8300 24216 8352 24268
rect 10140 24216 10192 24268
rect 6368 24012 6420 24064
rect 6828 24012 6880 24064
rect 8668 24012 8720 24064
rect 10048 24012 10100 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2780 23851 2832 23860
rect 2780 23817 2789 23851
rect 2789 23817 2823 23851
rect 2823 23817 2832 23851
rect 2780 23808 2832 23817
rect 6276 23808 6328 23860
rect 6460 23808 6512 23860
rect 8300 23851 8352 23860
rect 8300 23817 8309 23851
rect 8309 23817 8343 23851
rect 8343 23817 8352 23851
rect 8300 23808 8352 23817
rect 10140 23808 10192 23860
rect 15844 23808 15896 23860
rect 940 23740 992 23792
rect 2780 23604 2832 23656
rect 8668 23672 8720 23724
rect 6828 23647 6880 23656
rect 6828 23613 6837 23647
rect 6837 23613 6871 23647
rect 6871 23613 6880 23647
rect 6828 23604 6880 23613
rect 9128 23579 9180 23588
rect 2504 23468 2556 23520
rect 4528 23468 4580 23520
rect 9128 23545 9137 23579
rect 9137 23545 9171 23579
rect 9171 23545 9180 23579
rect 9128 23536 9180 23545
rect 8852 23468 8904 23520
rect 12808 23604 12860 23656
rect 18604 23604 18656 23656
rect 21364 23808 21416 23860
rect 23296 23808 23348 23860
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 25136 23604 25188 23656
rect 9956 23579 10008 23588
rect 9956 23545 9965 23579
rect 9965 23545 9999 23579
rect 9999 23545 10008 23579
rect 9956 23536 10008 23545
rect 21732 23536 21784 23588
rect 17776 23468 17828 23520
rect 18604 23511 18656 23520
rect 18604 23477 18613 23511
rect 18613 23477 18647 23511
rect 18647 23477 18656 23511
rect 18604 23468 18656 23477
rect 18696 23468 18748 23520
rect 19984 23468 20036 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 6828 23307 6880 23316
rect 6828 23273 6837 23307
rect 6837 23273 6871 23307
rect 6871 23273 6880 23307
rect 6828 23264 6880 23273
rect 5540 23239 5592 23248
rect 5540 23205 5549 23239
rect 5549 23205 5583 23239
rect 5583 23205 5592 23239
rect 5540 23196 5592 23205
rect 8116 23196 8168 23248
rect 9772 23196 9824 23248
rect 9956 23196 10008 23248
rect 1216 23128 1268 23180
rect 24676 23128 24728 23180
rect 4528 23060 4580 23112
rect 5448 23103 5500 23112
rect 5448 23069 5457 23103
rect 5457 23069 5491 23103
rect 5491 23069 5500 23103
rect 5448 23060 5500 23069
rect 6276 23060 6328 23112
rect 7840 23060 7892 23112
rect 8760 23103 8812 23112
rect 8760 23069 8769 23103
rect 8769 23069 8803 23103
rect 8803 23069 8812 23103
rect 8760 23060 8812 23069
rect 10140 23060 10192 23112
rect 18696 23060 18748 23112
rect 7564 23035 7616 23044
rect 7564 23001 7573 23035
rect 7573 23001 7607 23035
rect 7607 23001 7616 23035
rect 9128 23035 9180 23044
rect 7564 22992 7616 23001
rect 9128 23001 9137 23035
rect 9137 23001 9171 23035
rect 9171 23001 9180 23035
rect 9128 22992 9180 23001
rect 2320 22924 2372 22976
rect 22192 22924 22244 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1216 22720 1268 22772
rect 9772 22763 9824 22772
rect 9772 22729 9781 22763
rect 9781 22729 9815 22763
rect 9815 22729 9824 22763
rect 9772 22720 9824 22729
rect 10140 22763 10192 22772
rect 10140 22729 10149 22763
rect 10149 22729 10183 22763
rect 10183 22729 10192 22763
rect 10140 22720 10192 22729
rect 17684 22720 17736 22772
rect 24676 22763 24728 22772
rect 24676 22729 24685 22763
rect 24685 22729 24719 22763
rect 24719 22729 24728 22763
rect 24676 22720 24728 22729
rect 5540 22584 5592 22636
rect 6276 22584 6328 22636
rect 9128 22652 9180 22704
rect 8760 22584 8812 22636
rect 11244 22516 11296 22568
rect 6920 22491 6972 22500
rect 6920 22457 6929 22491
rect 6929 22457 6963 22491
rect 6963 22457 6972 22491
rect 6920 22448 6972 22457
rect 6552 22423 6604 22432
rect 6552 22389 6561 22423
rect 6561 22389 6595 22423
rect 6595 22389 6604 22423
rect 8944 22448 8996 22500
rect 8024 22423 8076 22432
rect 6552 22380 6604 22389
rect 8024 22389 8033 22423
rect 8033 22389 8067 22423
rect 8067 22389 8076 22423
rect 8024 22380 8076 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5448 22219 5500 22228
rect 5448 22185 5457 22219
rect 5457 22185 5491 22219
rect 5491 22185 5500 22219
rect 5448 22176 5500 22185
rect 6920 22219 6972 22228
rect 6920 22185 6929 22219
rect 6929 22185 6963 22219
rect 6963 22185 6972 22219
rect 6920 22176 6972 22185
rect 7840 22219 7892 22228
rect 7840 22185 7849 22219
rect 7849 22185 7883 22219
rect 7883 22185 7892 22219
rect 7840 22176 7892 22185
rect 8024 22151 8076 22160
rect 8024 22117 8033 22151
rect 8033 22117 8067 22151
rect 8067 22117 8076 22151
rect 8024 22108 8076 22117
rect 8944 22040 8996 22092
rect 11428 22040 11480 22092
rect 12072 22040 12124 22092
rect 13544 22040 13596 22092
rect 8944 21836 8996 21888
rect 11888 21836 11940 21888
rect 12532 21879 12584 21888
rect 12532 21845 12541 21879
rect 12541 21845 12575 21879
rect 12575 21845 12584 21879
rect 12532 21836 12584 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 11244 21632 11296 21684
rect 11428 21675 11480 21684
rect 11428 21641 11437 21675
rect 11437 21641 11471 21675
rect 11471 21641 11480 21675
rect 11428 21632 11480 21641
rect 13544 21675 13596 21684
rect 13544 21641 13553 21675
rect 13553 21641 13587 21675
rect 13587 21641 13596 21675
rect 13544 21632 13596 21641
rect 12440 21564 12492 21616
rect 12532 21539 12584 21548
rect 12532 21505 12541 21539
rect 12541 21505 12575 21539
rect 12575 21505 12584 21539
rect 12532 21496 12584 21505
rect 10784 21428 10836 21480
rect 12624 21403 12676 21412
rect 12624 21369 12633 21403
rect 12633 21369 12667 21403
rect 12667 21369 12676 21403
rect 12624 21360 12676 21369
rect 8944 21292 8996 21344
rect 9680 21335 9732 21344
rect 9680 21301 9689 21335
rect 9689 21301 9723 21335
rect 9723 21301 9732 21335
rect 9680 21292 9732 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 11888 21063 11940 21072
rect 11888 21029 11897 21063
rect 11897 21029 11931 21063
rect 11931 21029 11940 21063
rect 11888 21020 11940 21029
rect 12164 21020 12216 21072
rect 7288 20995 7340 21004
rect 7288 20961 7297 20995
rect 7297 20961 7331 20995
rect 7331 20961 7340 20995
rect 7288 20952 7340 20961
rect 10324 20995 10376 21004
rect 10324 20961 10333 20995
rect 10333 20961 10367 20995
rect 10367 20961 10376 20995
rect 10324 20952 10376 20961
rect 12440 20859 12492 20868
rect 12440 20825 12449 20859
rect 12449 20825 12483 20859
rect 12483 20825 12492 20859
rect 12440 20816 12492 20825
rect 8576 20748 8628 20800
rect 9956 20791 10008 20800
rect 9956 20757 9965 20791
rect 9965 20757 9999 20791
rect 9999 20757 10008 20791
rect 9956 20748 10008 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 7288 20587 7340 20596
rect 7288 20553 7297 20587
rect 7297 20553 7331 20587
rect 7331 20553 7340 20587
rect 7288 20544 7340 20553
rect 9680 20544 9732 20596
rect 9956 20587 10008 20596
rect 9956 20553 9965 20587
rect 9965 20553 9999 20587
rect 9999 20553 10008 20587
rect 9956 20544 10008 20553
rect 10324 20544 10376 20596
rect 11888 20544 11940 20596
rect 12624 20544 12676 20596
rect 8576 20451 8628 20460
rect 8576 20417 8585 20451
rect 8585 20417 8619 20451
rect 8619 20417 8628 20451
rect 8576 20408 8628 20417
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 8668 20315 8720 20324
rect 8668 20281 8677 20315
rect 8677 20281 8711 20315
rect 8711 20281 8720 20315
rect 8668 20272 8720 20281
rect 9220 20315 9272 20324
rect 9220 20281 9229 20315
rect 9229 20281 9263 20315
rect 9263 20281 9272 20315
rect 9220 20272 9272 20281
rect 9956 20204 10008 20256
rect 12164 20247 12216 20256
rect 12164 20213 12173 20247
rect 12173 20213 12207 20247
rect 12207 20213 12216 20247
rect 12164 20204 12216 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 4804 19839 4856 19848
rect 4804 19805 4813 19839
rect 4813 19805 4847 19839
rect 4847 19805 4856 19839
rect 4804 19796 4856 19805
rect 6276 20000 6328 20052
rect 6000 19975 6052 19984
rect 6000 19941 6009 19975
rect 6009 19941 6043 19975
rect 6043 19941 6052 19975
rect 6000 19932 6052 19941
rect 8116 19932 8168 19984
rect 10140 19932 10192 19984
rect 10784 19932 10836 19984
rect 13912 20000 13964 20052
rect 11336 19907 11388 19916
rect 11336 19873 11345 19907
rect 11345 19873 11379 19907
rect 11379 19873 11388 19907
rect 11336 19864 11388 19873
rect 12900 19907 12952 19916
rect 12900 19873 12909 19907
rect 12909 19873 12943 19907
rect 12943 19873 12952 19907
rect 12900 19864 12952 19873
rect 5448 19728 5500 19780
rect 7472 19660 7524 19712
rect 9220 19796 9272 19848
rect 10232 19796 10284 19848
rect 8668 19728 8720 19780
rect 11336 19728 11388 19780
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 6000 19456 6052 19508
rect 6460 19456 6512 19508
rect 8116 19499 8168 19508
rect 8116 19465 8125 19499
rect 8125 19465 8159 19499
rect 8159 19465 8168 19499
rect 8116 19456 8168 19465
rect 10140 19456 10192 19508
rect 10232 19456 10284 19508
rect 11336 19499 11388 19508
rect 11336 19465 11345 19499
rect 11345 19465 11379 19499
rect 11379 19465 11388 19499
rect 11336 19456 11388 19465
rect 14648 19499 14700 19508
rect 14648 19465 14657 19499
rect 14657 19465 14691 19499
rect 14691 19465 14700 19499
rect 14648 19456 14700 19465
rect 12900 19388 12952 19440
rect 3976 19320 4028 19372
rect 4804 19320 4856 19372
rect 5448 19320 5500 19372
rect 6460 19252 6512 19304
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 8576 19159 8628 19168
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 14648 19252 14700 19304
rect 13176 19116 13228 19168
rect 14096 19116 14148 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2504 18912 2556 18964
rect 3240 18912 3292 18964
rect 4252 18955 4304 18964
rect 4252 18921 4261 18955
rect 4261 18921 4295 18955
rect 4295 18921 4304 18955
rect 4252 18912 4304 18921
rect 6460 18955 6512 18964
rect 6460 18921 6469 18955
rect 6469 18921 6503 18955
rect 6503 18921 6512 18955
rect 6460 18912 6512 18921
rect 8024 18955 8076 18964
rect 8024 18921 8033 18955
rect 8033 18921 8067 18955
rect 8067 18921 8076 18955
rect 8024 18912 8076 18921
rect 12164 18955 12216 18964
rect 12164 18921 12173 18955
rect 12173 18921 12207 18955
rect 12207 18921 12216 18955
rect 12164 18912 12216 18921
rect 3976 18844 4028 18896
rect 6092 18844 6144 18896
rect 11704 18844 11756 18896
rect 1952 18776 2004 18828
rect 2504 18776 2556 18828
rect 4252 18776 4304 18828
rect 7564 18776 7616 18828
rect 8208 18819 8260 18828
rect 8208 18785 8217 18819
rect 8217 18785 8251 18819
rect 8251 18785 8260 18819
rect 8208 18776 8260 18785
rect 5540 18751 5592 18760
rect 5540 18717 5549 18751
rect 5549 18717 5583 18751
rect 5583 18717 5592 18751
rect 5540 18708 5592 18717
rect 10784 18708 10836 18760
rect 12992 18751 13044 18760
rect 12992 18717 13001 18751
rect 13001 18717 13035 18751
rect 13035 18717 13044 18751
rect 12992 18708 13044 18717
rect 2228 18640 2280 18692
rect 1676 18572 1728 18624
rect 8760 18615 8812 18624
rect 8760 18581 8769 18615
rect 8769 18581 8803 18615
rect 8803 18581 8812 18615
rect 8760 18572 8812 18581
rect 11428 18572 11480 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 2504 18411 2556 18420
rect 2504 18377 2513 18411
rect 2513 18377 2547 18411
rect 2547 18377 2556 18411
rect 2504 18368 2556 18377
rect 5448 18368 5500 18420
rect 8668 18368 8720 18420
rect 19524 18368 19576 18420
rect 4252 18343 4304 18352
rect 4252 18309 4261 18343
rect 4261 18309 4295 18343
rect 4295 18309 4304 18343
rect 4252 18300 4304 18309
rect 12624 18300 12676 18352
rect 3240 18275 3292 18284
rect 3240 18241 3249 18275
rect 3249 18241 3283 18275
rect 3283 18241 3292 18275
rect 3240 18232 3292 18241
rect 5540 18232 5592 18284
rect 8024 18275 8076 18284
rect 8024 18241 8033 18275
rect 8033 18241 8067 18275
rect 8067 18241 8076 18275
rect 8024 18232 8076 18241
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 12532 18232 12584 18241
rect 12992 18232 13044 18284
rect 1676 18164 1728 18216
rect 5172 18207 5224 18216
rect 5172 18173 5181 18207
rect 5181 18173 5215 18207
rect 5215 18173 5224 18207
rect 5172 18164 5224 18173
rect 6184 18164 6236 18216
rect 11428 18207 11480 18216
rect 11428 18173 11437 18207
rect 11437 18173 11471 18207
rect 11471 18173 11480 18207
rect 11428 18164 11480 18173
rect 18328 18164 18380 18216
rect 23756 18207 23808 18216
rect 23756 18173 23774 18207
rect 23774 18173 23808 18207
rect 23756 18164 23808 18173
rect 3332 18139 3384 18148
rect 3332 18105 3341 18139
rect 3341 18105 3375 18139
rect 3375 18105 3384 18139
rect 3332 18096 3384 18105
rect 3884 18139 3936 18148
rect 3884 18105 3893 18139
rect 3893 18105 3927 18139
rect 3927 18105 3936 18139
rect 3884 18096 3936 18105
rect 112 18028 164 18080
rect 6092 18028 6144 18080
rect 7564 18071 7616 18080
rect 7564 18037 7573 18071
rect 7573 18037 7607 18071
rect 7607 18037 7616 18071
rect 7564 18028 7616 18037
rect 7748 18028 7800 18080
rect 8576 18096 8628 18148
rect 13176 18139 13228 18148
rect 10784 18028 10836 18080
rect 11704 18028 11756 18080
rect 13176 18105 13185 18139
rect 13185 18105 13219 18139
rect 13219 18105 13228 18139
rect 13176 18096 13228 18105
rect 17500 18028 17552 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1676 17867 1728 17876
rect 1676 17833 1685 17867
rect 1685 17833 1719 17867
rect 1719 17833 1728 17867
rect 1676 17824 1728 17833
rect 6552 17867 6604 17876
rect 6552 17833 6561 17867
rect 6561 17833 6595 17867
rect 6595 17833 6604 17867
rect 6552 17824 6604 17833
rect 11428 17824 11480 17876
rect 12532 17867 12584 17876
rect 2228 17756 2280 17808
rect 2596 17799 2648 17808
rect 2596 17765 2605 17799
rect 2605 17765 2639 17799
rect 2639 17765 2648 17799
rect 2596 17756 2648 17765
rect 3332 17756 3384 17808
rect 5540 17756 5592 17808
rect 6092 17756 6144 17808
rect 8760 17799 8812 17808
rect 8760 17765 8769 17799
rect 8769 17765 8803 17799
rect 8803 17765 8812 17799
rect 8760 17756 8812 17765
rect 10508 17756 10560 17808
rect 11704 17756 11756 17808
rect 12532 17833 12541 17867
rect 12541 17833 12575 17867
rect 12575 17833 12584 17867
rect 12532 17824 12584 17833
rect 12624 17824 12676 17876
rect 18328 17867 18380 17876
rect 18328 17833 18337 17867
rect 18337 17833 18371 17867
rect 18371 17833 18380 17867
rect 18328 17824 18380 17833
rect 13452 17756 13504 17808
rect 4620 17731 4672 17740
rect 4620 17697 4629 17731
rect 4629 17697 4663 17731
rect 4663 17697 4672 17731
rect 4620 17688 4672 17697
rect 8024 17731 8076 17740
rect 8024 17697 8033 17731
rect 8033 17697 8067 17731
rect 8067 17697 8076 17731
rect 8024 17688 8076 17697
rect 3884 17620 3936 17672
rect 6000 17620 6052 17672
rect 6184 17484 6236 17536
rect 6828 17484 6880 17536
rect 8208 17620 8260 17672
rect 14372 17688 14424 17740
rect 18420 17688 18472 17740
rect 24676 17688 24728 17740
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 12900 17620 12952 17672
rect 13176 17663 13228 17672
rect 13176 17629 13185 17663
rect 13185 17629 13219 17663
rect 13219 17629 13228 17663
rect 13176 17620 13228 17629
rect 10508 17484 10560 17536
rect 22284 17484 22336 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2228 17280 2280 17332
rect 4620 17323 4672 17332
rect 4620 17289 4629 17323
rect 4629 17289 4663 17323
rect 4663 17289 4672 17323
rect 4620 17280 4672 17289
rect 6000 17323 6052 17332
rect 6000 17289 6009 17323
rect 6009 17289 6043 17323
rect 6043 17289 6052 17323
rect 6000 17280 6052 17289
rect 8944 17323 8996 17332
rect 8944 17289 8953 17323
rect 8953 17289 8987 17323
rect 8987 17289 8996 17323
rect 8944 17280 8996 17289
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 24676 17323 24728 17332
rect 24676 17289 24685 17323
rect 24685 17289 24719 17323
rect 24719 17289 24728 17323
rect 24676 17280 24728 17289
rect 2596 17212 2648 17264
rect 5172 17212 5224 17264
rect 6644 17212 6696 17264
rect 8024 17212 8076 17264
rect 11428 17212 11480 17264
rect 3700 17119 3752 17128
rect 3700 17085 3709 17119
rect 3709 17085 3743 17119
rect 3743 17085 3752 17119
rect 3700 17076 3752 17085
rect 8208 17076 8260 17128
rect 4620 17008 4672 17060
rect 5540 17008 5592 17060
rect 7748 17008 7800 17060
rect 10508 17144 10560 17196
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 18052 17051 18104 17060
rect 6828 16940 6880 16992
rect 10140 16983 10192 16992
rect 10140 16949 10149 16983
rect 10149 16949 10183 16983
rect 10183 16949 10192 16983
rect 10140 16940 10192 16949
rect 18052 17017 18061 17051
rect 18061 17017 18095 17051
rect 18095 17017 18104 17051
rect 18052 17008 18104 17017
rect 14372 16940 14424 16992
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 18236 16940 18288 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 3884 16736 3936 16788
rect 4804 16736 4856 16788
rect 6000 16736 6052 16788
rect 8852 16736 8904 16788
rect 12532 16779 12584 16788
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 7748 16668 7800 16720
rect 10876 16711 10928 16720
rect 10876 16677 10885 16711
rect 10885 16677 10919 16711
rect 10919 16677 10928 16711
rect 10876 16668 10928 16677
rect 11428 16711 11480 16720
rect 11428 16677 11437 16711
rect 11437 16677 11471 16711
rect 11471 16677 11480 16711
rect 11428 16668 11480 16677
rect 13912 16668 13964 16720
rect 14372 16711 14424 16720
rect 14372 16677 14381 16711
rect 14381 16677 14415 16711
rect 14415 16677 14424 16711
rect 14372 16668 14424 16677
rect 17592 16668 17644 16720
rect 18052 16668 18104 16720
rect 5540 16643 5592 16652
rect 5540 16609 5549 16643
rect 5549 16609 5583 16643
rect 5583 16609 5592 16643
rect 5540 16600 5592 16609
rect 6184 16600 6236 16652
rect 9404 16600 9456 16652
rect 10232 16643 10284 16652
rect 10232 16609 10241 16643
rect 10241 16609 10275 16643
rect 10275 16609 10284 16643
rect 10232 16600 10284 16609
rect 12900 16600 12952 16652
rect 3516 16396 3568 16448
rect 3700 16439 3752 16448
rect 3700 16405 3709 16439
rect 3709 16405 3743 16439
rect 3743 16405 3752 16439
rect 3700 16396 3752 16405
rect 11428 16532 11480 16584
rect 13728 16575 13780 16584
rect 13728 16541 13737 16575
rect 13737 16541 13771 16575
rect 13771 16541 13780 16575
rect 13728 16532 13780 16541
rect 17224 16532 17276 16584
rect 17500 16464 17552 16516
rect 18420 16464 18472 16516
rect 7932 16396 7984 16448
rect 14740 16439 14792 16448
rect 14740 16405 14749 16439
rect 14749 16405 14783 16439
rect 14783 16405 14792 16439
rect 14740 16396 14792 16405
rect 18236 16396 18288 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 5172 16192 5224 16244
rect 7748 16235 7800 16244
rect 7748 16201 7757 16235
rect 7757 16201 7791 16235
rect 7791 16201 7800 16235
rect 7748 16192 7800 16201
rect 11336 16235 11388 16244
rect 11336 16201 11345 16235
rect 11345 16201 11379 16235
rect 11379 16201 11388 16235
rect 11336 16192 11388 16201
rect 13728 16192 13780 16244
rect 17224 16235 17276 16244
rect 17224 16201 17233 16235
rect 17233 16201 17267 16235
rect 17267 16201 17276 16235
rect 17224 16192 17276 16201
rect 17592 16235 17644 16244
rect 17592 16201 17601 16235
rect 17601 16201 17635 16235
rect 17635 16201 17644 16235
rect 17592 16192 17644 16201
rect 25136 16235 25188 16244
rect 25136 16201 25145 16235
rect 25145 16201 25179 16235
rect 25179 16201 25188 16235
rect 25136 16192 25188 16201
rect 3700 16099 3752 16108
rect 3700 16065 3709 16099
rect 3709 16065 3743 16099
rect 3743 16065 3752 16099
rect 3700 16056 3752 16065
rect 3516 15988 3568 16040
rect 6920 16124 6972 16176
rect 4804 16099 4856 16108
rect 4804 16065 4813 16099
rect 4813 16065 4847 16099
rect 4847 16065 4856 16099
rect 4804 16056 4856 16065
rect 5264 16099 5316 16108
rect 5264 16065 5273 16099
rect 5273 16065 5307 16099
rect 5307 16065 5316 16099
rect 5264 16056 5316 16065
rect 5540 16056 5592 16108
rect 7564 16056 7616 16108
rect 10968 16124 11020 16176
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 5172 15852 5224 15904
rect 5540 15852 5592 15904
rect 6184 15895 6236 15904
rect 6184 15861 6193 15895
rect 6193 15861 6227 15895
rect 6227 15861 6236 15895
rect 6184 15852 6236 15861
rect 7196 15852 7248 15904
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 10140 16056 10192 16108
rect 14372 16056 14424 16108
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 10232 16031 10284 16040
rect 10232 15997 10241 16031
rect 10241 15997 10275 16031
rect 10275 15997 10284 16031
rect 10232 15988 10284 15997
rect 25136 15988 25188 16040
rect 7932 15895 7984 15904
rect 7932 15861 7941 15895
rect 7941 15861 7975 15895
rect 7975 15861 7984 15895
rect 7932 15852 7984 15861
rect 9036 15852 9088 15904
rect 9404 15852 9456 15904
rect 11428 15852 11480 15904
rect 13912 15852 13964 15904
rect 14464 15963 14516 15972
rect 14464 15929 14473 15963
rect 14473 15929 14507 15963
rect 14507 15929 14516 15963
rect 14464 15920 14516 15929
rect 14740 15852 14792 15904
rect 15108 15852 15160 15904
rect 18236 15963 18288 15972
rect 18236 15929 18245 15963
rect 18245 15929 18279 15963
rect 18279 15929 18288 15963
rect 18236 15920 18288 15929
rect 18696 15852 18748 15904
rect 25044 15852 25096 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 5540 15648 5592 15700
rect 8208 15691 8260 15700
rect 8208 15657 8217 15691
rect 8217 15657 8251 15691
rect 8251 15657 8260 15691
rect 8208 15648 8260 15657
rect 13912 15691 13964 15700
rect 13912 15657 13921 15691
rect 13921 15657 13955 15691
rect 13955 15657 13964 15691
rect 13912 15648 13964 15657
rect 14464 15648 14516 15700
rect 18236 15648 18288 15700
rect 4620 15580 4672 15632
rect 4528 15512 4580 15564
rect 6644 15555 6696 15564
rect 6644 15521 6653 15555
rect 6653 15521 6687 15555
rect 6687 15521 6696 15555
rect 6644 15512 6696 15521
rect 6920 15555 6972 15564
rect 6920 15521 6929 15555
rect 6929 15521 6963 15555
rect 6963 15521 6972 15555
rect 6920 15512 6972 15521
rect 8208 15555 8260 15564
rect 8208 15521 8217 15555
rect 8217 15521 8251 15555
rect 8251 15521 8260 15555
rect 8208 15512 8260 15521
rect 8392 15512 8444 15564
rect 8852 15512 8904 15564
rect 9036 15512 9088 15564
rect 11796 15512 11848 15564
rect 13728 15555 13780 15564
rect 13728 15521 13737 15555
rect 13737 15521 13771 15555
rect 13771 15521 13780 15555
rect 16120 15580 16172 15632
rect 18144 15623 18196 15632
rect 18144 15589 18153 15623
rect 18153 15589 18187 15623
rect 18187 15589 18196 15623
rect 18144 15580 18196 15589
rect 18696 15623 18748 15632
rect 18696 15589 18705 15623
rect 18705 15589 18739 15623
rect 18739 15589 18748 15623
rect 18696 15580 18748 15589
rect 24216 15580 24268 15632
rect 24860 15623 24912 15632
rect 24860 15589 24869 15623
rect 24869 15589 24903 15623
rect 24903 15589 24912 15623
rect 24860 15580 24912 15589
rect 13728 15512 13780 15521
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 11336 15444 11388 15496
rect 15844 15444 15896 15496
rect 17776 15444 17828 15496
rect 25044 15444 25096 15496
rect 5540 15376 5592 15428
rect 7656 15308 7708 15360
rect 10324 15351 10376 15360
rect 10324 15317 10333 15351
rect 10333 15317 10367 15351
rect 10367 15317 10376 15351
rect 10324 15308 10376 15317
rect 12440 15308 12492 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 6460 15147 6512 15156
rect 6460 15113 6469 15147
rect 6469 15113 6503 15147
rect 6503 15113 6512 15147
rect 6460 15104 6512 15113
rect 6644 15104 6696 15156
rect 8208 15104 8260 15156
rect 12808 15104 12860 15156
rect 13728 15104 13780 15156
rect 17776 15104 17828 15156
rect 25044 15147 25096 15156
rect 25044 15113 25053 15147
rect 25053 15113 25087 15147
rect 25087 15113 25096 15147
rect 25044 15104 25096 15113
rect 2964 14968 3016 15020
rect 8116 15079 8168 15088
rect 8116 15045 8125 15079
rect 8125 15045 8159 15079
rect 8159 15045 8168 15079
rect 8116 15036 8168 15045
rect 10048 15036 10100 15088
rect 5264 15011 5316 15020
rect 5264 14977 5273 15011
rect 5273 14977 5307 15011
rect 5307 14977 5316 15011
rect 5264 14968 5316 14977
rect 6368 14968 6420 15020
rect 7288 14968 7340 15020
rect 10324 15011 10376 15020
rect 10324 14977 10333 15011
rect 10333 14977 10367 15011
rect 10367 14977 10376 15011
rect 10324 14968 10376 14977
rect 4528 14900 4580 14952
rect 4068 14875 4120 14884
rect 4068 14841 4077 14875
rect 4077 14841 4111 14875
rect 4111 14841 4120 14875
rect 4068 14832 4120 14841
rect 5080 14875 5132 14884
rect 5080 14841 5089 14875
rect 5089 14841 5123 14875
rect 5123 14841 5132 14875
rect 5080 14832 5132 14841
rect 7656 14875 7708 14884
rect 7656 14841 7665 14875
rect 7665 14841 7699 14875
rect 7699 14841 7708 14875
rect 7656 14832 7708 14841
rect 12716 14900 12768 14952
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 6920 14764 6972 14816
rect 8668 14764 8720 14816
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 9404 14807 9456 14816
rect 9404 14773 9413 14807
rect 9413 14773 9447 14807
rect 9447 14773 9456 14807
rect 9404 14764 9456 14773
rect 9588 14764 9640 14816
rect 10692 14832 10744 14884
rect 13820 14900 13872 14952
rect 16120 15036 16172 15088
rect 18696 15079 18748 15088
rect 18696 15045 18705 15079
rect 18705 15045 18739 15079
rect 18739 15045 18748 15079
rect 18696 15036 18748 15045
rect 15844 14968 15896 15020
rect 16212 14832 16264 14884
rect 16580 14832 16632 14884
rect 24216 14968 24268 15020
rect 24032 14943 24084 14952
rect 24032 14909 24041 14943
rect 24041 14909 24075 14943
rect 24075 14909 24084 14943
rect 24032 14900 24084 14909
rect 18236 14875 18288 14884
rect 18236 14841 18245 14875
rect 18245 14841 18279 14875
rect 18279 14841 18288 14875
rect 18236 14832 18288 14841
rect 11796 14764 11848 14816
rect 15568 14807 15620 14816
rect 15568 14773 15577 14807
rect 15577 14773 15611 14807
rect 15611 14773 15620 14807
rect 15568 14764 15620 14773
rect 17040 14807 17092 14816
rect 17040 14773 17049 14807
rect 17049 14773 17083 14807
rect 17083 14773 17092 14807
rect 17040 14764 17092 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 4068 14560 4120 14612
rect 5080 14603 5132 14612
rect 5080 14569 5089 14603
rect 5089 14569 5123 14603
rect 5123 14569 5132 14603
rect 5080 14560 5132 14569
rect 5540 14603 5592 14612
rect 5540 14569 5549 14603
rect 5549 14569 5583 14603
rect 5583 14569 5592 14603
rect 5540 14560 5592 14569
rect 7656 14560 7708 14612
rect 12440 14603 12492 14612
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 12440 14560 12492 14569
rect 13820 14560 13872 14612
rect 16120 14603 16172 14612
rect 7288 14535 7340 14544
rect 7288 14501 7297 14535
rect 7297 14501 7331 14535
rect 7331 14501 7340 14535
rect 7288 14492 7340 14501
rect 7748 14535 7800 14544
rect 7748 14501 7757 14535
rect 7757 14501 7791 14535
rect 7791 14501 7800 14535
rect 7748 14492 7800 14501
rect 10048 14492 10100 14544
rect 11612 14535 11664 14544
rect 11612 14501 11621 14535
rect 11621 14501 11655 14535
rect 11655 14501 11664 14535
rect 11612 14492 11664 14501
rect 16120 14569 16129 14603
rect 16129 14569 16163 14603
rect 16163 14569 16172 14603
rect 16120 14560 16172 14569
rect 17040 14560 17092 14612
rect 18144 14560 18196 14612
rect 16672 14492 16724 14544
rect 18236 14492 18288 14544
rect 24124 14492 24176 14544
rect 24860 14492 24912 14544
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 4988 14424 5040 14476
rect 6000 14467 6052 14476
rect 6000 14433 6009 14467
rect 6009 14433 6043 14467
rect 6043 14433 6052 14467
rect 6000 14424 6052 14433
rect 7656 14424 7708 14476
rect 13084 14424 13136 14476
rect 13820 14424 13872 14476
rect 18420 14467 18472 14476
rect 18420 14433 18429 14467
rect 18429 14433 18463 14467
rect 18463 14433 18472 14467
rect 18420 14424 18472 14433
rect 7840 14356 7892 14408
rect 9864 14356 9916 14408
rect 11336 14356 11388 14408
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 16488 14356 16540 14408
rect 24860 14356 24912 14408
rect 4344 14263 4396 14272
rect 4344 14229 4353 14263
rect 4353 14229 4387 14263
rect 4387 14229 4396 14263
rect 4344 14220 4396 14229
rect 8392 14220 8444 14272
rect 9496 14220 9548 14272
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 17500 14263 17552 14272
rect 17500 14229 17509 14263
rect 17509 14229 17543 14263
rect 17543 14229 17552 14263
rect 17500 14220 17552 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1400 14016 1452 14068
rect 6000 14059 6052 14068
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 8208 14016 8260 14068
rect 10048 14059 10100 14068
rect 7840 13948 7892 14000
rect 8116 13991 8168 14000
rect 8116 13957 8125 13991
rect 8125 13957 8159 13991
rect 8159 13957 8168 13991
rect 8116 13948 8168 13957
rect 4436 13880 4488 13932
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 11336 14016 11388 14068
rect 16672 14059 16724 14068
rect 16672 14025 16681 14059
rect 16681 14025 16715 14059
rect 16715 14025 16724 14059
rect 16672 14016 16724 14025
rect 18420 14059 18472 14068
rect 18420 14025 18429 14059
rect 18429 14025 18463 14059
rect 18463 14025 18472 14059
rect 18420 14016 18472 14025
rect 11612 13923 11664 13932
rect 11612 13889 11621 13923
rect 11621 13889 11655 13923
rect 11655 13889 11664 13923
rect 11612 13880 11664 13889
rect 13176 13880 13228 13932
rect 13820 13880 13872 13932
rect 16488 13880 16540 13932
rect 9312 13812 9364 13864
rect 9496 13812 9548 13864
rect 10600 13812 10652 13864
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 13544 13855 13596 13864
rect 13544 13821 13553 13855
rect 13553 13821 13587 13855
rect 13587 13821 13596 13855
rect 13544 13812 13596 13821
rect 4068 13744 4120 13796
rect 4988 13744 5040 13796
rect 4620 13676 4672 13728
rect 7380 13744 7432 13796
rect 7656 13787 7708 13796
rect 7656 13753 7665 13787
rect 7665 13753 7699 13787
rect 7699 13753 7708 13787
rect 7656 13744 7708 13753
rect 9864 13744 9916 13796
rect 14372 13787 14424 13796
rect 14372 13753 14381 13787
rect 14381 13753 14415 13787
rect 14415 13753 14424 13787
rect 14372 13744 14424 13753
rect 12624 13719 12676 13728
rect 12624 13685 12633 13719
rect 12633 13685 12667 13719
rect 12667 13685 12676 13719
rect 12624 13676 12676 13685
rect 13084 13676 13136 13728
rect 14832 13676 14884 13728
rect 15476 13812 15528 13864
rect 15660 13812 15712 13864
rect 15844 13855 15896 13864
rect 15844 13821 15853 13855
rect 15853 13821 15887 13855
rect 15887 13821 15896 13855
rect 15844 13812 15896 13821
rect 24032 13719 24084 13728
rect 24032 13685 24041 13719
rect 24041 13685 24075 13719
rect 24075 13685 24084 13719
rect 24032 13676 24084 13685
rect 24860 13676 24912 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 7656 13472 7708 13524
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 9864 13515 9916 13524
rect 9864 13481 9873 13515
rect 9873 13481 9907 13515
rect 9907 13481 9916 13515
rect 9864 13472 9916 13481
rect 4344 13404 4396 13456
rect 7196 13447 7248 13456
rect 7196 13413 7205 13447
rect 7205 13413 7239 13447
rect 7239 13413 7248 13447
rect 13544 13472 13596 13524
rect 15568 13515 15620 13524
rect 15568 13481 15577 13515
rect 15577 13481 15611 13515
rect 15611 13481 15620 13515
rect 15568 13472 15620 13481
rect 7196 13404 7248 13413
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 6276 13336 6328 13345
rect 11888 13404 11940 13456
rect 12716 13447 12768 13456
rect 12716 13413 12725 13447
rect 12725 13413 12759 13447
rect 12759 13413 12768 13447
rect 12716 13404 12768 13413
rect 8392 13336 8444 13388
rect 11060 13379 11112 13388
rect 11060 13345 11069 13379
rect 11069 13345 11103 13379
rect 11103 13345 11112 13379
rect 11060 13336 11112 13345
rect 13636 13379 13688 13388
rect 13636 13345 13645 13379
rect 13645 13345 13679 13379
rect 13679 13345 13688 13379
rect 13636 13336 13688 13345
rect 14372 13336 14424 13388
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 15660 13336 15712 13388
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4436 13311 4488 13320
rect 4160 13268 4212 13277
rect 4436 13277 4445 13311
rect 4445 13277 4479 13311
rect 4479 13277 4488 13311
rect 4436 13268 4488 13277
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 9312 13200 9364 13252
rect 13084 13200 13136 13252
rect 8944 13132 8996 13184
rect 12256 13132 12308 13184
rect 12440 13132 12492 13184
rect 13176 13175 13228 13184
rect 13176 13141 13185 13175
rect 13185 13141 13219 13175
rect 13219 13141 13228 13175
rect 13176 13132 13228 13141
rect 13820 13175 13872 13184
rect 13820 13141 13829 13175
rect 13829 13141 13863 13175
rect 13863 13141 13872 13175
rect 13820 13132 13872 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 4344 12928 4396 12980
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 6276 12971 6328 12980
rect 6276 12937 6285 12971
rect 6285 12937 6319 12971
rect 6319 12937 6328 12971
rect 6276 12928 6328 12937
rect 8392 12928 8444 12980
rect 8760 12928 8812 12980
rect 10140 12928 10192 12980
rect 4068 12860 4120 12912
rect 1216 12792 1268 12844
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 8208 12860 8260 12912
rect 7564 12792 7616 12844
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 11888 12928 11940 12980
rect 13636 12928 13688 12980
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 15292 12971 15344 12980
rect 13820 12928 13872 12937
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 4712 12724 4764 12776
rect 4620 12656 4672 12708
rect 6276 12656 6328 12708
rect 3056 12588 3108 12640
rect 7288 12588 7340 12640
rect 10692 12724 10744 12776
rect 8944 12656 8996 12708
rect 12716 12792 12768 12844
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 14372 12835 14424 12844
rect 14372 12801 14381 12835
rect 14381 12801 14415 12835
rect 14415 12801 14424 12835
rect 14372 12792 14424 12801
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 12164 12656 12216 12708
rect 12256 12656 12308 12708
rect 12624 12699 12676 12708
rect 12624 12665 12633 12699
rect 12633 12665 12667 12699
rect 12667 12665 12676 12699
rect 12624 12656 12676 12665
rect 11060 12588 11112 12640
rect 13820 12588 13872 12640
rect 15660 12631 15712 12640
rect 15660 12597 15669 12631
rect 15669 12597 15703 12631
rect 15703 12597 15712 12631
rect 15660 12588 15712 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 4160 12384 4212 12436
rect 6276 12384 6328 12436
rect 12072 12384 12124 12436
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 14096 12384 14148 12436
rect 18144 12427 18196 12436
rect 18144 12393 18153 12427
rect 18153 12393 18187 12427
rect 18187 12393 18196 12427
rect 18144 12384 18196 12393
rect 19984 12384 20036 12436
rect 4620 12316 4672 12368
rect 5540 12316 5592 12368
rect 6736 12316 6788 12368
rect 7748 12316 7800 12368
rect 10692 12316 10744 12368
rect 13636 12316 13688 12368
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 9956 12248 10008 12300
rect 10876 12248 10928 12300
rect 15384 12291 15436 12300
rect 15384 12257 15393 12291
rect 15393 12257 15427 12291
rect 15427 12257 15436 12291
rect 15384 12248 15436 12257
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 6460 12180 6512 12232
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 9772 12180 9824 12232
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 12900 12112 12952 12164
rect 13728 12112 13780 12164
rect 14372 12112 14424 12164
rect 7196 12044 7248 12096
rect 8208 12044 8260 12096
rect 8576 12044 8628 12096
rect 9772 12044 9824 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 14280 12087 14332 12096
rect 14280 12053 14289 12087
rect 14289 12053 14323 12087
rect 14323 12053 14332 12087
rect 14280 12044 14332 12053
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 5540 11840 5592 11892
rect 6184 11840 6236 11892
rect 7748 11840 7800 11892
rect 7104 11772 7156 11824
rect 8576 11840 8628 11892
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 9772 11840 9824 11892
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 13636 11883 13688 11892
rect 13636 11849 13645 11883
rect 13645 11849 13679 11883
rect 13679 11849 13688 11883
rect 13636 11840 13688 11849
rect 15384 11840 15436 11892
rect 15752 11883 15804 11892
rect 15752 11849 15761 11883
rect 15761 11849 15795 11883
rect 15795 11849 15804 11883
rect 15752 11840 15804 11849
rect 8208 11772 8260 11824
rect 10692 11772 10744 11824
rect 6368 11704 6420 11756
rect 7840 11704 7892 11756
rect 16028 11704 16080 11756
rect 18144 11747 18196 11756
rect 18144 11713 18153 11747
rect 18153 11713 18187 11747
rect 18187 11713 18196 11747
rect 18144 11704 18196 11713
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 5540 11636 5592 11688
rect 8576 11636 8628 11688
rect 10140 11636 10192 11688
rect 7196 11568 7248 11620
rect 8944 11568 8996 11620
rect 10876 11568 10928 11620
rect 1400 11500 1452 11552
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 11520 11500 11572 11552
rect 14280 11636 14332 11688
rect 12164 11568 12216 11620
rect 13820 11500 13872 11552
rect 14556 11543 14608 11552
rect 14556 11509 14565 11543
rect 14565 11509 14599 11543
rect 14599 11509 14608 11543
rect 14556 11500 14608 11509
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 15752 11500 15804 11552
rect 17776 11543 17828 11552
rect 17776 11509 17785 11543
rect 17785 11509 17819 11543
rect 17819 11509 17828 11543
rect 17776 11500 17828 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 5448 11296 5500 11348
rect 6552 11296 6604 11348
rect 8760 11296 8812 11348
rect 9312 11296 9364 11348
rect 10140 11296 10192 11348
rect 12992 11339 13044 11348
rect 7196 11228 7248 11280
rect 8300 11228 8352 11280
rect 9680 11228 9732 11280
rect 10968 11228 11020 11280
rect 12992 11305 13001 11339
rect 13001 11305 13035 11339
rect 13035 11305 13044 11339
rect 12992 11296 13044 11305
rect 15384 11296 15436 11348
rect 15476 11339 15528 11348
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 17776 11339 17828 11348
rect 15476 11296 15528 11305
rect 17776 11305 17785 11339
rect 17785 11305 17819 11339
rect 17819 11305 17828 11339
rect 17776 11296 17828 11305
rect 14556 11228 14608 11280
rect 16304 11228 16356 11280
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 5172 11203 5224 11212
rect 5172 11169 5181 11203
rect 5181 11169 5215 11203
rect 5215 11169 5224 11203
rect 5172 11160 5224 11169
rect 5540 11160 5592 11212
rect 1584 11067 1636 11076
rect 1584 11033 1593 11067
rect 1593 11033 1627 11067
rect 1627 11033 1636 11067
rect 1584 11024 1636 11033
rect 9588 11160 9640 11212
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 12716 11160 12768 11212
rect 17592 11203 17644 11212
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 24676 11160 24728 11212
rect 11244 11092 11296 11144
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 8944 11067 8996 11076
rect 8944 11033 8953 11067
rect 8953 11033 8987 11067
rect 8987 11033 8996 11067
rect 8944 11024 8996 11033
rect 9772 11024 9824 11076
rect 10140 11024 10192 11076
rect 11428 11024 11480 11076
rect 11888 11024 11940 11076
rect 14096 11024 14148 11076
rect 6460 10999 6512 11008
rect 6460 10965 6469 10999
rect 6469 10965 6503 10999
rect 6503 10965 6512 10999
rect 6460 10956 6512 10965
rect 7288 10956 7340 11008
rect 8208 10956 8260 11008
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 8576 10956 8628 11008
rect 13636 10999 13688 11008
rect 13636 10965 13645 10999
rect 13645 10965 13679 10999
rect 13679 10965 13688 10999
rect 13636 10956 13688 10965
rect 23940 10956 23992 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1400 10752 1452 10804
rect 5172 10795 5224 10804
rect 5172 10761 5181 10795
rect 5181 10761 5215 10795
rect 5215 10761 5224 10795
rect 5172 10752 5224 10761
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 7840 10795 7892 10804
rect 7840 10761 7849 10795
rect 7849 10761 7883 10795
rect 7883 10761 7892 10795
rect 7840 10752 7892 10761
rect 8576 10795 8628 10804
rect 8576 10761 8585 10795
rect 8585 10761 8619 10795
rect 8619 10761 8628 10795
rect 8576 10752 8628 10761
rect 9588 10752 9640 10804
rect 11888 10795 11940 10804
rect 11888 10761 11897 10795
rect 11897 10761 11931 10795
rect 11931 10761 11940 10795
rect 11888 10752 11940 10761
rect 15752 10752 15804 10804
rect 17592 10795 17644 10804
rect 17592 10761 17601 10795
rect 17601 10761 17635 10795
rect 17635 10761 17644 10795
rect 17592 10752 17644 10761
rect 24676 10795 24728 10804
rect 24676 10761 24685 10795
rect 24685 10761 24719 10795
rect 24719 10761 24728 10795
rect 24676 10752 24728 10761
rect 7196 10684 7248 10736
rect 8760 10616 8812 10668
rect 11796 10616 11848 10668
rect 18420 10616 18472 10668
rect 6920 10412 6972 10464
rect 8484 10591 8536 10600
rect 8484 10557 8490 10591
rect 8490 10557 8536 10591
rect 8484 10548 8536 10557
rect 8300 10523 8352 10532
rect 8300 10489 8309 10523
rect 8309 10489 8343 10523
rect 8343 10489 8352 10523
rect 8300 10480 8352 10489
rect 7288 10412 7340 10464
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 9404 10455 9456 10464
rect 9404 10421 9413 10455
rect 9413 10421 9447 10455
rect 9447 10421 9456 10455
rect 9404 10412 9456 10421
rect 9772 10412 9824 10464
rect 11152 10548 11204 10600
rect 11428 10548 11480 10600
rect 11888 10548 11940 10600
rect 13452 10591 13504 10600
rect 13452 10557 13461 10591
rect 13461 10557 13495 10591
rect 13495 10557 13504 10591
rect 13452 10548 13504 10557
rect 14096 10591 14148 10600
rect 13636 10480 13688 10532
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14096 10548 14148 10557
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 15476 10523 15528 10532
rect 15476 10489 15485 10523
rect 15485 10489 15519 10523
rect 15519 10489 15528 10523
rect 15476 10480 15528 10489
rect 10784 10412 10836 10464
rect 12716 10455 12768 10464
rect 12716 10421 12725 10455
rect 12725 10421 12759 10455
rect 12759 10421 12768 10455
rect 12716 10412 12768 10421
rect 16304 10455 16356 10464
rect 16304 10421 16313 10455
rect 16313 10421 16347 10455
rect 16347 10421 16356 10455
rect 16304 10412 16356 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 6828 10251 6880 10260
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 8576 10208 8628 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 14280 10251 14332 10260
rect 14280 10217 14289 10251
rect 14289 10217 14323 10251
rect 14323 10217 14332 10251
rect 14280 10208 14332 10217
rect 23388 10208 23440 10260
rect 23940 10251 23992 10260
rect 23940 10217 23949 10251
rect 23949 10217 23983 10251
rect 23983 10217 23992 10251
rect 23940 10208 23992 10217
rect 7196 10140 7248 10192
rect 8852 10140 8904 10192
rect 9404 10140 9456 10192
rect 6644 10072 6696 10124
rect 7288 10072 7340 10124
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 7104 10004 7156 10056
rect 8208 10072 8260 10124
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 10876 10072 10928 10124
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 17592 10140 17644 10192
rect 18420 10140 18472 10192
rect 13452 10115 13504 10124
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 13636 10115 13688 10124
rect 13636 10081 13645 10115
rect 13645 10081 13679 10115
rect 13679 10081 13688 10115
rect 13636 10072 13688 10081
rect 14004 10115 14056 10124
rect 8116 10047 8168 10056
rect 6276 9936 6328 9988
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 9864 10004 9916 10056
rect 11612 10004 11664 10056
rect 14004 10081 14013 10115
rect 14013 10081 14047 10115
rect 14047 10081 14056 10115
rect 14004 10072 14056 10081
rect 14832 10072 14884 10124
rect 15660 10072 15712 10124
rect 15844 10115 15896 10124
rect 15844 10081 15853 10115
rect 15853 10081 15887 10115
rect 15887 10081 15896 10115
rect 15844 10072 15896 10081
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 8116 9868 8168 9920
rect 8760 9911 8812 9920
rect 8760 9877 8769 9911
rect 8769 9877 8803 9911
rect 8803 9877 8812 9911
rect 8760 9868 8812 9877
rect 12716 9868 12768 9920
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 6184 9664 6236 9716
rect 7840 9664 7892 9716
rect 8392 9707 8444 9716
rect 8392 9673 8401 9707
rect 8401 9673 8435 9707
rect 8435 9673 8444 9707
rect 8392 9664 8444 9673
rect 8484 9664 8536 9716
rect 10876 9707 10928 9716
rect 10876 9673 10885 9707
rect 10885 9673 10919 9707
rect 10919 9673 10928 9707
rect 10876 9664 10928 9673
rect 11244 9664 11296 9716
rect 13452 9707 13504 9716
rect 13452 9673 13461 9707
rect 13461 9673 13495 9707
rect 13495 9673 13504 9707
rect 13452 9664 13504 9673
rect 14004 9664 14056 9716
rect 14464 9707 14516 9716
rect 14464 9673 14473 9707
rect 14473 9673 14507 9707
rect 14507 9673 14516 9707
rect 14464 9664 14516 9673
rect 15660 9707 15712 9716
rect 15660 9673 15669 9707
rect 15669 9673 15703 9707
rect 15703 9673 15712 9707
rect 15660 9664 15712 9673
rect 17592 9664 17644 9716
rect 6276 9639 6328 9648
rect 6276 9605 6285 9639
rect 6285 9605 6319 9639
rect 6319 9605 6328 9639
rect 6276 9596 6328 9605
rect 6644 9639 6696 9648
rect 6644 9605 6653 9639
rect 6653 9605 6687 9639
rect 6687 9605 6696 9639
rect 6644 9596 6696 9605
rect 7196 9596 7248 9648
rect 8116 9639 8168 9648
rect 8116 9605 8140 9639
rect 8140 9605 8168 9639
rect 8116 9596 8168 9605
rect 8208 9639 8260 9648
rect 8208 9605 8217 9639
rect 8217 9605 8251 9639
rect 8251 9605 8260 9639
rect 8208 9596 8260 9605
rect 9128 9596 9180 9648
rect 10048 9596 10100 9648
rect 15752 9596 15804 9648
rect 8852 9528 8904 9580
rect 9404 9528 9456 9580
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 16120 9528 16172 9580
rect 23388 9528 23440 9580
rect 6552 9460 6604 9512
rect 7104 9460 7156 9512
rect 8024 9460 8076 9512
rect 8760 9460 8812 9512
rect 9680 9460 9732 9512
rect 14464 9460 14516 9512
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 15844 9460 15896 9512
rect 19064 9460 19116 9512
rect 7196 9392 7248 9444
rect 9772 9392 9824 9444
rect 12624 9435 12676 9444
rect 12624 9401 12633 9435
rect 12633 9401 12667 9435
rect 12667 9401 12676 9435
rect 12624 9392 12676 9401
rect 16212 9392 16264 9444
rect 16304 9392 16356 9444
rect 17408 9392 17460 9444
rect 18052 9435 18104 9444
rect 18052 9401 18061 9435
rect 18061 9401 18095 9435
rect 18095 9401 18104 9435
rect 18052 9392 18104 9401
rect 24584 9435 24636 9444
rect 7932 9324 7984 9376
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 23388 9367 23440 9376
rect 23388 9333 23397 9367
rect 23397 9333 23431 9367
rect 23431 9333 23440 9367
rect 24584 9401 24593 9435
rect 24593 9401 24627 9435
rect 24627 9401 24636 9435
rect 24584 9392 24636 9401
rect 23388 9324 23440 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 6184 9163 6236 9172
rect 6184 9129 6193 9163
rect 6193 9129 6227 9163
rect 6227 9129 6236 9163
rect 6184 9120 6236 9129
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 9772 9120 9824 9172
rect 8024 9095 8076 9104
rect 8024 9061 8033 9095
rect 8033 9061 8067 9095
rect 8067 9061 8076 9095
rect 8024 9052 8076 9061
rect 1676 8984 1728 9036
rect 2596 8984 2648 9036
rect 6092 8984 6144 9036
rect 7012 9027 7064 9036
rect 7012 8993 7021 9027
rect 7021 8993 7055 9027
rect 7055 8993 7064 9027
rect 7012 8984 7064 8993
rect 7104 8916 7156 8968
rect 8208 8984 8260 9036
rect 10048 9120 10100 9172
rect 10600 9027 10652 9036
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 8024 8916 8076 8968
rect 12440 9120 12492 9172
rect 11888 9052 11940 9104
rect 13820 9120 13872 9172
rect 16120 9120 16172 9172
rect 13636 9052 13688 9104
rect 17408 9052 17460 9104
rect 19524 9120 19576 9172
rect 24492 9120 24544 9172
rect 24860 9120 24912 9172
rect 19064 9052 19116 9104
rect 24032 9095 24084 9104
rect 24032 9061 24041 9095
rect 24041 9061 24075 9095
rect 24075 9061 24084 9095
rect 24032 9052 24084 9061
rect 11612 8984 11664 9036
rect 14464 8984 14516 9036
rect 15476 8984 15528 9036
rect 15752 9027 15804 9036
rect 15752 8993 15761 9027
rect 15761 8993 15795 9027
rect 15795 8993 15804 9027
rect 15752 8984 15804 8993
rect 16212 8984 16264 9036
rect 16764 8984 16816 9036
rect 22928 8984 22980 9036
rect 24584 9027 24636 9036
rect 24584 8993 24593 9027
rect 24593 8993 24627 9027
rect 24627 8993 24636 9027
rect 25504 9027 25556 9036
rect 24584 8984 24636 8993
rect 25504 8993 25522 9027
rect 25522 8993 25556 9027
rect 25504 8984 25556 8993
rect 27620 8984 27672 9036
rect 13452 8916 13504 8968
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 18788 8916 18840 8968
rect 23940 8959 23992 8968
rect 23940 8925 23949 8959
rect 23949 8925 23983 8959
rect 23983 8925 23992 8959
rect 23940 8916 23992 8925
rect 1584 8891 1636 8900
rect 1584 8857 1593 8891
rect 1593 8857 1627 8891
rect 1627 8857 1636 8891
rect 1584 8848 1636 8857
rect 7564 8848 7616 8900
rect 9128 8848 9180 8900
rect 15108 8848 15160 8900
rect 23388 8848 23440 8900
rect 1676 8780 1728 8832
rect 6552 8823 6604 8832
rect 6552 8789 6561 8823
rect 6561 8789 6595 8823
rect 6595 8789 6604 8823
rect 6552 8780 6604 8789
rect 8116 8780 8168 8832
rect 12624 8780 12676 8832
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 22836 8780 22888 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 7564 8576 7616 8628
rect 7840 8576 7892 8628
rect 8300 8576 8352 8628
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 14464 8576 14516 8628
rect 9128 8440 9180 8492
rect 11428 8508 11480 8560
rect 11520 8483 11572 8492
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 8116 8372 8168 8424
rect 8484 8372 8536 8424
rect 10876 8415 10928 8424
rect 10876 8381 10885 8415
rect 10885 8381 10919 8415
rect 10919 8381 10928 8415
rect 10876 8372 10928 8381
rect 11244 8372 11296 8424
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 15660 8576 15712 8628
rect 16764 8619 16816 8628
rect 16764 8585 16773 8619
rect 16773 8585 16807 8619
rect 16807 8585 16816 8619
rect 16764 8576 16816 8585
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 18052 8576 18104 8628
rect 19064 8619 19116 8628
rect 19064 8585 19073 8619
rect 19073 8585 19107 8619
rect 19107 8585 19116 8619
rect 19064 8576 19116 8585
rect 19524 8619 19576 8628
rect 19524 8585 19533 8619
rect 19533 8585 19567 8619
rect 19567 8585 19576 8619
rect 19524 8576 19576 8585
rect 22928 8619 22980 8628
rect 22928 8585 22937 8619
rect 22937 8585 22971 8619
rect 22971 8585 22980 8619
rect 22928 8576 22980 8585
rect 23388 8619 23440 8628
rect 23388 8585 23397 8619
rect 23397 8585 23431 8619
rect 23431 8585 23440 8619
rect 23388 8576 23440 8585
rect 25504 8619 25556 8628
rect 25504 8585 25513 8619
rect 25513 8585 25547 8619
rect 25547 8585 25556 8619
rect 25504 8576 25556 8585
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 18788 8440 18840 8449
rect 24032 8440 24084 8492
rect 6552 8304 6604 8356
rect 7564 8304 7616 8356
rect 8208 8347 8260 8356
rect 8208 8313 8217 8347
rect 8217 8313 8251 8347
rect 8251 8313 8260 8347
rect 8208 8304 8260 8313
rect 8944 8347 8996 8356
rect 8944 8313 8953 8347
rect 8953 8313 8987 8347
rect 8987 8313 8996 8347
rect 8944 8304 8996 8313
rect 11980 8304 12032 8356
rect 2596 8279 2648 8288
rect 2596 8245 2605 8279
rect 2605 8245 2639 8279
rect 2639 8245 2648 8279
rect 2596 8236 2648 8245
rect 6092 8279 6144 8288
rect 6092 8245 6101 8279
rect 6101 8245 6135 8279
rect 6135 8245 6144 8279
rect 6092 8236 6144 8245
rect 8024 8279 8076 8288
rect 8024 8245 8033 8279
rect 8033 8245 8067 8279
rect 8067 8245 8076 8279
rect 8024 8236 8076 8245
rect 11888 8236 11940 8288
rect 12716 8236 12768 8288
rect 13636 8236 13688 8288
rect 15752 8415 15804 8424
rect 15752 8381 15761 8415
rect 15761 8381 15795 8415
rect 15795 8381 15804 8415
rect 15752 8372 15804 8381
rect 23388 8372 23440 8424
rect 16672 8304 16724 8356
rect 18144 8304 18196 8356
rect 23940 8304 23992 8356
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 7196 8032 7248 8041
rect 8760 8075 8812 8084
rect 8760 8041 8769 8075
rect 8769 8041 8803 8075
rect 8803 8041 8812 8075
rect 8760 8032 8812 8041
rect 11152 8032 11204 8084
rect 12624 8032 12676 8084
rect 15752 8032 15804 8084
rect 23940 8032 23992 8084
rect 11980 8007 12032 8016
rect 11980 7973 11989 8007
rect 11989 7973 12023 8007
rect 12023 7973 12032 8007
rect 11980 7964 12032 7973
rect 15476 7964 15528 8016
rect 16396 7964 16448 8016
rect 6276 7896 6328 7948
rect 6092 7828 6144 7880
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 8024 7896 8076 7948
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 11612 7896 11664 7948
rect 12532 7939 12584 7948
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 12532 7896 12584 7905
rect 12808 7896 12860 7948
rect 13452 7939 13504 7948
rect 13452 7905 13461 7939
rect 13461 7905 13495 7939
rect 13495 7905 13504 7939
rect 13452 7896 13504 7905
rect 16028 7896 16080 7948
rect 18236 7939 18288 7948
rect 18236 7905 18245 7939
rect 18245 7905 18279 7939
rect 18279 7905 18288 7939
rect 18236 7896 18288 7905
rect 24768 7896 24820 7948
rect 8484 7871 8536 7880
rect 6552 7828 6604 7837
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 11336 7828 11388 7880
rect 12164 7828 12216 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 7012 7760 7064 7812
rect 17776 7760 17828 7812
rect 22284 7760 22336 7812
rect 6644 7692 6696 7744
rect 6828 7735 6880 7744
rect 6828 7701 6837 7735
rect 6837 7701 6871 7735
rect 6871 7701 6880 7735
rect 6828 7692 6880 7701
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 10876 7692 10928 7744
rect 18328 7735 18380 7744
rect 18328 7701 18337 7735
rect 18337 7701 18371 7735
rect 18371 7701 18380 7735
rect 18328 7692 18380 7701
rect 23756 7735 23808 7744
rect 23756 7701 23765 7735
rect 23765 7701 23799 7735
rect 23799 7701 23808 7735
rect 23756 7692 23808 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 6828 7488 6880 7540
rect 9680 7488 9732 7540
rect 10692 7531 10744 7540
rect 10692 7497 10701 7531
rect 10701 7497 10735 7531
rect 10735 7497 10744 7531
rect 10692 7488 10744 7497
rect 11980 7488 12032 7540
rect 12164 7531 12216 7540
rect 12164 7497 12173 7531
rect 12173 7497 12207 7531
rect 12207 7497 12216 7531
rect 12164 7488 12216 7497
rect 13452 7531 13504 7540
rect 13452 7497 13461 7531
rect 13461 7497 13495 7531
rect 13495 7497 13504 7531
rect 13452 7488 13504 7497
rect 16028 7488 16080 7540
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 6644 7420 6696 7472
rect 8944 7352 8996 7404
rect 13728 7352 13780 7404
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 18512 7395 18564 7404
rect 18512 7361 18521 7395
rect 18521 7361 18555 7395
rect 18555 7361 18564 7395
rect 18512 7352 18564 7361
rect 23756 7395 23808 7404
rect 112 7284 164 7336
rect 5080 7284 5132 7336
rect 6552 7327 6604 7336
rect 6552 7293 6561 7327
rect 6561 7293 6595 7327
rect 6595 7293 6604 7327
rect 6552 7284 6604 7293
rect 7196 7284 7248 7336
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 8484 7284 8536 7336
rect 10048 7284 10100 7336
rect 10692 7284 10744 7336
rect 11244 7327 11296 7336
rect 11244 7293 11253 7327
rect 11253 7293 11287 7327
rect 11287 7293 11296 7327
rect 11244 7284 11296 7293
rect 14832 7284 14884 7336
rect 6276 7216 6328 7268
rect 11520 7259 11572 7268
rect 11520 7225 11529 7259
rect 11529 7225 11563 7259
rect 11563 7225 11572 7259
rect 11520 7216 11572 7225
rect 14648 7259 14700 7268
rect 7012 7191 7064 7200
rect 7012 7157 7021 7191
rect 7021 7157 7055 7191
rect 7055 7157 7064 7191
rect 7012 7148 7064 7157
rect 9404 7148 9456 7200
rect 13452 7148 13504 7200
rect 14648 7225 14657 7259
rect 14657 7225 14691 7259
rect 14691 7225 14700 7259
rect 14648 7216 14700 7225
rect 18236 7259 18288 7268
rect 18236 7225 18245 7259
rect 18245 7225 18279 7259
rect 18279 7225 18288 7259
rect 18236 7216 18288 7225
rect 22100 7216 22152 7268
rect 23756 7361 23765 7395
rect 23765 7361 23799 7395
rect 23799 7361 23808 7395
rect 23756 7352 23808 7361
rect 23940 7352 23992 7404
rect 23848 7259 23900 7268
rect 23848 7225 23857 7259
rect 23857 7225 23891 7259
rect 23891 7225 23900 7259
rect 23848 7216 23900 7225
rect 14832 7148 14884 7200
rect 15384 7191 15436 7200
rect 15384 7157 15393 7191
rect 15393 7157 15427 7191
rect 15427 7157 15436 7191
rect 15384 7148 15436 7157
rect 16304 7191 16356 7200
rect 16304 7157 16313 7191
rect 16313 7157 16347 7191
rect 16347 7157 16356 7191
rect 16304 7148 16356 7157
rect 24768 7191 24820 7200
rect 24768 7157 24777 7191
rect 24777 7157 24811 7191
rect 24811 7157 24820 7191
rect 24768 7148 24820 7157
rect 25504 7148 25556 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 7932 6944 7984 6996
rect 8392 6944 8444 6996
rect 11244 6987 11296 6996
rect 11244 6953 11253 6987
rect 11253 6953 11287 6987
rect 11287 6953 11296 6987
rect 11244 6944 11296 6953
rect 13452 6944 13504 6996
rect 13728 6944 13780 6996
rect 15384 6944 15436 6996
rect 18236 6944 18288 6996
rect 7012 6876 7064 6928
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 6276 6808 6328 6860
rect 7656 6851 7708 6860
rect 7656 6817 7665 6851
rect 7665 6817 7699 6851
rect 7699 6817 7708 6851
rect 7656 6808 7708 6817
rect 11888 6876 11940 6928
rect 16304 6876 16356 6928
rect 18512 6919 18564 6928
rect 18512 6885 18521 6919
rect 18521 6885 18555 6919
rect 18555 6885 18564 6919
rect 18512 6876 18564 6885
rect 22836 6944 22888 6996
rect 19616 6876 19668 6928
rect 23020 6919 23072 6928
rect 23020 6885 23029 6919
rect 23029 6885 23063 6919
rect 23063 6885 23072 6919
rect 23020 6876 23072 6885
rect 23848 6876 23900 6928
rect 9680 6851 9732 6860
rect 9680 6817 9689 6851
rect 9689 6817 9723 6851
rect 9723 6817 9732 6851
rect 9680 6808 9732 6817
rect 16672 6851 16724 6860
rect 16672 6817 16681 6851
rect 16681 6817 16715 6851
rect 16715 6817 16724 6851
rect 16672 6808 16724 6817
rect 18236 6808 18288 6860
rect 24676 6851 24728 6860
rect 24676 6817 24685 6851
rect 24685 6817 24719 6851
rect 24719 6817 24728 6851
rect 24676 6808 24728 6817
rect 7104 6740 7156 6792
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 11520 6740 11572 6792
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 19156 6783 19208 6792
rect 19156 6749 19165 6783
rect 19165 6749 19199 6783
rect 19199 6749 19208 6783
rect 19156 6740 19208 6749
rect 24032 6740 24084 6792
rect 8392 6672 8444 6724
rect 9956 6715 10008 6724
rect 9956 6681 9965 6715
rect 9965 6681 9999 6715
rect 9999 6681 10008 6715
rect 9956 6672 10008 6681
rect 9496 6604 9548 6656
rect 10876 6647 10928 6656
rect 10876 6613 10885 6647
rect 10885 6613 10919 6647
rect 10919 6613 10928 6647
rect 10876 6604 10928 6613
rect 23848 6647 23900 6656
rect 23848 6613 23857 6647
rect 23857 6613 23891 6647
rect 23891 6613 23900 6647
rect 23848 6604 23900 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 8024 6400 8076 6452
rect 9496 6400 9548 6452
rect 10048 6400 10100 6452
rect 11520 6400 11572 6452
rect 13360 6443 13412 6452
rect 13360 6409 13369 6443
rect 13369 6409 13403 6443
rect 13403 6409 13412 6443
rect 13360 6400 13412 6409
rect 8392 6375 8444 6384
rect 8392 6341 8401 6375
rect 8401 6341 8435 6375
rect 8435 6341 8444 6375
rect 8392 6332 8444 6341
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 9956 6264 10008 6316
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 8024 6196 8076 6248
rect 8760 6196 8812 6248
rect 10876 6332 10928 6384
rect 14832 6400 14884 6452
rect 16672 6400 16724 6452
rect 19616 6443 19668 6452
rect 14096 6375 14148 6384
rect 14096 6341 14105 6375
rect 14105 6341 14139 6375
rect 14139 6341 14148 6375
rect 14096 6332 14148 6341
rect 13544 6264 13596 6316
rect 14004 6264 14056 6316
rect 15384 6264 15436 6316
rect 19156 6332 19208 6384
rect 19616 6409 19625 6443
rect 19625 6409 19659 6443
rect 19659 6409 19668 6443
rect 19616 6400 19668 6409
rect 24676 6443 24728 6452
rect 24676 6409 24685 6443
rect 24685 6409 24719 6443
rect 24719 6409 24728 6443
rect 24676 6400 24728 6409
rect 25596 6400 25648 6452
rect 17592 6264 17644 6316
rect 10968 6196 11020 6248
rect 23388 6332 23440 6384
rect 6644 6128 6696 6180
rect 7012 6128 7064 6180
rect 12716 6128 12768 6180
rect 23020 6239 23072 6248
rect 23020 6205 23029 6239
rect 23029 6205 23063 6239
rect 23063 6205 23072 6239
rect 23020 6196 23072 6205
rect 13544 6171 13596 6180
rect 13544 6137 13553 6171
rect 13553 6137 13587 6171
rect 13587 6137 13596 6171
rect 13544 6128 13596 6137
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 7564 6060 7616 6112
rect 8116 6060 8168 6112
rect 8208 6060 8260 6112
rect 8392 6060 8444 6112
rect 9680 6103 9732 6112
rect 9680 6069 9689 6103
rect 9689 6069 9723 6103
rect 9723 6069 9732 6103
rect 9680 6060 9732 6069
rect 11060 6103 11112 6112
rect 11060 6069 11069 6103
rect 11069 6069 11103 6103
rect 11103 6069 11112 6103
rect 11060 6060 11112 6069
rect 11888 6060 11940 6112
rect 12992 6103 13044 6112
rect 12992 6069 13001 6103
rect 13001 6069 13035 6103
rect 13035 6069 13044 6103
rect 12992 6060 13044 6069
rect 13360 6060 13412 6112
rect 16304 6128 16356 6180
rect 23848 6264 23900 6316
rect 24032 6307 24084 6316
rect 24032 6273 24041 6307
rect 24041 6273 24075 6307
rect 24075 6273 24084 6307
rect 24032 6264 24084 6273
rect 25228 6239 25280 6248
rect 25228 6205 25237 6239
rect 25237 6205 25271 6239
rect 25271 6205 25280 6239
rect 25228 6196 25280 6205
rect 15476 6103 15528 6112
rect 15476 6069 15485 6103
rect 15485 6069 15519 6103
rect 15519 6069 15528 6103
rect 15476 6060 15528 6069
rect 18420 6103 18472 6112
rect 18420 6069 18429 6103
rect 18429 6069 18463 6103
rect 18463 6069 18472 6103
rect 18420 6060 18472 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 6920 5856 6972 5908
rect 7656 5856 7708 5908
rect 8484 5856 8536 5908
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 11612 5856 11664 5908
rect 13544 5899 13596 5908
rect 8024 5831 8076 5840
rect 8024 5797 8033 5831
rect 8033 5797 8067 5831
rect 8067 5797 8076 5831
rect 8024 5788 8076 5797
rect 9956 5788 10008 5840
rect 11796 5831 11848 5840
rect 11796 5797 11805 5831
rect 11805 5797 11839 5831
rect 11839 5797 11848 5831
rect 11796 5788 11848 5797
rect 6184 5720 6236 5772
rect 6644 5720 6696 5772
rect 7748 5652 7800 5704
rect 9404 5720 9456 5772
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 13544 5856 13596 5865
rect 22100 5899 22152 5908
rect 12992 5788 13044 5840
rect 13728 5788 13780 5840
rect 15476 5788 15528 5840
rect 18328 5788 18380 5840
rect 22100 5865 22109 5899
rect 22109 5865 22143 5899
rect 22143 5865 22152 5899
rect 22100 5856 22152 5865
rect 22836 5899 22888 5908
rect 22836 5865 22845 5899
rect 22845 5865 22879 5899
rect 22879 5865 22888 5899
rect 22836 5856 22888 5865
rect 25228 5856 25280 5908
rect 23388 5788 23440 5840
rect 23940 5788 23992 5840
rect 13084 5720 13136 5772
rect 9772 5652 9824 5704
rect 12072 5652 12124 5704
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 12716 5652 12768 5704
rect 14648 5720 14700 5772
rect 25412 5720 25464 5772
rect 16580 5652 16632 5704
rect 8116 5584 8168 5636
rect 8300 5627 8352 5636
rect 8300 5593 8309 5627
rect 8309 5593 8343 5627
rect 8343 5593 8352 5627
rect 8300 5584 8352 5593
rect 18512 5652 18564 5704
rect 24032 5652 24084 5704
rect 9036 5559 9088 5568
rect 9036 5525 9045 5559
rect 9045 5525 9079 5559
rect 9079 5525 9088 5559
rect 9036 5516 9088 5525
rect 10692 5516 10744 5568
rect 10968 5516 11020 5568
rect 18604 5516 18656 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 8300 5355 8352 5364
rect 8300 5321 8309 5355
rect 8309 5321 8343 5355
rect 8343 5321 8352 5355
rect 8300 5312 8352 5321
rect 9404 5355 9456 5364
rect 9404 5321 9413 5355
rect 9413 5321 9447 5355
rect 9447 5321 9456 5355
rect 9404 5312 9456 5321
rect 9864 5312 9916 5364
rect 12716 5355 12768 5364
rect 12716 5321 12725 5355
rect 12725 5321 12759 5355
rect 12759 5321 12768 5355
rect 12716 5312 12768 5321
rect 13084 5355 13136 5364
rect 13084 5321 13093 5355
rect 13093 5321 13127 5355
rect 13127 5321 13136 5355
rect 13084 5312 13136 5321
rect 8024 5176 8076 5228
rect 12164 5244 12216 5296
rect 10692 5176 10744 5228
rect 11796 5176 11848 5228
rect 12072 5219 12124 5228
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 6736 5108 6788 5160
rect 8116 5108 8168 5160
rect 9036 5108 9088 5160
rect 15476 5312 15528 5364
rect 16580 5355 16632 5364
rect 16580 5321 16589 5355
rect 16589 5321 16623 5355
rect 16623 5321 16632 5355
rect 16580 5312 16632 5321
rect 18420 5355 18472 5364
rect 18420 5321 18429 5355
rect 18429 5321 18463 5355
rect 18463 5321 18472 5355
rect 18420 5312 18472 5321
rect 23848 5312 23900 5364
rect 24032 5312 24084 5364
rect 25412 5355 25464 5364
rect 25412 5321 25421 5355
rect 25421 5321 25455 5355
rect 25455 5321 25464 5355
rect 25412 5312 25464 5321
rect 14832 5244 14884 5296
rect 14096 5151 14148 5160
rect 14096 5117 14105 5151
rect 14105 5117 14139 5151
rect 14139 5117 14148 5151
rect 18328 5244 18380 5296
rect 23388 5287 23440 5296
rect 23388 5253 23397 5287
rect 23397 5253 23431 5287
rect 23431 5253 23440 5287
rect 23388 5244 23440 5253
rect 14096 5108 14148 5117
rect 18236 5151 18288 5160
rect 6828 5083 6880 5092
rect 6828 5049 6837 5083
rect 6837 5049 6871 5083
rect 6871 5049 6880 5083
rect 6828 5040 6880 5049
rect 8392 5083 8444 5092
rect 8392 5049 8401 5083
rect 8401 5049 8435 5083
rect 8435 5049 8444 5083
rect 8392 5040 8444 5049
rect 9128 5083 9180 5092
rect 9128 5049 9137 5083
rect 9137 5049 9171 5083
rect 9171 5049 9180 5083
rect 9128 5040 9180 5049
rect 10232 5083 10284 5092
rect 10232 5049 10241 5083
rect 10241 5049 10275 5083
rect 10275 5049 10284 5083
rect 10232 5040 10284 5049
rect 14372 5083 14424 5092
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 9864 5015 9916 5024
rect 9864 4981 9873 5015
rect 9873 4981 9907 5015
rect 9907 4981 9916 5015
rect 9864 4972 9916 4981
rect 9956 4972 10008 5024
rect 14372 5049 14381 5083
rect 14381 5049 14415 5083
rect 14415 5049 14424 5083
rect 14372 5040 14424 5049
rect 18236 5117 18245 5151
rect 18245 5117 18279 5151
rect 18279 5117 18288 5151
rect 18236 5108 18288 5117
rect 19156 5108 19208 5160
rect 24124 5040 24176 5092
rect 27620 5040 27672 5092
rect 15292 5015 15344 5024
rect 15292 4981 15301 5015
rect 15301 4981 15335 5015
rect 15335 4981 15344 5015
rect 15292 4972 15344 4981
rect 19984 4972 20036 5024
rect 24032 4972 24084 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 6828 4768 6880 4820
rect 7748 4811 7800 4820
rect 7748 4777 7757 4811
rect 7757 4777 7791 4811
rect 7791 4777 7800 4811
rect 7748 4768 7800 4777
rect 8024 4768 8076 4820
rect 9128 4768 9180 4820
rect 10968 4768 11020 4820
rect 11244 4768 11296 4820
rect 14096 4768 14148 4820
rect 18236 4811 18288 4820
rect 18236 4777 18245 4811
rect 18245 4777 18279 4811
rect 18279 4777 18288 4811
rect 18236 4768 18288 4777
rect 8300 4700 8352 4752
rect 9864 4700 9916 4752
rect 11796 4700 11848 4752
rect 15476 4700 15528 4752
rect 17224 4743 17276 4752
rect 17224 4709 17233 4743
rect 17233 4709 17267 4743
rect 17267 4709 17276 4743
rect 17224 4700 17276 4709
rect 1584 4632 1636 4684
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 6736 4632 6788 4684
rect 11060 4675 11112 4684
rect 11060 4641 11069 4675
rect 11069 4641 11103 4675
rect 11103 4641 11112 4675
rect 11060 4632 11112 4641
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 18604 4675 18656 4684
rect 18604 4641 18613 4675
rect 18613 4641 18647 4675
rect 18647 4641 18656 4675
rect 18604 4632 18656 4641
rect 19984 4632 20036 4684
rect 8392 4564 8444 4616
rect 17776 4564 17828 4616
rect 10232 4496 10284 4548
rect 14556 4496 14608 4548
rect 17684 4539 17736 4548
rect 17684 4505 17693 4539
rect 17693 4505 17727 4539
rect 17727 4505 17736 4539
rect 17684 4496 17736 4505
rect 9956 4428 10008 4480
rect 11980 4471 12032 4480
rect 11980 4437 11989 4471
rect 11989 4437 12023 4471
rect 12023 4437 12032 4471
rect 11980 4428 12032 4437
rect 16488 4428 16540 4480
rect 21364 4428 21416 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1584 4267 1636 4276
rect 1584 4233 1593 4267
rect 1593 4233 1627 4267
rect 1627 4233 1636 4267
rect 1584 4224 1636 4233
rect 6828 4224 6880 4276
rect 8116 4267 8168 4276
rect 8116 4233 8125 4267
rect 8125 4233 8159 4267
rect 8159 4233 8168 4267
rect 8116 4224 8168 4233
rect 10232 4267 10284 4276
rect 10232 4233 10241 4267
rect 10241 4233 10275 4267
rect 10275 4233 10284 4267
rect 10232 4224 10284 4233
rect 3792 4156 3844 4208
rect 6736 4156 6788 4208
rect 8300 4156 8352 4208
rect 10140 4156 10192 4208
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 6276 4020 6328 4072
rect 6828 4020 6880 4072
rect 10692 4020 10744 4072
rect 11612 4224 11664 4276
rect 10876 4156 10928 4208
rect 17776 4199 17828 4208
rect 17776 4165 17785 4199
rect 17785 4165 17819 4199
rect 17819 4165 17828 4199
rect 17776 4156 17828 4165
rect 11796 4088 11848 4140
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 11244 4020 11296 4029
rect 11980 4020 12032 4072
rect 13452 4020 13504 4072
rect 11428 3952 11480 4004
rect 12440 3995 12492 4004
rect 12440 3961 12449 3995
rect 12449 3961 12483 3995
rect 12483 3961 12492 3995
rect 12440 3952 12492 3961
rect 14464 4063 14516 4072
rect 14464 4029 14473 4063
rect 14473 4029 14507 4063
rect 14507 4029 14516 4063
rect 14464 4020 14516 4029
rect 16488 4063 16540 4072
rect 16488 4029 16497 4063
rect 16497 4029 16531 4063
rect 16531 4029 16540 4063
rect 16488 4020 16540 4029
rect 18788 4224 18840 4276
rect 19984 4224 20036 4276
rect 24860 4267 24912 4276
rect 24860 4233 24869 4267
rect 24869 4233 24903 4267
rect 24903 4233 24912 4267
rect 24860 4224 24912 4233
rect 15476 3952 15528 4004
rect 17224 3952 17276 4004
rect 572 3884 624 3936
rect 6276 3884 6328 3936
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 12164 3884 12216 3936
rect 13268 3884 13320 3936
rect 15384 3927 15436 3936
rect 15384 3893 15393 3927
rect 15393 3893 15427 3927
rect 15427 3893 15436 3927
rect 15384 3884 15436 3893
rect 26884 3884 26936 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 11060 3723 11112 3732
rect 11060 3689 11069 3723
rect 11069 3689 11103 3723
rect 11103 3689 11112 3723
rect 11060 3680 11112 3689
rect 11796 3723 11848 3732
rect 11796 3689 11805 3723
rect 11805 3689 11839 3723
rect 11839 3689 11848 3723
rect 11796 3680 11848 3689
rect 14464 3723 14516 3732
rect 14464 3689 14473 3723
rect 14473 3689 14507 3723
rect 14507 3689 14516 3723
rect 14464 3680 14516 3689
rect 15292 3680 15344 3732
rect 13084 3612 13136 3664
rect 13268 3655 13320 3664
rect 13268 3621 13277 3655
rect 13277 3621 13311 3655
rect 13311 3621 13320 3655
rect 13268 3612 13320 3621
rect 13452 3612 13504 3664
rect 16488 3655 16540 3664
rect 16488 3621 16497 3655
rect 16497 3621 16531 3655
rect 16531 3621 16540 3655
rect 16488 3612 16540 3621
rect 16672 3612 16724 3664
rect 17684 3612 17736 3664
rect 5264 3544 5316 3596
rect 6000 3544 6052 3596
rect 18512 3587 18564 3596
rect 18512 3553 18521 3587
rect 18521 3553 18555 3587
rect 18555 3553 18564 3587
rect 18512 3544 18564 3553
rect 10692 3476 10744 3528
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 16580 3476 16632 3528
rect 10968 3340 11020 3392
rect 12348 3383 12400 3392
rect 12348 3349 12357 3383
rect 12357 3349 12391 3383
rect 12391 3349 12400 3383
rect 12348 3340 12400 3349
rect 12532 3340 12584 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 6000 3179 6052 3188
rect 6000 3145 6009 3179
rect 6009 3145 6043 3179
rect 6043 3145 6052 3179
rect 6000 3136 6052 3145
rect 6460 3136 6512 3188
rect 9956 3136 10008 3188
rect 12164 3136 12216 3188
rect 12440 3136 12492 3188
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 16488 3179 16540 3188
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 18512 3179 18564 3188
rect 18512 3145 18521 3179
rect 18521 3145 18555 3179
rect 18555 3145 18564 3179
rect 18512 3136 18564 3145
rect 13084 3068 13136 3120
rect 204 3000 256 3052
rect 13544 3000 13596 3052
rect 8668 2796 8720 2848
rect 12348 2932 12400 2984
rect 13268 2932 13320 2984
rect 16672 3000 16724 3052
rect 17592 3000 17644 3052
rect 16212 2975 16264 2984
rect 16212 2941 16221 2975
rect 16221 2941 16255 2975
rect 16255 2941 16264 2975
rect 16212 2932 16264 2941
rect 10784 2907 10836 2916
rect 10784 2873 10793 2907
rect 10793 2873 10827 2907
rect 10827 2873 10836 2907
rect 10784 2864 10836 2873
rect 12532 2907 12584 2916
rect 12532 2873 12541 2907
rect 12541 2873 12575 2907
rect 12575 2873 12584 2907
rect 12532 2864 12584 2873
rect 11612 2796 11664 2848
rect 11796 2839 11848 2848
rect 11796 2805 11805 2839
rect 11805 2805 11839 2839
rect 11839 2805 11848 2839
rect 11796 2796 11848 2805
rect 12440 2796 12492 2848
rect 15384 2839 15436 2848
rect 15384 2805 15393 2839
rect 15393 2805 15427 2839
rect 15427 2805 15436 2839
rect 18512 2864 18564 2916
rect 15384 2796 15436 2805
rect 16396 2796 16448 2848
rect 17500 2796 17552 2848
rect 17592 2796 17644 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 7104 2592 7156 2644
rect 7472 2592 7524 2644
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 10692 2524 10744 2576
rect 11428 2592 11480 2644
rect 12348 2635 12400 2644
rect 12348 2601 12357 2635
rect 12357 2601 12391 2635
rect 12391 2601 12400 2635
rect 12348 2592 12400 2601
rect 12624 2592 12676 2644
rect 12716 2592 12768 2644
rect 12900 2592 12952 2644
rect 13544 2592 13596 2644
rect 15292 2524 15344 2576
rect 16580 2592 16632 2644
rect 16948 2592 17000 2644
rect 17500 2592 17552 2644
rect 16212 2567 16264 2576
rect 16212 2533 16221 2567
rect 16221 2533 16255 2567
rect 16255 2533 16264 2567
rect 16212 2524 16264 2533
rect 17776 2524 17828 2576
rect 7472 2456 7524 2508
rect 10876 2456 10928 2508
rect 18328 2499 18380 2508
rect 10140 2388 10192 2440
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 11520 2320 11572 2372
rect 11612 2363 11664 2372
rect 11612 2329 11621 2363
rect 11621 2329 11655 2363
rect 11655 2329 11664 2363
rect 17592 2388 17644 2440
rect 11612 2320 11664 2329
rect 15660 2320 15712 2372
rect 7472 2295 7524 2304
rect 7472 2261 7481 2295
rect 7481 2261 7515 2295
rect 7515 2261 7524 2295
rect 7472 2252 7524 2261
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 19984 2320 20036 2372
rect 18420 2252 18472 2304
rect 19708 2252 19760 2304
rect 22652 2252 22704 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 938 27520 994 28000
rect 2778 27520 2834 28000
rect 4264 27526 4568 27554
rect 952 23798 980 27520
rect 1214 24304 1270 24313
rect 1214 24239 1270 24248
rect 940 23792 992 23798
rect 940 23734 992 23740
rect 1228 23186 1256 24239
rect 2792 23866 2820 27520
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2792 23662 2820 23802
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2504 23520 2556 23526
rect 2504 23462 2556 23468
rect 1216 23180 1268 23186
rect 1216 23122 1268 23128
rect 1228 22778 1256 23122
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 1216 22772 1268 22778
rect 1216 22714 1268 22720
rect 1950 19816 2006 19825
rect 1950 19751 2006 19760
rect 1964 18834 1992 19751
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1688 18222 1716 18566
rect 1964 18426 1992 18770
rect 2228 18692 2280 18698
rect 2228 18634 2280 18640
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1676 18216 1728 18222
rect 110 18184 166 18193
rect 1676 18158 1728 18164
rect 110 18119 166 18128
rect 124 18086 152 18119
rect 112 18080 164 18086
rect 112 18022 164 18028
rect 1688 17882 1716 18158
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 2240 17814 2268 18634
rect 2228 17808 2280 17814
rect 2228 17750 2280 17756
rect 2240 17338 2268 17750
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 1582 15464 1638 15473
rect 1582 15399 1638 15408
rect 1596 14618 1624 15399
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1412 14074 1440 14418
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1214 13696 1270 13705
rect 1214 13631 1270 13640
rect 1228 12850 1256 13631
rect 1216 12844 1268 12850
rect 1216 12786 1268 12792
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 1412 11218 1440 11494
rect 1582 11248 1638 11257
rect 1400 11212 1452 11218
rect 1582 11183 1638 11192
rect 1400 11154 1452 11160
rect 1412 10810 1440 11154
rect 1596 11082 1624 11183
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 2240 10713 2268 11494
rect 2226 10704 2282 10713
rect 2226 10639 2282 10648
rect 1582 9208 1638 9217
rect 1582 9143 1638 9152
rect 1596 8906 1624 9143
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1584 8900 1636 8906
rect 1584 8842 1636 8848
rect 1688 8838 1716 8978
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8634 1716 8774
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 2332 7993 2360 22918
rect 2516 18970 2544 23462
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 2516 18426 2544 18770
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 3252 18290 3280 18906
rect 3988 18902 4016 19314
rect 4264 18970 4292 27526
rect 4540 27418 4568 27526
rect 4618 27520 4674 28000
rect 6458 27520 6514 28000
rect 8390 27554 8446 28000
rect 8312 27526 8446 27554
rect 4632 27418 4660 27520
rect 4540 27390 4660 27418
rect 6274 26344 6330 26353
rect 6274 26279 6330 26288
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6288 24274 6316 26279
rect 6276 24268 6328 24274
rect 6276 24210 6328 24216
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6288 23866 6316 24210
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 4528 23520 4580 23526
rect 4528 23462 4580 23468
rect 4540 23118 4568 23462
rect 5540 23248 5592 23254
rect 5540 23190 5592 23196
rect 4528 23112 4580 23118
rect 4528 23054 4580 23060
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5460 22234 5488 23054
rect 5552 22642 5580 23190
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6288 22642 6316 23054
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 6276 22636 6328 22642
rect 6276 22578 6328 22584
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6288 20058 6316 22578
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6000 19984 6052 19990
rect 6000 19926 6052 19932
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4816 19378 4844 19790
rect 5448 19780 5500 19786
rect 5448 19722 5500 19728
rect 5460 19378 5488 19722
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6012 19514 6040 19926
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 3976 18896 4028 18902
rect 3976 18838 4028 18844
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4264 18358 4292 18770
rect 5460 18426 5488 19314
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 4252 18352 4304 18358
rect 4252 18294 4304 18300
rect 5552 18290 5580 18702
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 3884 18148 3936 18154
rect 3884 18090 3936 18096
rect 3344 17814 3372 18090
rect 2596 17808 2648 17814
rect 2596 17750 2648 17756
rect 3332 17808 3384 17814
rect 3332 17750 3384 17756
rect 2608 17270 2636 17750
rect 3896 17678 3924 18090
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3712 16454 3740 17070
rect 3896 16794 3924 17614
rect 4632 17338 4660 17682
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 5184 17270 5212 18158
rect 6104 18086 6132 18838
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6104 17814 6132 18022
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 6092 17808 6144 17814
rect 6092 17750 6144 17756
rect 5172 17264 5224 17270
rect 5172 17206 5224 17212
rect 5552 17066 5580 17750
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6012 17338 6040 17614
rect 6196 17542 6224 18158
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 4620 17060 4672 17066
rect 4620 17002 4672 17008
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3528 16046 3556 16390
rect 3712 16114 3740 16390
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15570 4568 15846
rect 4632 15638 4660 17002
rect 6012 16794 6040 17274
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 4816 16114 4844 16730
rect 6196 16658 6224 17478
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 5184 15910 5212 16186
rect 5552 16114 5580 16594
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 4620 15632 4672 15638
rect 4620 15574 4672 15580
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2976 15026 3004 15438
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 4540 14958 4568 15506
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4080 14618 4108 14826
rect 4632 14822 4660 15574
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 4080 12918 4108 13738
rect 4356 13462 4384 14214
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4344 13456 4396 13462
rect 4344 13398 4396 13404
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 12345 3096 12582
rect 4172 12442 4200 13262
rect 4356 12986 4384 13398
rect 4448 13326 4476 13874
rect 4632 13734 4660 14758
rect 5092 14618 5120 14826
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 5000 13802 5028 14418
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4632 12714 4660 13670
rect 5000 12986 5028 13738
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4632 12374 4660 12650
rect 4620 12368 4672 12374
rect 3054 12336 3110 12345
rect 4620 12310 4672 12316
rect 3054 12271 3110 12280
rect 4724 11558 4752 12718
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 5184 11218 5212 15846
rect 5276 15026 5304 16050
rect 5552 15910 5580 16050
rect 6196 15910 6224 16594
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5552 15434 5580 15642
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 10810 5212 11154
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2608 8294 2636 8978
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2318 7984 2374 7993
rect 2318 7919 2374 7928
rect 2608 7857 2636 8230
rect 2594 7848 2650 7857
rect 2594 7783 2650 7792
rect 110 7440 166 7449
rect 110 7375 166 7384
rect 124 7342 152 7375
rect 112 7336 164 7342
rect 112 7278 164 7284
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 1582 4720 1638 4729
rect 1582 4655 1584 4664
rect 1636 4655 1638 4664
rect 1584 4626 1636 4632
rect 1596 4282 1624 4626
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 572 3936 624 3942
rect 572 3878 624 3884
rect 110 3088 166 3097
rect 166 3058 244 3074
rect 166 3052 256 3058
rect 166 3046 204 3052
rect 110 3023 166 3032
rect 204 2994 256 3000
rect 584 82 612 3878
rect 2318 2000 2374 2009
rect 2318 1935 2374 1944
rect 662 82 718 480
rect 584 54 718 82
rect 662 0 718 54
rect 2042 82 2098 480
rect 2332 82 2360 1935
rect 2042 54 2360 82
rect 3422 82 3478 480
rect 3804 82 3832 4150
rect 3422 54 3832 82
rect 4802 82 4858 480
rect 5092 82 5120 7278
rect 5276 3602 5304 14962
rect 5552 14618 5580 15370
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6012 14074 6040 14418
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5460 11354 5488 12174
rect 5552 11898 5580 12310
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6196 11898 6224 15846
rect 6380 15026 6408 24006
rect 6472 23866 6500 27520
rect 8312 24274 8340 27526
rect 8390 27520 8446 27526
rect 10230 27520 10286 28000
rect 12070 27520 12126 28000
rect 13910 27520 13966 28000
rect 15842 27520 15898 28000
rect 17682 27520 17738 28000
rect 19522 27520 19578 28000
rect 21362 27520 21418 28000
rect 23294 27520 23350 28000
rect 23756 27532 23808 27538
rect 10244 25786 10272 27520
rect 10152 25758 10272 25786
rect 10152 24274 10180 25758
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 7564 24268 7616 24274
rect 7564 24210 7616 24216
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 10140 24268 10192 24274
rect 10140 24210 10192 24216
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6460 23860 6512 23866
rect 6460 23802 6512 23808
rect 6840 23662 6868 24006
rect 6828 23656 6880 23662
rect 6828 23598 6880 23604
rect 6840 23322 6868 23598
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 7576 23050 7604 24210
rect 8312 23866 8340 24210
rect 8668 24064 8720 24070
rect 8668 24006 8720 24012
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 8680 23730 8708 24006
rect 8668 23724 8720 23730
rect 8668 23666 8720 23672
rect 9128 23588 9180 23594
rect 9128 23530 9180 23536
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 8116 23248 8168 23254
rect 8036 23208 8116 23236
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 6920 22500 6972 22506
rect 6920 22442 6972 22448
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6472 19310 6500 19450
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6472 18970 6500 19246
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6564 17882 6592 22374
rect 6932 22234 6960 22442
rect 7852 22234 7880 23054
rect 8036 22438 8064 23208
rect 8116 23190 8168 23196
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8772 22642 8800 23054
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 6932 22137 6960 22170
rect 8036 22166 8064 22374
rect 8024 22160 8076 22166
rect 6918 22128 6974 22137
rect 8024 22102 8076 22108
rect 6918 22063 6974 22072
rect 7286 21992 7342 22001
rect 7286 21927 7342 21936
rect 7300 21010 7328 21927
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 7300 20602 7328 20946
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 7288 20596 7340 20602
rect 7288 20538 7340 20544
rect 8588 20466 8616 20742
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8668 20324 8720 20330
rect 8668 20266 8720 20272
rect 8116 19984 8168 19990
rect 8116 19926 8168 19932
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 6552 17876 6604 17882
rect 6552 17818 6604 17824
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6656 15570 6684 17206
rect 6840 16998 6868 17478
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6656 15162 6684 15506
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6472 13841 6500 15098
rect 6458 13832 6514 13841
rect 6380 13786 6458 13814
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6288 12986 6316 13330
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6288 12714 6316 12922
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 6288 12442 6316 12650
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6380 11762 6408 13786
rect 6458 13767 6514 13776
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6748 12374 6776 13262
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5552 11218 5580 11630
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 10810 5580 11154
rect 6472 11014 6500 12174
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6196 9178 6224 9658
rect 6288 9654 6316 9930
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6104 8294 6132 8978
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6104 7886 6132 8230
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6288 7274 6316 7890
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6288 6866 6316 7210
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6196 6118 6224 6802
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5778 6224 6054
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6196 5030 6224 5714
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 3194 6040 3538
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6196 1601 6224 4966
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6288 4078 6316 4626
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6288 3942 6316 4014
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6472 3194 6500 10950
rect 6564 10062 6592 11290
rect 6840 10266 6868 16934
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6932 15570 6960 16118
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6932 14822 6960 15506
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 7208 13462 7236 15846
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7300 14550 7328 14962
rect 7288 14544 7340 14550
rect 7288 14486 7340 14492
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6932 12753 6960 12786
rect 6918 12744 6974 12753
rect 6918 12679 6974 12688
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 12186 7328 12582
rect 7116 12158 7328 12186
rect 7116 11830 7144 12158
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7208 11626 7236 12038
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7208 11286 7236 11562
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7208 10742 7236 11222
rect 7300 11014 7328 12158
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6564 9518 6592 9998
rect 6656 9654 6684 10066
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6564 8362 6592 8774
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6564 7342 6592 7822
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6656 7478 6684 7686
rect 6840 7546 6868 7686
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6656 5778 6684 6122
rect 6932 5914 6960 10406
rect 7208 10198 7236 10678
rect 7300 10470 7328 10950
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7116 9518 7144 9998
rect 7208 9654 7236 10134
rect 7300 10130 7328 10406
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7024 8634 7052 8978
rect 7116 8974 7144 9454
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 9178 7236 9386
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7208 8090 7236 8366
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 7024 7206 7052 7754
rect 7208 7342 7236 8026
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7024 6934 7052 7142
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7024 6186 7052 6870
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7116 6254 7144 6734
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6644 5772 6696 5778
rect 6564 5732 6644 5760
rect 6564 5030 6592 5732
rect 6644 5714 6696 5720
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6182 1592 6238 1601
rect 6182 1527 6238 1536
rect 4802 54 5120 82
rect 6182 82 6238 480
rect 6564 82 6592 4966
rect 6748 4690 6776 5102
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6840 4826 6868 5034
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6748 4214 6776 4626
rect 6840 4282 6868 4762
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 7392 4154 7420 13738
rect 7116 4126 7420 4154
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6840 3738 6868 4014
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 7116 2650 7144 4126
rect 7484 2650 7512 19654
rect 8128 19514 8156 19926
rect 8680 19786 8708 20266
rect 8668 19780 8720 19786
rect 8668 19722 8720 19728
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7576 18086 7604 18770
rect 8036 18290 8064 18906
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7576 16114 7604 18022
rect 7760 17066 7788 18022
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8036 17270 8064 17682
rect 8220 17678 8248 18770
rect 8588 18154 8616 19110
rect 8680 18426 8708 19722
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8772 18630 8800 19246
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8772 17814 8800 18566
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 7760 16726 7788 17002
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7760 16250 7788 16662
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7668 14890 7696 15302
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7668 14618 7696 14826
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7760 14550 7788 16186
rect 7944 15910 7972 16390
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 8220 15706 8248 17070
rect 8864 16794 8892 23462
rect 9140 23050 9168 23530
rect 9968 23254 9996 23530
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 9956 23248 10008 23254
rect 9956 23190 10008 23196
rect 9128 23044 9180 23050
rect 9128 22986 9180 22992
rect 9140 22710 9168 22986
rect 9784 22778 9812 23190
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 8944 22500 8996 22506
rect 8944 22442 8996 22448
rect 8956 22098 8984 22442
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8956 21894 8984 22034
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8956 21350 8984 21830
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 8956 17338 8984 21286
rect 9692 20602 9720 21286
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9968 20602 9996 20742
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 9220 20324 9272 20330
rect 9220 20266 9272 20272
rect 9232 19854 9260 20266
rect 9968 20262 9996 20538
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 10060 18612 10088 24006
rect 10152 23866 10180 24210
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10152 22778 10180 23054
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 11256 21690 11284 22510
rect 12084 22098 12112 27520
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 11428 22092 11480 22098
rect 11428 22034 11480 22040
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 11440 21690 11468 22034
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 10784 21480 10836 21486
rect 10784 21422 10836 21428
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10336 20602 10364 20946
rect 10324 20596 10376 20602
rect 10152 20556 10324 20584
rect 10152 19990 10180 20556
rect 10324 20538 10376 20544
rect 10796 20466 10824 21422
rect 11900 21078 11928 21830
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 11888 21072 11940 21078
rect 11888 21014 11940 21020
rect 12164 21072 12216 21078
rect 12164 21014 12216 21020
rect 11900 20602 11928 21014
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10796 19990 10824 20402
rect 12176 20262 12204 21014
rect 12452 20874 12480 21558
rect 12544 21554 12572 21830
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12624 21412 12676 21418
rect 12624 21354 12676 21360
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 10140 19984 10192 19990
rect 10140 19926 10192 19932
rect 10784 19984 10836 19990
rect 10784 19926 10836 19932
rect 10152 19514 10180 19926
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10244 19514 10272 19790
rect 11348 19786 11376 19858
rect 11336 19780 11388 19786
rect 11336 19722 11388 19728
rect 11348 19514 11376 19722
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 12176 18970 12204 20198
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 9784 18584 10088 18612
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8404 15570 8432 15982
rect 9416 15910 9444 16594
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9048 15570 9076 15846
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 8220 15162 8248 15506
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7668 13802 7696 14418
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7852 14006 7880 14350
rect 8128 14006 8156 15030
rect 8220 14074 8248 15098
rect 8864 14822 8892 15506
rect 8668 14816 8720 14822
rect 8852 14816 8904 14822
rect 8720 14776 8800 14804
rect 8668 14758 8720 14764
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7668 13530 7696 13738
rect 7852 13530 7880 13942
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 8404 13394 8432 14214
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8404 12986 8432 13330
rect 8772 12986 8800 14776
rect 8852 14758 8904 14764
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7576 12238 7604 12786
rect 8220 12646 8248 12854
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7760 11898 7788 12310
rect 8220 12102 8248 12582
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 8220 11830 8248 12038
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 11150 7880 11698
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7852 10810 7880 11086
rect 8220 11014 8248 11766
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7852 9722 7880 10746
rect 8220 10470 8248 10950
rect 8312 10538 8340 11222
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10130 8248 10406
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8116 10056 8168 10062
rect 7944 10016 8116 10044
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7576 8634 7604 8842
rect 7852 8634 7880 9658
rect 7944 9382 7972 10016
rect 8116 9998 8168 10004
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8128 9654 8156 9862
rect 8220 9654 8248 10066
rect 8404 9722 8432 12922
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8588 11898 8616 12038
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8588 11014 8616 11630
rect 8772 11354 8800 12786
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8496 10606 8524 10950
rect 8588 10810 8616 10950
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8496 9722 8524 10542
rect 8588 10266 8616 10746
rect 8772 10674 8800 11290
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8772 10010 8800 10610
rect 8864 10198 8892 14758
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8956 12714 8984 13126
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8956 11626 8984 12650
rect 9048 11898 9076 15506
rect 9416 14822 9444 15846
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9312 13864 9364 13870
rect 9416 13841 9444 14758
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 13870 9536 14214
rect 9496 13864 9548 13870
rect 9312 13806 9364 13812
rect 9402 13832 9458 13841
rect 9324 13258 9352 13806
rect 9496 13806 9548 13812
rect 9402 13767 9458 13776
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8956 11082 8984 11562
rect 9324 11354 9352 13194
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9600 11218 9628 14758
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9692 11898 9720 12242
rect 9784 12238 9812 18584
rect 10796 18086 10824 18702
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11440 18222 11468 18566
rect 11428 18216 11480 18222
rect 11428 18158 11480 18164
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10520 17542 10548 17750
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17202 10548 17478
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16114 10180 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10244 16046 10272 16594
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 10060 14550 10088 15030
rect 10336 15026 10364 15302
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 13802 9904 14350
rect 10060 14074 10088 14486
rect 10600 14272 10652 14278
rect 10704 14260 10732 14826
rect 10652 14232 10732 14260
rect 10600 14214 10652 14220
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 9954 13832 10010 13841
rect 9864 13796 9916 13802
rect 10060 13814 10088 14010
rect 10612 13870 10640 14214
rect 10600 13864 10652 13870
rect 10060 13786 10180 13814
rect 10600 13806 10652 13812
rect 9954 13767 10010 13776
rect 9864 13738 9916 13744
rect 9876 13530 9904 13738
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9968 12306 9996 13767
rect 10152 12986 10180 13786
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12374 10732 12718
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 9784 11898 9812 12038
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 10704 11830 10732 12038
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 10152 11354 10180 11630
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 9600 10810 9628 11154
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8772 9982 8892 10010
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8208 9648 8260 9654
rect 8260 9608 8340 9636
rect 8208 9590 8260 9596
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 8956 7972 9318
rect 8036 9110 8064 9454
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8024 8968 8076 8974
rect 7944 8928 8024 8956
rect 8024 8910 8076 8916
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7576 7750 7604 8298
rect 8036 8294 8064 8910
rect 8128 8838 8156 9590
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8128 8430 8156 8774
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8220 8362 8248 8978
rect 8312 8634 8340 9608
rect 8772 9518 8800 9862
rect 8864 9586 8892 9982
rect 9140 9654 9168 10202
rect 9416 10198 9444 10406
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9692 10130 9720 11222
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 9784 10470 9812 11018
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8484 8424 8536 8430
rect 8404 8384 8484 8412
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8036 7954 8064 8230
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 6118 7604 7686
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7944 7002 7972 7278
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7668 5914 7696 6802
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8036 6458 8064 6734
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 8036 5846 8064 6190
rect 8220 6118 8248 8298
rect 8404 7342 8432 8384
rect 8484 8366 8536 8372
rect 8772 8090 8800 9454
rect 9140 8906 9168 9590
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9416 9178 9444 9522
rect 9692 9518 9720 10066
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9784 9450 9812 10406
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9784 9178 9812 9386
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9140 8498 9168 8842
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8496 7342 8524 7822
rect 8392 7336 8444 7342
rect 8312 7296 8392 7324
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7760 4826 7788 5646
rect 8036 5234 8064 5782
rect 8128 5642 8156 6054
rect 8312 5642 8340 7296
rect 8392 7278 8444 7284
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8404 6730 8432 6938
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8404 6390 8432 6666
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8496 6322 8524 7278
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8036 4826 8064 5170
rect 8128 5166 8156 5578
rect 8312 5370 8340 5578
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8128 4282 8156 5102
rect 8312 4758 8340 5306
rect 8404 5098 8432 6054
rect 8496 5914 8524 6258
rect 8772 6254 8800 8026
rect 8956 7721 8984 8298
rect 8942 7712 8998 7721
rect 8942 7647 8998 7656
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8956 7313 8984 7346
rect 8942 7304 8998 7313
rect 8942 7239 8998 7248
rect 9416 7206 9444 9114
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 7546 9720 7890
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 9416 5778 9444 7142
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6458 9536 6598
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9508 5914 9536 6394
rect 9692 6118 9720 6802
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9876 5778 9904 9998
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10060 9178 10088 9590
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10060 6798 10088 7278
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 9968 6322 9996 6666
rect 10060 6458 10088 6734
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9048 5166 9076 5510
rect 9416 5370 9444 5714
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9784 5545 9812 5646
rect 9770 5536 9826 5545
rect 9770 5471 9826 5480
rect 9876 5370 9904 5714
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9968 5250 9996 5782
rect 9876 5222 9996 5250
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8312 4214 8340 4694
rect 8404 4622 8432 5034
rect 9140 4826 9168 5034
rect 9876 5030 9904 5222
rect 10152 5148 10180 11018
rect 10796 10470 10824 18022
rect 11440 17882 11468 18158
rect 11716 18086 11744 18838
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11716 17814 11744 18022
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10888 16726 10916 17614
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11440 16726 11468 17206
rect 10876 16720 10928 16726
rect 11428 16720 11480 16726
rect 10876 16662 10928 16668
rect 11348 16680 11428 16708
rect 11348 16250 11376 16680
rect 11428 16662 11480 16668
rect 12452 16674 12480 20810
rect 12636 20602 12664 21354
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12544 17882 12572 18226
rect 12636 17882 12664 18294
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12544 17105 12572 17138
rect 12530 17096 12586 17105
rect 12530 17031 12586 17040
rect 12544 16794 12572 17031
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12452 16646 12572 16674
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 11626 10916 12242
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10888 10130 10916 11562
rect 10980 11286 11008 16118
rect 11440 15910 11468 16526
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11348 14414 11376 15438
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 14074 11376 14350
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 11072 12646 11100 13330
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10888 9722 10916 10066
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 11164 9042 11192 10542
rect 11256 10130 11284 11086
rect 11440 11082 11468 15846
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11808 14822 11836 15506
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11624 13938 11652 14486
rect 11808 14414 11836 14758
rect 12452 14618 12480 15302
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 12452 13870 12480 14554
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11900 12986 11928 13398
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 12084 12442 12112 13262
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12268 12714 12296 13126
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12176 11898 12204 12650
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12176 11626 12204 11834
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11256 9722 11284 10066
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 10612 8634 10640 8978
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10704 7546 10732 7890
rect 10888 7750 10916 8366
rect 11164 8090 11192 8978
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10704 7342 10732 7482
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10888 6662 10916 7686
rect 11256 7342 11284 8366
rect 11348 7886 11376 9318
rect 11440 8566 11468 10542
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11532 8498 11560 11494
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11900 10810 11928 11018
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11808 10577 11836 10610
rect 11900 10606 11928 10746
rect 11888 10600 11940 10606
rect 11794 10568 11850 10577
rect 11888 10542 11940 10548
rect 11794 10503 11850 10512
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11624 9042 11652 9998
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11624 7954 11652 8978
rect 11900 8294 11928 9046
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11256 7002 11284 7278
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11532 6798 11560 7210
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10888 6390 10916 6598
rect 11532 6458 11560 6734
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10980 5574 11008 6190
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10704 5234 10732 5510
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10060 5120 10180 5148
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9876 4758 9904 4966
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 9968 4486 9996 4966
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 9968 4146 9996 4422
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9956 3188 10008 3194
rect 10060 3176 10088 5120
rect 10232 5092 10284 5098
rect 10152 5052 10232 5080
rect 10152 4536 10180 5052
rect 10232 5034 10284 5040
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10232 4548 10284 4554
rect 10152 4508 10232 4536
rect 10232 4490 10284 4496
rect 10244 4282 10272 4490
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10152 3641 10180 4150
rect 10704 4078 10732 5170
rect 10980 4826 11008 5510
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 11072 4690 11100 6054
rect 11624 5914 11652 7890
rect 11900 6934 11928 8230
rect 11992 8022 12020 8298
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11992 7546 12020 7958
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7546 12204 7822
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 11900 6118 11928 6870
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10138 3632 10194 3641
rect 10138 3567 10194 3576
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10008 3148 10088 3176
rect 9956 3130 10008 3136
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7484 2310 7512 2450
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 6182 54 6592 82
rect 7484 82 7512 2246
rect 7654 82 7710 480
rect 7484 54 7710 82
rect 8680 82 8708 2790
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2582 10732 3470
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10796 2650 10824 2858
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 10888 2514 10916 4150
rect 11072 3738 11100 4626
rect 11256 4078 11284 4762
rect 11624 4282 11652 5850
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11808 5234 11836 5782
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11796 4752 11848 4758
rect 11900 4740 11928 6054
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12164 5704 12216 5710
rect 12268 5692 12296 12650
rect 12452 9178 12480 13126
rect 12544 10266 12572 16646
rect 12820 15162 12848 23598
rect 13544 22092 13596 22098
rect 13544 22034 13596 22040
rect 13556 22001 13584 22034
rect 13542 21992 13598 22001
rect 13542 21927 13598 21936
rect 13556 21690 13584 21927
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 13924 20058 13952 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15856 23866 15884 27520
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 17696 22778 17724 27520
rect 18604 23656 18656 23662
rect 18602 23624 18604 23633
rect 18656 23624 18658 23633
rect 18602 23559 18658 23568
rect 18616 23526 18644 23559
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 17684 22772 17736 22778
rect 17684 22714 17736 22720
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14646 20496 14702 20505
rect 14646 20431 14702 20440
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12912 19446 12940 19858
rect 14660 19514 14688 20431
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 12900 19440 12952 19446
rect 12900 19382 12952 19388
rect 14660 19310 14688 19450
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 14096 19168 14148 19174
rect 14096 19110 14148 19116
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 13004 18290 13032 18702
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13188 18154 13216 19110
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 13188 17678 13216 18090
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 12912 17202 12940 17614
rect 13464 17338 13492 17750
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12912 16658 12940 17138
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13740 16250 13768 16526
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13924 15910 13952 16662
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15706 13952 15846
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13740 15162 13768 15506
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 12622 13832 12678 13841
rect 12622 13767 12678 13776
rect 12636 13734 12664 13767
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12728 13462 12756 14894
rect 13832 14618 13860 14894
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13096 13734 13124 14418
rect 13832 13938 13860 14418
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12728 12850 12756 13398
rect 13096 13258 13124 13670
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 13188 13190 13216 13874
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13556 13530 13584 13806
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13648 12986 13676 13330
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12986 13860 13126
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12636 12442 12664 12650
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 13648 12374 13676 12922
rect 13832 12646 13860 12922
rect 14108 12850 14136 19110
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14384 16998 14412 17682
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 17512 17105 17540 18022
rect 17498 17096 17554 17105
rect 17498 17031 17554 17040
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 14384 16726 14412 16934
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14384 16114 14412 16662
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14464 15972 14516 15978
rect 14464 15914 14516 15920
rect 14476 15706 14504 15914
rect 14752 15910 14780 16390
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 17236 16250 17264 16526
rect 17512 16522 17540 16934
rect 17592 16720 17644 16726
rect 17592 16662 17644 16668
rect 17500 16516 17552 16522
rect 17500 16458 17552 16464
rect 17604 16250 17632 16662
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 15106 16008 15162 16017
rect 15106 15943 15162 15952
rect 15120 15910 15148 15943
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15856 15026 15884 15438
rect 16132 15094 16160 15574
rect 17788 15502 17816 23462
rect 18708 23118 18736 23462
rect 18696 23112 18748 23118
rect 18696 23054 18748 23060
rect 19536 18426 19564 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 21376 23866 21404 27520
rect 23308 23866 23336 27520
rect 25134 27532 25190 28000
rect 25134 27520 25136 27532
rect 23756 27474 23808 27480
rect 25188 27520 25190 27532
rect 26974 27520 27030 28000
rect 25136 27474 25188 27480
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 21732 23588 21784 23594
rect 21732 23530 21784 23536
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18340 17882 18368 18158
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18052 17060 18104 17066
rect 18052 17002 18104 17008
rect 18064 16726 18092 17002
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 18248 16454 18276 16934
rect 18432 16522 18460 17682
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 18420 16516 18472 16522
rect 18420 16458 18472 16464
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 18248 15978 18276 16390
rect 18432 16114 18460 16458
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18236 15972 18288 15978
rect 18236 15914 18288 15920
rect 18248 15706 18276 15914
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18708 15638 18736 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 18144 15632 18196 15638
rect 18144 15574 18196 15580
rect 18696 15632 18748 15638
rect 18696 15574 18748 15580
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17788 15162 17816 15438
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15488 13870 15516 14214
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14384 13394 14412 13738
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14372 13388 14424 13394
rect 14424 13348 14504 13376
rect 14372 13330 14424 13336
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 14108 12442 14136 12786
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 13636 12368 13688 12374
rect 12990 12336 13046 12345
rect 13636 12310 13688 12316
rect 12990 12271 13046 12280
rect 13004 12238 13032 12271
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12728 10470 12756 11154
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12544 9586 12572 10202
rect 12728 9926 12756 10406
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12636 8838 12664 9386
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8430 12664 8774
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12636 8090 12664 8366
rect 12728 8294 12756 9862
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12820 7954 12848 9522
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12544 7857 12572 7890
rect 12530 7848 12586 7857
rect 12530 7783 12586 7792
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12728 5710 12756 6122
rect 12216 5664 12296 5692
rect 12716 5704 12768 5710
rect 12164 5646 12216 5652
rect 12716 5646 12768 5652
rect 12084 5234 12112 5646
rect 12176 5302 12204 5646
rect 12728 5370 12756 5646
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12164 5296 12216 5302
rect 12164 5238 12216 5244
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12084 5137 12112 5170
rect 12070 5128 12126 5137
rect 12070 5063 12126 5072
rect 11848 4712 11928 4740
rect 11796 4694 11848 4700
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11808 4146 11836 4694
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11440 3534 11468 3946
rect 11808 3942 11836 4082
rect 11992 4078 12020 4422
rect 12912 4154 12940 12106
rect 13004 11354 13032 12174
rect 13648 11898 13676 12310
rect 14384 12170 14412 12786
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 14372 12164 14424 12170
rect 14372 12106 14424 12112
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 10130 13492 10542
rect 13648 10538 13676 10950
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13648 10130 13676 10474
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13464 9722 13492 10066
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13648 9110 13676 10066
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13464 8634 13492 8910
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13372 6458 13400 7822
rect 13464 7546 13492 7890
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13464 7206 13492 7482
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13464 7002 13492 7142
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13372 6118 13400 6394
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 6186 13584 6258
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13004 5846 13032 6054
rect 13556 5914 13584 6122
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 12992 5840 13044 5846
rect 13648 5828 13676 8230
rect 13740 7410 13768 12106
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14292 11694 14320 12038
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 9178 13860 11494
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14108 10606 14136 11018
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14292 10266 14320 11630
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14016 9722 14044 10066
rect 14476 9722 14504 13348
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14568 11286 14596 11494
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14844 10130 14872 13670
rect 15580 13530 15608 14758
rect 15856 13870 15884 14962
rect 16132 14872 16160 15030
rect 16212 14884 16264 14890
rect 16132 14844 16212 14872
rect 16132 14618 16160 14844
rect 16212 14826 16264 14832
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16500 13938 16528 14350
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15672 13394 15700 13806
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12986 15332 13330
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15672 12646 15700 13330
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15396 11898 15424 12242
rect 15384 11892 15436 11898
rect 15436 11852 15516 11880
rect 15384 11834 15436 11840
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 11354 15424 11494
rect 15488 11354 15516 11852
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15488 10538 15516 11290
rect 15672 10577 15700 12582
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15764 11898 15792 12038
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15764 11558 15792 11834
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15764 10810 15792 11086
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 16040 10713 16068 11698
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16026 10704 16082 10713
rect 16026 10639 16082 10648
rect 16040 10606 16068 10639
rect 16028 10600 16080 10606
rect 15658 10568 15714 10577
rect 15476 10532 15528 10538
rect 16028 10542 16080 10548
rect 15658 10503 15714 10512
rect 15476 10474 15528 10480
rect 16316 10470 16344 11222
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15672 9722 15700 10066
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 14476 9518 14504 9658
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 14476 9042 14504 9454
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14476 8634 14504 8978
rect 15120 8906 15148 9454
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14660 7721 14688 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15488 8022 15516 8978
rect 15672 8634 15700 9658
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15764 9042 15792 9590
rect 15856 9518 15884 10066
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16132 9586 16160 9998
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 16132 9178 16160 9522
rect 16316 9450 16344 10406
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16224 9042 16252 9386
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15764 8430 15792 8978
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15764 8090 15792 8366
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 16040 7954 16068 8910
rect 16396 8016 16448 8022
rect 16316 7976 16396 8004
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 14646 7712 14702 7721
rect 14646 7647 14702 7656
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 16040 7546 16068 7890
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 13740 7002 13768 7346
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14016 6322 14044 6734
rect 14108 6390 14136 7346
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 13728 5840 13780 5846
rect 13648 5800 13728 5828
rect 12992 5782 13044 5788
rect 13728 5782 13780 5788
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 13096 5370 13124 5714
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 12912 4126 13124 4154
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 11808 3738 11836 3878
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 9034 82 9090 480
rect 8680 54 9090 82
rect 10152 82 10180 2382
rect 10980 1873 11008 3334
rect 11440 2650 11468 3470
rect 11808 2854 11836 3674
rect 12176 3194 12204 3878
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12360 2990 12388 3334
rect 12452 3194 12480 3946
rect 13096 3670 13124 4126
rect 13280 3942 13308 4626
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13464 3670 13492 4014
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11624 2378 11652 2790
rect 11520 2372 11572 2378
rect 11520 2314 11572 2320
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 10966 1864 11022 1873
rect 10966 1799 11022 1808
rect 10414 82 10470 480
rect 10152 54 10470 82
rect 11532 82 11560 2314
rect 11808 2009 11836 2790
rect 12360 2650 12388 2926
rect 12452 2854 12480 3130
rect 12544 2922 12572 3334
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 11794 2000 11850 2009
rect 11794 1935 11850 1944
rect 12544 1737 12572 2858
rect 12624 2644 12676 2650
rect 12716 2644 12768 2650
rect 12676 2604 12716 2632
rect 12624 2586 12676 2592
rect 12716 2586 12768 2592
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 12716 2440 12768 2446
rect 12912 2428 12940 2586
rect 12768 2400 12940 2428
rect 12716 2382 12768 2388
rect 12530 1728 12586 1737
rect 12530 1663 12586 1672
rect 11794 82 11850 480
rect 11532 54 11850 82
rect 13096 82 13124 3062
rect 13280 2990 13308 3606
rect 13464 3194 13492 3606
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13556 3058 13584 3470
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13556 2650 13584 2994
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 13174 82 13230 480
rect 13740 105 13768 5782
rect 14660 5778 14688 7210
rect 14844 7206 14872 7278
rect 16316 7206 16344 7976
rect 16396 7958 16448 7964
rect 16592 7313 16620 14826
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 17052 14618 17080 14758
rect 18156 14618 18184 15574
rect 18708 15094 18736 15574
rect 18696 15088 18748 15094
rect 18696 15030 18748 15036
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18248 14550 18276 14826
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 16672 14544 16724 14550
rect 16672 14486 16724 14492
rect 18236 14544 18288 14550
rect 18236 14486 18288 14492
rect 16684 14074 16712 14486
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 17512 13433 17540 14214
rect 18432 14074 18460 14418
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 17498 13424 17554 13433
rect 17498 13359 17554 13368
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19996 12442 20024 23462
rect 21744 22137 21772 23530
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 21730 22128 21786 22137
rect 21730 22063 21786 22072
rect 22204 12753 22232 22918
rect 23768 18222 23796 27474
rect 25148 27443 25176 27474
rect 25134 26480 25190 26489
rect 25134 26415 25190 26424
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24674 24440 24730 24449
rect 24674 24375 24730 24384
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23186 24716 24375
rect 25148 23866 25176 26415
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25148 23662 25176 23802
rect 25136 23656 25188 23662
rect 26988 23633 27016 27520
rect 25136 23598 25188 23604
rect 26974 23624 27030 23633
rect 26974 23559 27030 23568
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22778 24716 23122
rect 27618 22944 27674 22953
rect 27618 22879 27674 22888
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 27632 22001 27660 22879
rect 27618 21992 27674 22001
rect 27618 21927 27674 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24674 18456 24730 18465
rect 24674 18391 24730 18400
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 24688 17746 24716 18391
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22190 12744 22246 12753
rect 22190 12679 22246 12688
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 18156 11762 18184 12378
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17788 11354 17816 11494
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17604 10810 17632 11154
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17604 10198 17632 10746
rect 18432 10674 18460 11698
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18432 10198 18460 10610
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16776 8634 16804 8978
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16578 7304 16634 7313
rect 16578 7239 16634 7248
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 14844 6458 14872 7142
rect 15396 7002 15424 7142
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14094 5536 14150 5545
rect 14094 5471 14150 5480
rect 14108 5166 14136 5471
rect 14844 5302 14872 6394
rect 15396 6322 15424 6938
rect 16316 6934 16344 7142
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 16316 6186 16344 6870
rect 16684 6866 16712 8298
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16684 6458 16712 6802
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16304 6180 16356 6186
rect 16304 6122 16356 6128
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15488 5846 15516 6054
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15488 5370 15516 5782
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16592 5370 16620 5646
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 14832 5296 14884 5302
rect 14832 5238 14884 5244
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14108 4826 14136 5102
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14384 4060 14412 5034
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15304 4690 15332 4966
rect 15488 4758 15516 5306
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 14556 4548 14608 4554
rect 14556 4490 14608 4496
rect 14464 4072 14516 4078
rect 14384 4032 14464 4060
rect 14464 4014 14516 4020
rect 14476 3738 14504 4014
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 13096 54 13230 82
rect 2042 0 2098 54
rect 3422 0 3478 54
rect 4802 0 4858 54
rect 6182 0 6238 54
rect 7654 0 7710 54
rect 9034 0 9090 54
rect 10414 0 10470 54
rect 11794 0 11850 54
rect 13174 0 13230 54
rect 13726 96 13782 105
rect 14568 82 14596 4490
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 3738 15332 4626
rect 15488 4010 15516 4694
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16500 4078 16528 4422
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15304 2582 15332 3470
rect 15396 2854 15424 3878
rect 16500 3670 16528 4014
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 16224 2582 16252 2926
rect 16408 2854 16436 3470
rect 16500 3194 16528 3606
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16592 2650 16620 3470
rect 16684 3058 16712 3606
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16960 2650 16988 9862
rect 17604 9722 17632 10134
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 17420 9110 17448 9386
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 17420 8634 17448 9046
rect 18064 8634 18092 9386
rect 19076 9110 19104 9454
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18064 8344 18092 8570
rect 18156 8498 18184 8774
rect 18800 8498 18828 8910
rect 19076 8634 19104 9046
rect 19536 8634 19564 9114
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18144 8356 18196 8362
rect 18064 8316 18144 8344
rect 18144 8298 18196 8304
rect 17406 7984 17462 7993
rect 17406 7919 17462 7928
rect 18236 7948 18288 7954
rect 17420 7546 17448 7919
rect 18236 7890 18288 7896
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 17236 4010 17264 4694
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 17604 3058 17632 6258
rect 17788 4622 17816 7754
rect 18248 7274 18276 7890
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18236 7268 18288 7274
rect 18236 7210 18288 7216
rect 18248 7002 18276 7210
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18248 5166 18276 6802
rect 18340 5846 18368 7686
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18524 6934 18552 7346
rect 18512 6928 18564 6934
rect 18512 6870 18564 6876
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 18340 5302 18368 5782
rect 18432 5370 18460 6054
rect 18524 5710 18552 6870
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 18248 4826 18276 5102
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18616 4690 18644 5510
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 17776 4616 17828 4622
rect 18616 4593 18644 4626
rect 17776 4558 17828 4564
rect 18602 4584 18658 4593
rect 17684 4548 17736 4554
rect 17684 4490 17736 4496
rect 17696 3670 17724 4490
rect 17788 4214 17816 4558
rect 18602 4519 18658 4528
rect 18800 4282 18828 8434
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 22296 7818 22324 17478
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17338 24716 17682
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 25134 16416 25190 16425
rect 24289 16348 24585 16368
rect 25134 16351 25190 16360
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 25148 16250 25176 16351
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25148 16046 25176 16186
rect 25136 16040 25188 16046
rect 24858 16008 24914 16017
rect 25136 15982 25188 15988
rect 24858 15943 24914 15952
rect 24872 15638 24900 15943
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 24216 15632 24268 15638
rect 24216 15574 24268 15580
rect 24860 15632 24912 15638
rect 24860 15574 24912 15580
rect 24228 15026 24256 15574
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 24044 14532 24072 14894
rect 24872 14550 24900 15574
rect 25056 15502 25084 15846
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 25056 15162 25084 15438
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 27618 15056 27674 15065
rect 27618 14991 27674 15000
rect 24124 14544 24176 14550
rect 24044 14504 24124 14532
rect 24044 13734 24072 14504
rect 24124 14486 24176 14492
rect 24860 14544 24912 14550
rect 24860 14486 24912 14492
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24872 13734 24900 14350
rect 27632 13841 27660 14991
rect 27618 13832 27674 13841
rect 27618 13767 27674 13776
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 24860 13728 24912 13734
rect 24860 13670 24912 13676
rect 24044 13433 24072 13670
rect 24030 13424 24086 13433
rect 24030 13359 24086 13368
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24674 12472 24730 12481
rect 24674 12407 24730 12416
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11218 24716 12407
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 23940 11008 23992 11014
rect 23940 10950 23992 10956
rect 22926 10432 22982 10441
rect 22926 10367 22982 10376
rect 22940 9042 22968 10367
rect 23952 10266 23980 10950
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10810 24716 11154
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23940 10260 23992 10266
rect 23940 10202 23992 10208
rect 23400 9586 23428 10202
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 24584 9444 24636 9450
rect 24584 9386 24636 9392
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 22928 9036 22980 9042
rect 22928 8978 22980 8984
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22284 7812 22336 7818
rect 22284 7754 22336 7760
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19616 6928 19668 6934
rect 19616 6870 19668 6876
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19168 6390 19196 6734
rect 19628 6458 19656 6870
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19156 6384 19208 6390
rect 19156 6326 19208 6332
rect 19168 5166 19196 6326
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 22112 5914 22140 7210
rect 22848 7002 22876 8774
rect 22940 8634 22968 8978
rect 23400 8906 23428 9318
rect 24492 9172 24544 9178
rect 24596 9160 24624 9386
rect 24872 9178 24900 13670
rect 24544 9132 24624 9160
rect 24492 9114 24544 9120
rect 24032 9104 24084 9110
rect 24032 9046 24084 9052
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 23400 8634 23428 8842
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23400 8430 23428 8570
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23952 8362 23980 8910
rect 24044 8498 24072 9046
rect 24596 9042 24624 9132
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24584 9036 24636 9042
rect 24584 8978 24636 8984
rect 25504 9036 25556 9042
rect 25504 8978 25556 8984
rect 27620 9036 27672 9042
rect 27620 8978 27672 8984
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 25516 8634 25544 8978
rect 27632 8945 27660 8978
rect 27618 8936 27674 8945
rect 27618 8871 27674 8880
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23952 8090 23980 8298
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 24768 7948 24820 7954
rect 24768 7890 24820 7896
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23768 7410 23796 7686
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23940 7404 23992 7410
rect 23940 7346 23992 7352
rect 23848 7268 23900 7274
rect 23848 7210 23900 7216
rect 22836 6996 22888 7002
rect 22836 6938 22888 6944
rect 22848 5914 22876 6938
rect 23860 6934 23888 7210
rect 23020 6928 23072 6934
rect 23020 6870 23072 6876
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23032 6254 23060 6870
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 23020 6248 23072 6254
rect 23020 6190 23072 6196
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22836 5908 22888 5914
rect 22836 5850 22888 5856
rect 23400 5846 23428 6326
rect 23860 6322 23888 6598
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 23400 5302 23428 5782
rect 23860 5370 23888 6258
rect 23952 5846 23980 7346
rect 24780 7206 24808 7890
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 24044 6322 24072 6734
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6458 24716 6802
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 23940 5840 23992 5846
rect 23940 5782 23992 5788
rect 24044 5710 24072 6258
rect 25228 6248 25280 6254
rect 25228 6190 25280 6196
rect 25240 5914 25268 6190
rect 25228 5908 25280 5914
rect 25228 5850 25280 5856
rect 25412 5772 25464 5778
rect 25412 5714 25464 5720
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24044 5370 24072 5646
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 25424 5370 25452 5714
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 25412 5364 25464 5370
rect 25412 5306 25464 5312
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 24858 5128 24914 5137
rect 24124 5092 24176 5098
rect 24858 5063 24914 5072
rect 24124 5034 24176 5040
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4690 20024 4966
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19996 4282 20024 4626
rect 24044 4593 24072 4966
rect 24030 4584 24086 4593
rect 24030 4519 24086 4528
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18524 3194 18552 3538
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 18524 2922 18552 3130
rect 18512 2916 18564 2922
rect 18512 2858 18564 2864
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17592 2848 17644 2854
rect 17592 2790 17644 2796
rect 17512 2650 17540 2790
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 17604 2446 17632 2790
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14646 82 14702 480
rect 14568 54 14702 82
rect 15672 82 15700 2314
rect 16026 82 16082 480
rect 15672 54 16082 82
rect 13726 31 13782 40
rect 14646 0 14702 54
rect 16026 0 16082 54
rect 17406 82 17462 480
rect 17788 82 17816 2518
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 18340 1873 18368 2450
rect 19984 2372 20036 2378
rect 19984 2314 20036 2320
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 19708 2304 19760 2310
rect 19708 2246 19760 2252
rect 18326 1864 18382 1873
rect 18326 1799 18382 1808
rect 17406 54 17816 82
rect 18432 82 18460 2246
rect 19720 1737 19748 2246
rect 19706 1728 19762 1737
rect 19706 1663 19762 1672
rect 18786 82 18842 480
rect 18432 54 18842 82
rect 19996 82 20024 2314
rect 20166 82 20222 480
rect 19996 54 20222 82
rect 21376 82 21404 4422
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 21638 82 21694 480
rect 21376 54 21694 82
rect 22664 82 22692 2246
rect 23018 82 23074 480
rect 22664 54 23074 82
rect 24136 82 24164 5034
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24872 4282 24900 5063
rect 24860 4276 24912 4282
rect 24860 4218 24912 4224
rect 25516 4154 25544 7142
rect 25594 6624 25650 6633
rect 25594 6559 25650 6568
rect 25608 6458 25636 6559
rect 25596 6452 25648 6458
rect 25596 6394 25648 6400
rect 27620 5092 27672 5098
rect 27620 5034 27672 5040
rect 27632 5001 27660 5034
rect 27618 4992 27674 5001
rect 27618 4927 27674 4936
rect 25516 4126 25636 4154
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24398 82 24454 480
rect 24136 54 24454 82
rect 25608 82 25636 4126
rect 26884 3936 26936 3942
rect 26884 3878 26936 3884
rect 25778 82 25834 480
rect 25608 54 25834 82
rect 26896 82 26924 3878
rect 27618 1048 27674 1057
rect 27618 983 27674 992
rect 27158 82 27214 480
rect 27632 105 27660 983
rect 26896 54 27214 82
rect 17406 0 17462 54
rect 18786 0 18842 54
rect 20166 0 20222 54
rect 21638 0 21694 54
rect 23018 0 23074 54
rect 24398 0 24454 54
rect 25778 0 25834 54
rect 27158 0 27214 54
rect 27618 96 27674 105
rect 27618 31 27674 40
<< via2 >>
rect 1214 24248 1270 24304
rect 1950 19760 2006 19816
rect 110 18128 166 18184
rect 1582 15408 1638 15464
rect 1214 13640 1270 13696
rect 1582 11192 1638 11248
rect 2226 10648 2282 10704
rect 1582 9152 1638 9208
rect 6274 26288 6330 26344
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 3054 12280 3110 12336
rect 2318 7928 2374 7984
rect 2594 7792 2650 7848
rect 110 7384 166 7440
rect 1582 4684 1638 4720
rect 1582 4664 1584 4684
rect 1584 4664 1636 4684
rect 1636 4664 1638 4684
rect 110 3032 166 3088
rect 2318 1944 2374 2000
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 6918 22072 6974 22128
rect 7286 21936 7342 21992
rect 6458 13776 6514 13832
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6918 12688 6974 12744
rect 6182 1536 6238 1592
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 9402 13776 9458 13832
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 9954 13776 10010 13832
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 8942 7656 8998 7712
rect 8942 7248 8998 7304
rect 9770 5480 9826 5536
rect 12530 17040 12586 17096
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 11794 10512 11850 10568
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3576 10194 3632
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 13542 21936 13598 21992
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 18602 23604 18604 23624
rect 18604 23604 18656 23624
rect 18656 23604 18658 23624
rect 18602 23568 18658 23604
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14646 20440 14702 20496
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 12622 13776 12678 13832
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 17498 17040 17554 17096
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15106 15952 15162 16008
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 12990 12280 13046 12336
rect 12530 7792 12586 7848
rect 12070 5072 12126 5128
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 16026 10648 16082 10704
rect 15658 10512 15714 10568
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14646 7656 14702 7712
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 10966 1808 11022 1864
rect 11794 1944 11850 2000
rect 12530 1672 12586 1728
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 17498 13368 17554 13424
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 21730 22072 21786 22128
rect 25134 26424 25190 26480
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24674 24384 24730 24440
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 26974 23568 27030 23624
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 27618 22888 27674 22944
rect 27618 21936 27674 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24674 18400 24730 18456
rect 22190 12688 22246 12744
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 16578 7248 16634 7304
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14094 5480 14150 5536
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 13726 40 13782 96
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 17406 7928 17462 7984
rect 18602 4528 18658 4584
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 25134 16360 25190 16416
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24858 15952 24914 16008
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 27618 15000 27674 15056
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 27618 13776 27674 13832
rect 24030 13368 24086 13424
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24674 12416 24730 12472
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 22926 10376 22982 10432
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 27618 8880 27674 8936
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24858 5072 24914 5128
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 24030 4528 24086 4584
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 18326 1808 18382 1864
rect 19706 1672 19762 1728
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25594 6568 25650 6624
rect 27618 4936 27674 4992
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 27618 992 27674 1048
rect 27618 40 27674 96
<< metal3 >>
rect 27520 26936 28000 27056
rect 0 26800 480 26920
rect 62 26346 122 26800
rect 25129 26482 25195 26485
rect 27662 26482 27722 26936
rect 25129 26480 27722 26482
rect 25129 26424 25134 26480
rect 25190 26424 27722 26480
rect 25129 26422 27722 26424
rect 25129 26419 25195 26422
rect 6269 26346 6335 26349
rect 62 26344 6335 26346
rect 62 26288 6274 26344
rect 6330 26288 6335 26344
rect 62 26286 6335 26288
rect 6269 26283 6335 26286
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 27520 24896 28000 25016
rect 0 24624 480 24744
rect 62 24306 122 24624
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 24669 24442 24735 24445
rect 27662 24442 27722 24896
rect 24669 24440 27722 24442
rect 24669 24384 24674 24440
rect 24730 24384 27722 24440
rect 24669 24382 27722 24384
rect 24669 24379 24735 24382
rect 1209 24306 1275 24309
rect 62 24304 1275 24306
rect 62 24248 1214 24304
rect 1270 24248 1275 24304
rect 62 24246 1275 24248
rect 1209 24243 1275 24246
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 18597 23626 18663 23629
rect 26969 23626 27035 23629
rect 18597 23624 27035 23626
rect 18597 23568 18602 23624
rect 18658 23568 26974 23624
rect 27030 23568 27035 23624
rect 18597 23566 27035 23568
rect 18597 23563 18663 23566
rect 26969 23563 27035 23566
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 27520 22944 28000 22976
rect 27520 22888 27618 22944
rect 27674 22888 28000 22944
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 27520 22856 28000 22888
rect 24277 22815 24597 22816
rect 0 22448 480 22568
rect 62 21994 122 22448
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 6913 22130 6979 22133
rect 21725 22130 21791 22133
rect 6913 22128 21791 22130
rect 6913 22072 6918 22128
rect 6974 22072 21730 22128
rect 21786 22072 21791 22128
rect 6913 22070 21791 22072
rect 6913 22067 6979 22070
rect 21725 22067 21791 22070
rect 7281 21994 7347 21997
rect 62 21992 7347 21994
rect 62 21936 7286 21992
rect 7342 21936 7347 21992
rect 62 21934 7347 21936
rect 7281 21931 7347 21934
rect 13537 21994 13603 21997
rect 27613 21994 27679 21997
rect 13537 21992 27679 21994
rect 13537 21936 13542 21992
rect 13598 21936 27618 21992
rect 27674 21936 27679 21992
rect 13537 21934 27679 21936
rect 13537 21931 13603 21934
rect 27613 21931 27679 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 27520 20952 28000 21072
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 14641 20498 14707 20501
rect 27662 20498 27722 20952
rect 14641 20496 27722 20498
rect 14641 20440 14646 20496
rect 14702 20440 27722 20496
rect 14641 20438 27722 20440
rect 14641 20435 14707 20438
rect 0 20272 480 20392
rect 62 19818 122 20272
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1945 19818 2011 19821
rect 62 19816 2011 19818
rect 62 19760 1950 19816
rect 2006 19760 2011 19816
rect 62 19758 2011 19760
rect 1945 19755 2011 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 27520 18912 28000 19032
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 24669 18458 24735 18461
rect 27662 18458 27722 18912
rect 24669 18456 27722 18458
rect 24669 18400 24674 18456
rect 24730 18400 27722 18456
rect 24669 18398 27722 18400
rect 24669 18395 24735 18398
rect 0 18184 480 18216
rect 0 18128 110 18184
rect 166 18128 480 18184
rect 0 18096 480 18128
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 12525 17098 12591 17101
rect 17493 17098 17559 17101
rect 12525 17096 17559 17098
rect 12525 17040 12530 17096
rect 12586 17040 17498 17096
rect 17554 17040 17559 17096
rect 12525 17038 17559 17040
rect 12525 17035 12591 17038
rect 17493 17035 17559 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 27520 16872 28000 16992
rect 19610 16831 19930 16832
rect 25129 16418 25195 16421
rect 27662 16418 27722 16872
rect 25129 16416 27722 16418
rect 25129 16360 25134 16416
rect 25190 16360 27722 16416
rect 25129 16358 27722 16360
rect 25129 16355 25195 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 15920 480 16040
rect 15101 16010 15167 16013
rect 24853 16010 24919 16013
rect 15101 16008 24919 16010
rect 15101 15952 15106 16008
rect 15162 15952 24858 16008
rect 24914 15952 24919 16008
rect 15101 15950 24919 15952
rect 15101 15947 15167 15950
rect 24853 15947 24919 15950
rect 62 15466 122 15920
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 1577 15466 1643 15469
rect 62 15464 1643 15466
rect 62 15408 1582 15464
rect 1638 15408 1643 15464
rect 62 15406 1643 15408
rect 1577 15403 1643 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 27520 15056 28000 15088
rect 27520 15000 27618 15056
rect 27674 15000 28000 15056
rect 27520 14968 28000 15000
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13880 480 14000
rect 62 13698 122 13880
rect 6453 13834 6519 13837
rect 9397 13834 9463 13837
rect 9949 13834 10015 13837
rect 6453 13832 10015 13834
rect 6453 13776 6458 13832
rect 6514 13776 9402 13832
rect 9458 13776 9954 13832
rect 10010 13776 10015 13832
rect 6453 13774 10015 13776
rect 6453 13771 6519 13774
rect 9397 13771 9463 13774
rect 9949 13771 10015 13774
rect 12617 13834 12683 13837
rect 27613 13834 27679 13837
rect 12617 13832 27679 13834
rect 12617 13776 12622 13832
rect 12678 13776 27618 13832
rect 27674 13776 27679 13832
rect 12617 13774 27679 13776
rect 12617 13771 12683 13774
rect 27613 13771 27679 13774
rect 1209 13698 1275 13701
rect 62 13696 1275 13698
rect 62 13640 1214 13696
rect 1270 13640 1275 13696
rect 62 13638 1275 13640
rect 1209 13635 1275 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 17493 13426 17559 13429
rect 24025 13426 24091 13429
rect 17493 13424 24091 13426
rect 17493 13368 17498 13424
rect 17554 13368 24030 13424
rect 24086 13368 24091 13424
rect 17493 13366 24091 13368
rect 17493 13363 17559 13366
rect 24025 13363 24091 13366
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 27520 12928 28000 13048
rect 6913 12746 6979 12749
rect 22185 12746 22251 12749
rect 6913 12744 22251 12746
rect 6913 12688 6918 12744
rect 6974 12688 22190 12744
rect 22246 12688 22251 12744
rect 6913 12686 22251 12688
rect 6913 12683 6979 12686
rect 22185 12683 22251 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 24669 12474 24735 12477
rect 27662 12474 27722 12928
rect 24669 12472 27722 12474
rect 24669 12416 24674 12472
rect 24730 12416 27722 12472
rect 24669 12414 27722 12416
rect 24669 12411 24735 12414
rect 3049 12338 3115 12341
rect 12985 12338 13051 12341
rect 3049 12336 13051 12338
rect 3049 12280 3054 12336
rect 3110 12280 12990 12336
rect 13046 12280 13051 12336
rect 3049 12278 13051 12280
rect 3049 12275 3115 12278
rect 12985 12275 13051 12278
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11704 480 11824
rect 62 11250 122 11704
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 1577 11250 1643 11253
rect 62 11248 1643 11250
rect 62 11192 1582 11248
rect 1638 11192 1643 11248
rect 62 11190 1643 11192
rect 1577 11187 1643 11190
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 27520 10888 28000 11008
rect 24277 10847 24597 10848
rect 2221 10706 2287 10709
rect 16021 10706 16087 10709
rect 2221 10704 16087 10706
rect 2221 10648 2226 10704
rect 2282 10648 16026 10704
rect 16082 10648 16087 10704
rect 2221 10646 16087 10648
rect 2221 10643 2287 10646
rect 16021 10643 16087 10646
rect 11789 10570 11855 10573
rect 15653 10570 15719 10573
rect 11789 10568 15719 10570
rect 11789 10512 11794 10568
rect 11850 10512 15658 10568
rect 15714 10512 15719 10568
rect 11789 10510 15719 10512
rect 11789 10507 11855 10510
rect 15653 10507 15719 10510
rect 22921 10434 22987 10437
rect 27662 10434 27722 10888
rect 22921 10432 27722 10434
rect 22921 10376 22926 10432
rect 22982 10376 27722 10432
rect 22921 10374 27722 10376
rect 22921 10371 22987 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 0 9528 480 9648
rect 62 9210 122 9528
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 1577 9210 1643 9213
rect 62 9208 1643 9210
rect 62 9152 1582 9208
rect 1638 9152 1643 9208
rect 62 9150 1643 9152
rect 1577 9147 1643 9150
rect 27520 8936 28000 8968
rect 27520 8880 27618 8936
rect 27674 8880 28000 8936
rect 27520 8848 28000 8880
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 2313 7986 2379 7989
rect 17401 7986 17467 7989
rect 2313 7984 17467 7986
rect 2313 7928 2318 7984
rect 2374 7928 17406 7984
rect 17462 7928 17467 7984
rect 2313 7926 17467 7928
rect 2313 7923 2379 7926
rect 17401 7923 17467 7926
rect 2589 7850 2655 7853
rect 12525 7850 12591 7853
rect 2589 7848 12591 7850
rect 2589 7792 2594 7848
rect 2650 7792 12530 7848
rect 12586 7792 12591 7848
rect 2589 7790 12591 7792
rect 2589 7787 2655 7790
rect 12525 7787 12591 7790
rect 8937 7714 9003 7717
rect 14641 7714 14707 7717
rect 8937 7712 14707 7714
rect 8937 7656 8942 7712
rect 8998 7656 14646 7712
rect 14702 7656 14707 7712
rect 8937 7654 14707 7656
rect 8937 7651 9003 7654
rect 14641 7651 14707 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 0 7440 480 7472
rect 0 7384 110 7440
rect 166 7384 480 7440
rect 0 7352 480 7384
rect 8937 7306 9003 7309
rect 16573 7306 16639 7309
rect 8937 7304 16639 7306
rect 8937 7248 8942 7304
rect 8998 7248 16578 7304
rect 16634 7248 16639 7304
rect 8937 7246 16639 7248
rect 8937 7243 9003 7246
rect 16573 7243 16639 7246
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 27520 6944 28000 7064
rect 25589 6626 25655 6629
rect 27662 6626 27722 6944
rect 25589 6624 27722 6626
rect 25589 6568 25594 6624
rect 25650 6568 27722 6624
rect 25589 6566 27722 6568
rect 25589 6563 25655 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 9765 5538 9831 5541
rect 14089 5538 14155 5541
rect 9765 5536 14155 5538
rect 9765 5480 9770 5536
rect 9826 5480 14094 5536
rect 14150 5480 14155 5536
rect 9765 5478 14155 5480
rect 9765 5475 9831 5478
rect 14089 5475 14155 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 0 5176 480 5296
rect 62 4722 122 5176
rect 12065 5130 12131 5133
rect 24853 5130 24919 5133
rect 12065 5128 24919 5130
rect 12065 5072 12070 5128
rect 12126 5072 24858 5128
rect 24914 5072 24919 5128
rect 12065 5070 24919 5072
rect 12065 5067 12131 5070
rect 24853 5067 24919 5070
rect 27520 4992 28000 5024
rect 27520 4936 27618 4992
rect 27674 4936 28000 4992
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 27520 4904 28000 4936
rect 19610 4863 19930 4864
rect 1577 4722 1643 4725
rect 62 4720 1643 4722
rect 62 4664 1582 4720
rect 1638 4664 1643 4720
rect 62 4662 1643 4664
rect 1577 4659 1643 4662
rect 18597 4586 18663 4589
rect 24025 4586 24091 4589
rect 18597 4584 24091 4586
rect 18597 4528 18602 4584
rect 18658 4528 24030 4584
rect 24086 4528 24091 4584
rect 18597 4526 24091 4528
rect 18597 4523 18663 4526
rect 24025 4523 24091 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 10133 3634 10199 3637
rect 10133 3632 27722 3634
rect 10133 3576 10138 3632
rect 10194 3576 27722 3632
rect 10133 3574 27722 3576
rect 10133 3571 10199 3574
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 0 3088 480 3120
rect 0 3032 110 3088
rect 166 3032 480 3088
rect 0 3000 480 3032
rect 27662 2984 27722 3574
rect 27520 2864 28000 2984
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 2313 2002 2379 2005
rect 11789 2002 11855 2005
rect 2313 2000 11855 2002
rect 2313 1944 2318 2000
rect 2374 1944 11794 2000
rect 11850 1944 11855 2000
rect 2313 1942 11855 1944
rect 2313 1939 2379 1942
rect 11789 1939 11855 1942
rect 10961 1866 11027 1869
rect 18321 1866 18387 1869
rect 10961 1864 18387 1866
rect 10961 1808 10966 1864
rect 11022 1808 18326 1864
rect 18382 1808 18387 1864
rect 10961 1806 18387 1808
rect 10961 1803 11027 1806
rect 18321 1803 18387 1806
rect 12525 1730 12591 1733
rect 19701 1730 19767 1733
rect 12525 1728 19767 1730
rect 12525 1672 12530 1728
rect 12586 1672 19706 1728
rect 19762 1672 19767 1728
rect 12525 1670 19767 1672
rect 12525 1667 12591 1670
rect 19701 1667 19767 1670
rect 6177 1594 6243 1597
rect 62 1592 6243 1594
rect 62 1536 6182 1592
rect 6238 1536 6243 1592
rect 62 1534 6243 1536
rect 62 1080 122 1534
rect 6177 1531 6243 1534
rect 0 960 480 1080
rect 27520 1048 28000 1080
rect 27520 992 27618 1048
rect 27674 992 28000 1048
rect 27520 960 28000 992
rect 13721 98 13787 101
rect 27613 98 27679 101
rect 13721 96 27679 98
rect 13721 40 13726 96
rect 13782 40 27618 96
rect 27674 40 27679 96
rect 13721 38 27679 40
rect 13721 35 13787 38
rect 27613 35 27679 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_1_54 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_62 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_60
timestamp 1586364061
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_67
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_66
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_70
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_90
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _234_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_99
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _198_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_148
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_144
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_152
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_165 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_165
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_173
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_169
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_173
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_181
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_187
timestamp 1586364061
transform 1 0 18308 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_191
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_191
timestamp 1586364061
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_195
timestamp 1586364061
transform 1 0 19044 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_202
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_206
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_198
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_202
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_214
timestamp 1586364061
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_226
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_237
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_0_245
timestamp 1586364061
transform 1 0 23644 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_238
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_6  FILLER_2_55
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_61
timestamp 1586364061
transform 1 0 6716 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use scs8hd_conb_1  _216_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_110
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_2_123
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_140
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_147
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 590 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_157
timestamp 1586364061
transform 1 0 15548 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_161
timestamp 1586364061
transform 1 0 15916 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_174
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_12  FILLER_2_191
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_203
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_54
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_58
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 774 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_85
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _158_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 130 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_182
timestamp 1586364061
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_187
timestamp 1586364061
transform 1 0 18308 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_191
timestamp 1586364061
transform 1 0 18676 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_216
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_228
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_253
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_262
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_3_274
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_69
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_73
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_77
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_100
timestamp 1586364061
transform 1 0 10304 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_136
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_187
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_191
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 406 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_69
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_or4_4  _157_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_73
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_97
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_107
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_120
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_128
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_145
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_162
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 314 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 18124 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_194
timestamp 1586364061
transform 1 0 18952 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_205
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_209
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23828 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_249
timestamp 1586364061
transform 1 0 24012 0 1 4896
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_262
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_266
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_274
timestamp 1586364061
transform 1 0 26312 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_60
timestamp 1586364061
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_68
timestamp 1586364061
transform 1 0 7360 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_1  _139_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 314 592
use scs8hd_or2_4  _099_
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 682 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_73
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_89
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_85
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_103
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_131
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_126
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_130
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_168
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_172
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_176
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_181
timestamp 1586364061
transform 1 0 17756 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_185
timestamp 1586364061
transform 1 0 18124 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_180
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_195
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_199
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_199
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 866 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_231
timestamp 1586364061
transform 1 0 22356 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_235
timestamp 1586364061
transform 1 0 22724 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_222
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_238
timestamp 1586364061
transform 1 0 23000 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_248
timestamp 1586364061
transform 1 0 23920 0 -1 5984
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_259
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_271
timestamp 1586364061
transform 1 0 26036 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_266
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_270
timestamp 1586364061
transform 1 0 25944 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_276
timestamp 1586364061
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 6072 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_52
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_63
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_67
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_8_111
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_132
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_137
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 314 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_143
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_151
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_159
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_8_167
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_180
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_197
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_209
timestamp 1586364061
transform 1 0 20332 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_235
timestamp 1586364061
transform 1 0 22724 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22816 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_245
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_249
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_8_262
timestamp 1586364061
transform 1 0 25208 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_46
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_50
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 7728 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_70
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 590 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_102
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_131
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_161
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_167
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_229
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_270
timestamp 1586364061
transform 1 0 25944 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_276
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_52
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_81
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_85
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_96
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_109
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_113
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_142
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_150
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_158
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_162
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_176
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_3  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_253
timestamp 1586364061
transform 1 0 24380 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_265
timestamp 1586364061
transform 1 0 25484 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_273
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_41
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 406 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 590 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_145
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_163
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_167
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_201
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_11_233
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 314 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_238
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_254
timestamp 1586364061
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_262
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_266
timestamp 1586364061
transform 1 0 25576 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_11_274
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_52
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 406 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_71
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_nor3_4  _168_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_101
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_12_116
timestamp 1586364061
transform 1 0 11776 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_135
timestamp 1586364061
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_12_167
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_235
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_12_256
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 6900 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_70
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_71
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_81
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_87
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_85
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_104
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_108
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_113
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_nor3_4  _170_
timestamp 1586364061
transform 1 0 13156 0 -1 10336
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_144
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_152
timestamp 1586364061
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 15364 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_160
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_164
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_183
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_205
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_195
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_207
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_241
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_249
timestamp 1586364061
transform 1 0 24012 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_256
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_261
timestamp 1586364061
transform 1 0 25116 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_268
timestamp 1586364061
transform 1 0 25760 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_273
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_45
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_49
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 774 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_70
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 314 592
use scs8hd_nor3_4  _169_
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_145
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_150
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_163
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_177
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_180
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_253
timestamp 1586364061
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_3  FILLER_16_40
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_52
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_60
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 9752 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 10580 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_101
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_114
timestamp 1586364061
transform 1 0 11592 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_134
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 406 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_158
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_170
timestamp 1586364061
transform 1 0 16744 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_258
timestamp 1586364061
transform 1 0 24840 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_270
timestamp 1586364061
transform 1 0 25944 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_9
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_13
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_25
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_33
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 406 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_88
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_109
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_138
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_157
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_170
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_229
timestamp 1586364061
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_241
timestamp 1586364061
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_75
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_81
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 590 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_148
timestamp 1586364061
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_183
timestamp 1586364061
transform 1 0 17940 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_186
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_198
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_6
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_10
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_24
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_28
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_43
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_49
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_81
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_96
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_85
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 10396 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_110
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_120
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_127
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_133
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_19_149
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_153
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_175
timestamp 1586364061
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_21
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_26
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_43
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_54
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_58
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_78
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_82
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_116
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_120
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 13156 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_133
timestamp 1586364061
transform 1 0 13340 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_144
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_148
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_167
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_170
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_182
timestamp 1586364061
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_189
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_201
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_213
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_225
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_237
timestamp 1586364061
transform 1 0 22908 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_243
timestamp 1586364061
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_251
timestamp 1586364061
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_255
timestamp 1586364061
transform 1 0 24564 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_267
timestamp 1586364061
transform 1 0 25668 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_275
timestamp 1586364061
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_45
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_49
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_61
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_6  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_6  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_158
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_162
timestamp 1586364061
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_165
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_22_179
timestamp 1586364061
transform 1 0 17572 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_185
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_196
timestamp 1586364061
transform 1 0 19136 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_208
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_258
timestamp 1586364061
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_270
timestamp 1586364061
transform 1 0 25944 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_21
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_33
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_37
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_50
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_54
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_78
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_82
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_108
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_115
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_119
timestamp 1586364061
transform 1 0 12052 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_128
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_151
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_178
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_201
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_213
timestamp 1586364061
transform 1 0 20700 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_225
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 1142 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_237
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_241
timestamp 1586364061
transform 1 0 23276 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_262
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_23_274
timestamp 1586364061
transform 1 0 26312 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_8  FILLER_24_49
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_101
timestamp 1586364061
transform 1 0 10396 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_116
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_128
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_162
timestamp 1586364061
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_175
timestamp 1586364061
transform 1 0 17204 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_192
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_247
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_19
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_56
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_60
timestamp 1586364061
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_69
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_82
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_103
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_116
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 590 592
use scs8hd_decap_8  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_131
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_139
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_152
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_164
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_172
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_176
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_180
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_209
timestamp 1586364061
transform 1 0 20332 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_233
timestamp 1586364061
transform 1 0 22540 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_241
timestamp 1586364061
transform 1 0 23276 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_262
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_25_274
timestamp 1586364061
transform 1 0 26312 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 3128 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_21
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_24
timestamp 1586364061
transform 1 0 3312 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_20
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 590 592
use scs8hd_decap_6  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_30
timestamp 1586364061
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_38
timestamp 1586364061
transform 1 0 4600 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 5520 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_43
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_55
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_57
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_26_69
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_67
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_90
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_6  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_135
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_165
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_187
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_191
timestamp 1586364061
transform 1 0 18676 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 1142 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_198
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_205
timestamp 1586364061
transform 1 0 19964 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_229
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_241
timestamp 1586364061
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_13
timestamp 1586364061
transform 1 0 2300 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_46
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_60
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 1142 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_101
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_134
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_200
timestamp 1586364061
transform 1 0 19504 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_258
timestamp 1586364061
transform 1 0 24840 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_270
timestamp 1586364061
transform 1 0 25944 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_274
timestamp 1586364061
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_31
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_67
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_102
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_144
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_168
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 18584 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_188
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_192
timestamp 1586364061
transform 1 0 18768 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_204
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_216
timestamp 1586364061
transform 1 0 20976 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_228
timestamp 1586364061
transform 1 0 22080 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_248
timestamp 1586364061
transform 1 0 23920 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_252
timestamp 1586364061
transform 1 0 24288 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_264
timestamp 1586364061
transform 1 0 25392 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_29_276
timestamp 1586364061
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_17
timestamp 1586364061
transform 1 0 2668 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_21
timestamp 1586364061
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_24
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 590 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_46
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_59
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 1142 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_71
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_81
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_85
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_121
timestamp 1586364061
transform 1 0 12236 0 -1 19040
box -38 -48 774 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_132
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_144
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_31_77
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_102
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_112
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_120
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_126
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_130
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_134
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_140
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_144
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_148
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_160
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_172
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_180
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 4784 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_43
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_32_60
timestamp 1586364061
transform 1 0 6624 0 -1 20128
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_72
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_32_119
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_127
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_132
timestamp 1586364061
transform 1 0 13248 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_144
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_66
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_69
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_64
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_70
timestamp 1586364061
transform 1 0 7544 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_78
timestamp 1586364061
transform 1 0 8280 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_82
timestamp 1586364061
transform 1 0 8648 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_89
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_93
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_90
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_106
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_114
timestamp 1586364061
transform 1 0 11592 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_137
timestamp 1586364061
transform 1 0 13708 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_144
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_156
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_168
timestamp 1586364061
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_180
timestamp 1586364061
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_77
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 1142 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_89
timestamp 1586364061
transform 1 0 9292 0 1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_35_96
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_104
timestamp 1586364061
transform 1 0 10672 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_113
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_117
timestamp 1586364061
transform 1 0 11868 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_148
timestamp 1586364061
transform 1 0 14720 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_160
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_172
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_48
timestamp 1586364061
transform 1 0 5520 0 -1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_60
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_64
timestamp 1586364061
transform 1 0 6992 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_72
timestamp 1586364061
transform 1 0 7728 0 -1 22304
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_109
timestamp 1586364061
transform 1 0 11132 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_113
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_121
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 314 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  FILLER_37_77
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_89
timestamp 1586364061
transform 1 0 9292 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_99
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 1142 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_111
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_37_119
timestamp 1586364061
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 12972 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_127
timestamp 1586364061
transform 1 0 12788 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_131
timestamp 1586364061
transform 1 0 13156 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_143
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_155
timestamp 1586364061
transform 1 0 15364 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_167
timestamp 1586364061
transform 1 0 16468 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_18
timestamp 1586364061
transform 1 0 2760 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_30
timestamp 1586364061
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5336 0 -1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_55
timestamp 1586364061
transform 1 0 6164 0 -1 23392
box -38 -48 590 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_61
timestamp 1586364061
transform 1 0 6716 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_67
timestamp 1586364061
transform 1 0 7268 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_38_71
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_88
timestamp 1586364061
transform 1 0 9200 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_114
timestamp 1586364061
transform 1 0 11592 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_126
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_138
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_38_150
timestamp 1586364061
transform 1 0 14904 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_258
timestamp 1586364061
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_270
timestamp 1586364061
transform 1 0 25944 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_274
timestamp 1586364061
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_19
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_31
timestamp 1586364061
transform 1 0 3956 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_36
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_40
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_52
timestamp 1586364061
transform 1 0 5888 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_56
timestamp 1586364061
transform 1 0 6256 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6348 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_60
timestamp 1586364061
transform 1 0 6624 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_71
timestamp 1586364061
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_75
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_71
timestamp 1586364061
transform 1 0 7636 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_82
timestamp 1586364061
transform 1 0 8648 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_88
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_90
timestamp 1586364061
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_105
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_109
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_97
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_101
timestamp 1586364061
transform 1 0 10396 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_113
timestamp 1586364061
transform 1 0 11500 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_137
timestamp 1586364061
transform 1 0 13708 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_146
timestamp 1586364061
transform 1 0 14536 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_149
timestamp 1586364061
transform 1 0 14812 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_182
timestamp 1586364061
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_187
timestamp 1586364061
transform 1 0 18308 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_191
timestamp 1586364061
transform 1 0 18676 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_202
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_206
timestamp 1586364061
transform 1 0 20056 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_218
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal3 s 27520 960 28000 1080 6 address[0]
port 0 nsew default input
rlabel metal2 s 3422 0 3478 480 6 address[1]
port 1 nsew default input
rlabel metal3 s 27520 2864 28000 2984 6 address[2]
port 2 nsew default input
rlabel metal2 s 4802 0 4858 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 6182 0 6238 480 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 960 480 1080 6 address[5]
port 5 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chanx_right_in[0]
port 6 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_right_in[1]
port 7 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chanx_right_in[2]
port 8 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_right_in[3]
port 9 nsew default input
rlabel metal2 s 938 27520 994 28000 6 chanx_right_in[4]
port 10 nsew default input
rlabel metal2 s 2778 27520 2834 28000 6 chanx_right_in[5]
port 11 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chanx_right_in[6]
port 12 nsew default input
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_in[7]
port 13 nsew default input
rlabel metal3 s 0 7352 480 7472 6 chanx_right_in[8]
port 14 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chanx_right_out[0]
port 15 nsew default tristate
rlabel metal2 s 4618 27520 4674 28000 6 chanx_right_out[1]
port 16 nsew default tristate
rlabel metal2 s 6458 27520 6514 28000 6 chanx_right_out[2]
port 17 nsew default tristate
rlabel metal2 s 13174 0 13230 480 6 chanx_right_out[3]
port 18 nsew default tristate
rlabel metal2 s 14646 0 14702 480 6 chanx_right_out[4]
port 19 nsew default tristate
rlabel metal3 s 27520 6944 28000 7064 6 chanx_right_out[5]
port 20 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 chanx_right_out[6]
port 21 nsew default tristate
rlabel metal3 s 0 9528 480 9648 6 chanx_right_out[7]
port 22 nsew default tristate
rlabel metal3 s 0 11704 480 11824 6 chanx_right_out[8]
port 23 nsew default tristate
rlabel metal3 s 27520 8848 28000 8968 6 chany_top_in[0]
port 24 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 17406 0 17462 480 6 chany_top_in[2]
port 26 nsew default input
rlabel metal2 s 10230 27520 10286 28000 6 chany_top_in[3]
port 27 nsew default input
rlabel metal3 s 27520 10888 28000 11008 6 chany_top_in[4]
port 28 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 12070 27520 12126 28000 6 chany_top_in[6]
port 30 nsew default input
rlabel metal2 s 18786 0 18842 480 6 chany_top_in[7]
port 31 nsew default input
rlabel metal3 s 27520 12928 28000 13048 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal2 s 15842 27520 15898 28000 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal3 s 0 18096 480 18216 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal2 s 20166 0 20222 480 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal2 s 17682 27520 17738 28000 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal2 s 21638 0 21694 480 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal2 s 19522 27520 19578 28000 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal3 s 27520 14968 28000 15088 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 2042 0 2098 480 6 data_in
port 42 nsew default input
rlabel metal2 s 662 0 718 480 6 enable
port 43 nsew default input
rlabel metal3 s 27520 20952 28000 21072 6 right_bottom_grid_pin_11_
port 44 nsew default input
rlabel metal3 s 27520 22856 28000 22976 6 right_bottom_grid_pin_13_
port 45 nsew default input
rlabel metal2 s 23294 27520 23350 28000 6 right_bottom_grid_pin_15_
port 46 nsew default input
rlabel metal3 s 27520 16872 28000 16992 6 right_bottom_grid_pin_1_
port 47 nsew default input
rlabel metal2 s 21362 27520 21418 28000 6 right_bottom_grid_pin_3_
port 48 nsew default input
rlabel metal3 s 27520 18912 28000 19032 6 right_bottom_grid_pin_5_
port 49 nsew default input
rlabel metal2 s 23018 0 23074 480 6 right_bottom_grid_pin_7_
port 50 nsew default input
rlabel metal2 s 24398 0 24454 480 6 right_bottom_grid_pin_9_
port 51 nsew default input
rlabel metal2 s 25778 0 25834 480 6 right_top_grid_pin_10_
port 52 nsew default input
rlabel metal3 s 0 22448 480 22568 6 top_left_grid_pin_11_
port 53 nsew default input
rlabel metal3 s 0 24624 480 24744 6 top_left_grid_pin_13_
port 54 nsew default input
rlabel metal2 s 26974 27520 27030 28000 6 top_left_grid_pin_15_
port 55 nsew default input
rlabel metal2 s 25134 27520 25190 28000 6 top_left_grid_pin_1_
port 56 nsew default input
rlabel metal3 s 27520 24896 28000 25016 6 top_left_grid_pin_3_
port 57 nsew default input
rlabel metal2 s 27158 0 27214 480 6 top_left_grid_pin_5_
port 58 nsew default input
rlabel metal3 s 27520 26936 28000 27056 6 top_left_grid_pin_7_
port 59 nsew default input
rlabel metal3 s 0 20272 480 20392 6 top_left_grid_pin_9_
port 60 nsew default input
rlabel metal3 s 0 26800 480 26920 6 top_right_grid_pin_11_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
