* NGSPICE file created from sb_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

.subckt sb_1__0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11]
+ chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16]
+ chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11]
+ chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16]
+ chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11]
+ chanx_right_out[12] chanx_right_out[13] chanx_right_out[14] chanx_right_out[15]
+ chanx_right_out[16] chanx_right_out[17] chanx_right_out[18] chanx_right_out[19]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_top_in[0]
+ chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14]
+ chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19]
+ chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5]
+ chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0]
+ chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14]
+ chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19]
+ chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9] left_bottom_grid_pin_1_
+ left_top_grid_pin_42_ left_top_grid_pin_43_ left_top_grid_pin_44_ left_top_grid_pin_45_
+ left_top_grid_pin_46_ left_top_grid_pin_47_ left_top_grid_pin_48_ left_top_grid_pin_49_
+ prog_clk right_bottom_grid_pin_1_ right_top_grid_pin_42_ right_top_grid_pin_43_
+ right_top_grid_pin_44_ right_top_grid_pin_45_ right_top_grid_pin_46_ right_top_grid_pin_47_
+ right_top_grid_pin_48_ right_top_grid_pin_49_ top_left_grid_pin_34_ top_left_grid_pin_35_
+ top_left_grid_pin_36_ top_left_grid_pin_37_ top_left_grid_pin_38_ top_left_grid_pin_39_
+ top_left_grid_pin_40_ top_left_grid_pin_41_ vpwr vgnd
XFILLER_39_266 vpwr vgnd scs8hd_fill_2
Xmem_right_track_2.scs8hd_dfxbp_1_3_ prog_clk mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l4_in_0_/S
+ mem_right_track_2.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_0.mux_l2_in_3__A0 _060_/HI vgnd vpwr scs8hd_diode_2
XFILLER_26_74 vgnd vpwr scs8hd_fill_1
XFILLER_13_133 vpwr vgnd scs8hd_fill_2
XFILLER_42_51 vpwr vgnd scs8hd_fill_2
XFILLER_9_115 vpwr vgnd scs8hd_fill_2
XFILLER_13_177 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A1 mux_left_track_25.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_228 vpwr vgnd scs8hd_fill_2
XFILLER_27_214 vgnd vpwr scs8hd_fill_1
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_36.mux_l2_in_0__A0 _048_/HI vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_32_250 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 top_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_15_206 vgnd vpwr scs8hd_decap_4
XFILLER_23_272 vgnd vpwr scs8hd_decap_4
X_062_ _062_/HI _062_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_23_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l1_in_2__A1 left_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_209 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.mux_l3_in_0_ mux_top_track_10.mux_l2_in_1_/X mux_top_track_10.mux_l2_in_0_/X
+ mux_top_track_10.mux_l3_in_0_/S mux_top_track_10.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_28.mux_l2_in_0__A1 mux_top_track_28.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_3__S mux_left_track_25.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_1.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_1.mux_l2_in_2_/S mux_left_track_1.mux_l3_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_42 vpwr vgnd scs8hd_fill_2
XFILLER_18_64 vpwr vgnd scs8hd_fill_2
XFILLER_18_75 vpwr vgnd scs8hd_fill_2
XFILLER_11_220 vpwr vgnd scs8hd_fill_2
XFILLER_11_231 vpwr vgnd scs8hd_fill_2
XFILLER_11_275 vpwr vgnd scs8hd_fill_2
X_114_ _114_/A chany_top_out[11] vgnd vpwr scs8hd_buf_2
X_045_ _045_/HI _045_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_106 vpwr vgnd scs8hd_fill_2
Xmem_top_track_14.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_12.mux_l2_in_0_/S mux_top_track_14.mux_l1_in_0_/S
+ mem_top_track_14.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_33.mux_l2_in_1__A1 mux_left_track_33.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__S mux_left_track_17.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__D mux_right_track_16.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_41 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.mux_l2_in_1_ _035_/HI chanx_left_in[9] mux_top_track_10.mux_l2_in_0_/S
+ mux_top_track_10.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_36.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__S mux_right_track_16.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_33.scs8hd_buf_4_0__A mux_left_track_33.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_161 vgnd vpwr scs8hd_decap_4
XFILLER_34_164 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_40_167 vgnd vpwr scs8hd_decap_6
XFILLER_40_145 vpwr vgnd scs8hd_fill_2
XFILLER_40_134 vgnd vpwr scs8hd_decap_6
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_20 vgnd vpwr scs8hd_decap_4
XFILLER_25_197 vpwr vgnd scs8hd_fill_2
XFILLER_31_97 vpwr vgnd scs8hd_fill_2
XFILLER_31_75 vgnd vpwr scs8hd_decap_4
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.scs8hd_dfxbp_1_1__D mux_top_track_10.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l2_in_1__S mux_top_track_0.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_16_186 vgnd vpwr scs8hd_fill_1
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_33.mux_l3_in_0__A1 mux_left_track_33.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_234 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_30.scs8hd_dfxbp_1_1__D mux_top_track_30.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_112 vpwr vgnd scs8hd_fill_2
XFILLER_22_123 vgnd vpwr scs8hd_decap_3
XFILLER_22_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_2__A0 left_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l1_in_2__S mux_top_track_6.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l3_in_0_/S
+ mem_right_track_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_0.mux_l2_in_3__A1 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_13_123 vgnd vpwr scs8hd_fill_1
XFILLER_13_156 vpwr vgnd scs8hd_fill_2
XFILLER_42_85 vpwr vgnd scs8hd_fill_2
XFILLER_9_127 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D mux_top_track_8.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_193 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_6.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_4
XFILLER_10_126 vpwr vgnd scs8hd_fill_2
XFILLER_10_137 vpwr vgnd scs8hd_fill_2
XFILLER_10_159 vpwr vgnd scs8hd_fill_2
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_99 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_36.mux_l2_in_0__A1 mux_top_track_36.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_215 vpwr vgnd scs8hd_fill_2
XFILLER_41_240 vpwr vgnd scs8hd_fill_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l3_in_1__A0 mux_left_track_9.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_270 vpwr vgnd scs8hd_fill_2
XFILLER_24_207 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XFILLER_23_240 vpwr vgnd scs8hd_fill_2
X_061_ _061_/HI _061_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XFILLER_14_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_30.mux_l2_in_0__S mux_top_track_30.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_9.scs8hd_dfxbp_1_3_ prog_clk mux_left_track_9.mux_l3_in_1_/S mux_left_track_9.mux_l4_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_210 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_2__S mux_left_track_1.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_243 vpwr vgnd scs8hd_fill_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_1.mux_l1_in_0_/S mux_left_track_1.mux_l2_in_2_/S
+ mem_left_track_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_32 vgnd vpwr scs8hd_decap_4
XFILLER_18_87 vpwr vgnd scs8hd_fill_2
X_113_ _113_/A chany_top_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_34_97 vpwr vgnd scs8hd_fill_2
XFILLER_11_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l4_in_0__A0 mux_left_track_9.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.scs8hd_buf_4_0__A mux_top_track_12.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_2__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_044_ _044_/HI _044_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_12.scs8hd_dfxbp_1_0__D mux_top_track_10.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__S mux_left_track_5.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_195 vpwr vgnd scs8hd_fill_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D mux_top_track_30.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l3_in_0__S mux_right_track_8.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_11 vpwr vgnd scs8hd_fill_2
XFILLER_20_66 vpwr vgnd scs8hd_fill_2
XFILLER_20_88 vgnd vpwr scs8hd_fill_1
XFILLER_29_86 vpwr vgnd scs8hd_fill_2
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.mux_l2_in_0_ chanx_right_in[19] mux_top_track_10.mux_l1_in_0_/X
+ mux_top_track_10.mux_l2_in_0_/S mux_top_track_10.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_38.scs8hd_buf_4_0__A mux_top_track_38.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_6.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l3_in_0_/S
+ mem_top_track_6.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_40_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_77 vpwr vgnd scs8hd_fill_2
Xmux_top_track_18.scs8hd_buf_4_0_ mux_top_track_18.mux_l2_in_0_/X _116_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
Xmux_right_track_8.mux_l2_in_3_ _033_/HI chanx_left_in[16] mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_121 vpwr vgnd scs8hd_fill_2
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_3_ _034_/HI chanx_left_in[2] mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_9.mux_l2_in_2__A1 left_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l2_in_1_/S
+ mem_right_track_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_10 vpwr vgnd scs8hd_fill_2
XFILLER_26_43 vpwr vgnd scs8hd_fill_2
XFILLER_9_139 vgnd vpwr scs8hd_decap_8
XFILLER_42_75 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_33.mux_l1_in_1__S mux_left_track_33.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l2_in_1__S mux_right_track_32.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l2_in_0__A0 chanx_right_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_8_183 vpwr vgnd scs8hd_fill_2
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_3__A0 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XFILLER_37_20 vpwr vgnd scs8hd_fill_2
XFILLER_18_227 vpwr vgnd scs8hd_fill_2
XFILLER_38_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l3_in_1__A1 mux_left_track_9.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_260 vpwr vgnd scs8hd_fill_2
XFILLER_24_219 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S mux_right_track_8.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_66 vgnd vpwr scs8hd_decap_4
X_060_ _060_/HI _060_/LO vgnd vpwr scs8hd_conb_1
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S mux_top_track_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_16.mux_l2_in_0__S mux_top_track_16.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_14_274 vgnd vpwr scs8hd_fill_1
XFILLER_36_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_2__A0 mux_right_track_4.mux_l1_in_5_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_9.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_9.mux_l2_in_0_/S mux_left_track_9.mux_l3_in_1_/S
+ mem_left_track_9.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_11 vpwr vgnd scs8hd_fill_2
XFILLER_18_22 vgnd vpwr scs8hd_decap_6
XFILLER_34_10 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_32.mux_l3_in_0_/S mux_left_track_1.mux_l1_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
X_112_ top_left_grid_pin_35_ chany_top_out[13] vgnd vpwr scs8hd_buf_2
X_043_ _043_/HI _043_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_9.mux_l4_in_0__A1 mux_left_track_9.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_23 vgnd vpwr scs8hd_decap_4
XFILLER_20_45 vpwr vgnd scs8hd_fill_2
XFILLER_29_65 vgnd vpwr scs8hd_decap_3
XFILLER_29_21 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l3_in_1__A0 mux_right_track_4.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_111 vpwr vgnd scs8hd_fill_2
XFILLER_34_188 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D mux_right_track_0.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_6.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_6.mux_l1_in_0_/S mux_top_track_6.mux_l2_in_0_/S
+ mem_top_track_6.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_25_155 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_25.mux_l2_in_1__S mux_left_track_25.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_2_ chanx_left_in[6] right_bottom_grid_pin_1_ mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_100 vgnd vpwr scs8hd_decap_4
XFILLER_31_169 vpwr vgnd scs8hd_fill_2
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_177 vgnd vpwr scs8hd_decap_3
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_2_ chanx_left_in[0] chanx_right_in[2] mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmem_top_track_22.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_22.mux_l1_in_1_/S mux_top_track_22.mux_l2_in_0_/S
+ mem_top_track_22.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_191 vgnd vpwr scs8hd_decap_4
Xmux_top_track_10.mux_l1_in_0_ chanx_right_in[9] top_left_grid_pin_35_ mux_top_track_10.mux_l1_in_0_/S
+ mux_top_track_10.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 top_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l4_in_0__A0 mux_right_track_4.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_0.mux_l4_in_0_/S mux_right_track_2.mux_l1_in_1_/S
+ mem_right_track_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_66 vpwr vgnd scs8hd_fill_2
XFILLER_42_32 vgnd vpwr scs8hd_decap_3
XFILLER_42_10 vpwr vgnd scs8hd_fill_2
Xmux_top_track_22.mux_l2_in_0_ mux_top_track_22.mux_l1_in_1_/X mux_top_track_22.mux_l1_in_0_/X
+ mux_top_track_22.mux_l2_in_0_/S mux_top_track_22.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_88 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_21_180 vgnd vpwr scs8hd_fill_1
XFILLER_36_206 vpwr vgnd scs8hd_fill_2
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_239 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l2_in_0__A1 mux_top_track_10.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_209 vpwr vgnd scs8hd_fill_2
XFILLER_27_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0__S mux_left_track_3.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_272 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_3__A1 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_18_206 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_fill_1
XFILLER_37_98 vpwr vgnd scs8hd_fill_2
XFILLER_37_43 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_2__S mux_top_track_2.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0__A0 mux_top_track_2.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
Xmux_top_track_22.mux_l1_in_1_ _042_/HI chanx_left_in[17] mux_top_track_22.mux_l1_in_1_/S
+ mux_top_track_22.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l2_in_0__S mux_top_track_6.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_23_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l2_in_2__A1 mux_right_track_4.mux_l1_in_4_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_9.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_top_track_34.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_top_track_34.scs8hd_buf_4_0_ mux_top_track_34.mux_l2_in_0_/X _108_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D mux_right_track_2.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_2__A0 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_256 vgnd vpwr scs8hd_decap_8
XFILLER_20_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_88 vpwr vgnd scs8hd_fill_2
XFILLER_34_77 vpwr vgnd scs8hd_fill_2
XFILLER_34_55 vpwr vgnd scs8hd_fill_2
X_111_ _111_/A chany_top_out[14] vgnd vpwr scs8hd_buf_2
X_042_ _042_/HI _042_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_249 vgnd vpwr scs8hd_decap_12
XFILLER_11_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D mux_top_track_16.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_37_131 vpwr vgnd scs8hd_fill_2
XFILLER_29_109 vgnd vpwr scs8hd_decap_3
XFILLER_37_175 vpwr vgnd scs8hd_fill_2
XFILLER_37_164 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__072__A chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_28_197 vgnd vpwr scs8hd_decap_3
XFILLER_28_164 vpwr vgnd scs8hd_fill_2
XFILLER_28_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_36.scs8hd_dfxbp_1_1__D mux_top_track_36.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l3_in_1__A1 mux_right_track_4.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l3_in_1__A0 mux_top_track_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_20.mux_l1_in_0__S mux_top_track_20.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_145 vpwr vgnd scs8hd_fill_2
XFILLER_34_134 vpwr vgnd scs8hd_fill_2
XFILLER_34_101 vgnd vpwr scs8hd_fill_1
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
Xmem_top_track_6.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_4.mux_l3_in_0_/S mux_top_track_6.mux_l1_in_0_/S
+ mem_top_track_6.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_0.mux_l2_in_2__S mux_right_track_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__S mux_left_track_1.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__067__A chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_31_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D mux_left_track_25.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
Xmux_right_track_8.mux_l2_in_1_ right_top_grid_pin_46_ right_top_grid_pin_42_ mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_134 vgnd vpwr scs8hd_decap_8
XFILLER_16_145 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ chanx_right_in[1] top_left_grid_pin_40_ mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_top_track_22.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_20.mux_l2_in_0_/S mux_top_track_22.mux_l1_in_1_/S
+ mem_top_track_22.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l4_in_0__A1 mux_right_track_4.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A1 top_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_42_99 vpwr vgnd scs8hd_fill_2
XFILLER_42_55 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_4
XFILLER_9_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l4_in_0__A0 mux_top_track_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_170 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.scs8hd_buf_4_0_ mux_left_track_9.mux_l4_in_0_/X _081_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_36_218 vgnd vpwr scs8hd_decap_3
XFILLER_29_270 vpwr vgnd scs8hd_fill_2
XFILLER_8_196 vgnd vpwr scs8hd_decap_4
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XFILLER_12_170 vpwr vgnd scs8hd_fill_2
XFILLER_35_262 vpwr vgnd scs8hd_fill_2
XFILLER_35_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D mux_right_track_2.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__080__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_37_66 vgnd vpwr scs8hd_decap_3
XFILLER_37_33 vpwr vgnd scs8hd_fill_2
XFILLER_41_254 vpwr vgnd scs8hd_fill_2
XFILLER_41_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_2.scs8hd_buf_4_0_ mux_top_track_2.mux_l3_in_0_/X _124_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_17_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_0__A1 mux_top_track_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_32_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_18.scs8hd_dfxbp_1_0__D mux_top_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0__A0 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A0 mux_left_track_1.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_22.mux_l1_in_0_ chanx_right_in[17] top_left_grid_pin_41_ mux_top_track_22.mux_l1_in_1_/S
+ mux_top_track_22.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__075__A chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_23_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_34.mux_l2_in_0_ _047_/HI mux_top_track_34.mux_l1_in_0_/X mux_top_track_34.mux_l2_in_0_/S
+ mux_top_track_34.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_38.scs8hd_dfxbp_1_0__D mux_top_track_36.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
Xmem_left_track_9.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_5.mux_l4_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_0.mux_l2_in_2__A1 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_18_46 vgnd vpwr scs8hd_decap_3
XFILLER_18_79 vpwr vgnd scs8hd_fill_2
X_110_ _110_/A chany_top_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_34_23 vpwr vgnd scs8hd_fill_2
XFILLER_11_224 vgnd vpwr scs8hd_decap_4
XFILLER_11_235 vpwr vgnd scs8hd_fill_2
X_041_ _041_/HI _041_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_12.mux_l2_in_0__S mux_top_track_12.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_45 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_14.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_18.mux_l1_in_1__S mux_top_track_18.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_154 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l3_in_1__A1 mux_top_track_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_110 vgnd vpwr scs8hd_decap_8
XFILLER_19_165 vgnd vpwr scs8hd_fill_1
XFILLER_34_168 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__D mux_right_track_4.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_149 vpwr vgnd scs8hd_fill_2
XFILLER_31_24 vgnd vpwr scs8hd_fill_1
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XANTENNA__083__A _083_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_ chany_top_in[16] mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_138 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ top_left_grid_pin_38_ mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_20.scs8hd_buf_4_0__A mux_top_track_20.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_116 vpwr vgnd scs8hd_fill_2
XFILLER_22_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_13_127 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l4_in_0__A1 mux_top_track_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA__078__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_42_89 vgnd vpwr scs8hd_decap_4
XFILLER_42_67 vpwr vgnd scs8hd_fill_2
XFILLER_42_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_6__A0 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_22.mux_l1_in_0__A0 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_16_90 vpwr vgnd scs8hd_fill_2
XFILLER_12_193 vpwr vgnd scs8hd_fill_2
XFILLER_35_230 vgnd vpwr scs8hd_decap_4
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l3_in_0__A0 mux_right_track_8.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_266 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XFILLER_17_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_14.mux_l1_in_0__A1 top_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A1 mux_left_track_1.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_23_36 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_14_222 vgnd vpwr scs8hd_fill_1
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
XFILLER_14_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l1_in_0__A0 top_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_28.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_58 vgnd vpwr scs8hd_decap_4
XANTENNA__086__A chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_11_203 vpwr vgnd scs8hd_fill_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
X_040_ _040_/HI _040_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_2.mux_l2_in_0__S mux_top_track_2.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
XFILLER_37_199 vgnd vpwr scs8hd_fill_1
XFILLER_37_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 chanx_right_in[7] vgnd vpwr scs8hd_diode_2
Xmux_top_track_34.mux_l1_in_0_ chanx_left_in[7] top_left_grid_pin_39_ mux_top_track_34.mux_l1_in_0_/S
+ mux_top_track_34.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_29_13 vpwr vgnd scs8hd_fill_2
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
XFILLER_19_144 vpwr vgnd scs8hd_fill_2
XFILLER_19_199 vpwr vgnd scs8hd_fill_2
XFILLER_42_191 vgnd vpwr scs8hd_decap_12
XFILLER_40_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D mux_right_track_24.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XFILLER_25_136 vpwr vgnd scs8hd_fill_2
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_31_36 vpwr vgnd scs8hd_fill_2
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_30.mux_l1_in_0__A0 chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A0 mux_top_track_4.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_22_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_38_261 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA__094__A chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_26_36 vgnd vpwr scs8hd_decap_4
XFILLER_13_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_6__A1 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_22.mux_l1_in_0__A1 top_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XFILLER_8_154 vgnd vpwr scs8hd_decap_3
XFILLER_8_187 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_1__S mux_left_track_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[9] chany_top_in[2] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D mux_right_track_8.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l3_in_0__A1 mux_right_track_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_38.mux_l1_in_0__S mux_top_track_38.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A _089_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A0 mux_top_track_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_223 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_36_ top_left_grid_pin_34_ mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l4_in_0__S mux_top_track_0.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_32_223 vgnd vpwr scs8hd_decap_3
XFILLER_32_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_30.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 mux_right_track_16.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_245 vpwr vgnd scs8hd_fill_2
XFILLER_23_256 vpwr vgnd scs8hd_fill_2
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XFILLER_14_201 vpwr vgnd scs8hd_fill_2
XFILLER_14_245 vpwr vgnd scs8hd_fill_2
Xmem_top_track_30.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_30.mux_l1_in_0_/S mux_top_track_30.mux_l2_in_0_/S
+ mem_top_track_30.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0__A1 top_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_20_215 vpwr vgnd scs8hd_fill_2
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
XFILLER_11_248 vpwr vgnd scs8hd_fill_2
XFILLER_11_259 vpwr vgnd scs8hd_fill_2
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_3 vgnd vpwr scs8hd_decap_4
X_099_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_37_123 vpwr vgnd scs8hd_fill_2
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_49 vpwr vgnd scs8hd_fill_2
XFILLER_28_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_20.scs8hd_dfxbp_1_0__D mux_top_track_18.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_115 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vgnd vpwr scs8hd_fill_1
XFILLER_42_170 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_24.mux_l1_in_1__A0 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XFILLER_33_192 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l3_in_0_/S
+ mem_right_track_16.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_30.mux_l1_in_0__A1 top_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_6_ chanx_left_in[14] chanx_left_in[5] mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_6_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_104 vgnd vpwr scs8hd_fill_1
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_28.scs8hd_buf_4_0__A mux_top_track_28.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A1 mux_top_track_4.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_1__S mux_top_track_14.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 _038_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_1__A0 left_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_38_273 vpwr vgnd scs8hd_fill_2
XFILLER_38_240 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_4
XFILLER_29_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 mux_right_track_24.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_166 vpwr vgnd scs8hd_fill_2
XFILLER_35_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_3__A0 _053_/HI vgnd vpwr scs8hd_diode_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_232 vgnd vpwr scs8hd_decap_4
XFILLER_26_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A1 mux_top_track_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A0 mux_top_track_16.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A0 mux_left_track_3.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_3.mux_l2_in_3_ _056_/HI left_top_grid_pin_49_ mux_left_track_3.mux_l2_in_2_/S
+ mux_left_track_3.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XFILLER_17_254 vgnd vpwr scs8hd_decap_4
Xmux_right_track_4.scs8hd_buf_4_0_ mux_right_track_4.mux_l4_in_0_/X _103_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D mux_left_track_1.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_224 vpwr vgnd scs8hd_fill_2
XFILLER_23_268 vpwr vgnd scs8hd_fill_2
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_33.mux_l3_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
Xmem_top_track_30.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_28.mux_l2_in_0_/S mux_top_track_30.mux_l1_in_0_/S
+ mem_top_track_30.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_18_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_59 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_10.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l3_in_0_/S
+ mem_left_track_17.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_40_80 vpwr vgnd scs8hd_fill_2
XFILLER_10_260 vgnd vpwr scs8hd_decap_12
X_098_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_32.mux_l1_in_1__A0 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2__S mux_right_track_16.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_179 vpwr vgnd scs8hd_fill_2
XFILLER_37_135 vpwr vgnd scs8hd_fill_2
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S mux_left_track_3.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_28_168 vpwr vgnd scs8hd_fill_2
XFILLER_28_135 vpwr vgnd scs8hd_fill_2
XFILLER_28_102 vgnd vpwr scs8hd_decap_3
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l1_in_1__A0 _043_/HI vgnd vpwr scs8hd_diode_2
XFILLER_19_102 vpwr vgnd scs8hd_fill_2
XFILLER_34_149 vpwr vgnd scs8hd_fill_2
XFILLER_19_81 vpwr vgnd scs8hd_fill_2
XFILLER_19_168 vpwr vgnd scs8hd_fill_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_25_149 vgnd vpwr scs8hd_decap_6
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_31_16 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_16.mux_l1_in_3_/S mux_right_track_16.mux_l2_in_0_/S
+ mem_right_track_16.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_4.mux_l1_in_5_ right_bottom_grid_pin_1_ right_top_grid_pin_49_ mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_5_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A0 mux_right_track_32.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_1__S mux_top_track_4.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_21_60 vgnd vpwr scs8hd_fill_1
XFILLER_21_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_30_174 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 mux_top_track_24.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D mux_left_track_3.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_59 vgnd vpwr scs8hd_decap_3
XFILLER_42_48 vgnd vpwr scs8hd_fill_1
XFILLER_21_130 vpwr vgnd scs8hd_fill_2
XFILLER_21_174 vgnd vpwr scs8hd_decap_6
XFILLER_29_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_12.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_12.mux_l1_in_0_/S mux_top_track_12.mux_l2_in_0_/S
+ mem_top_track_12.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_1.mux_l2_in_3__A1 left_bottom_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_37_37 vgnd vpwr scs8hd_decap_4
XFILLER_41_236 vpwr vgnd scs8hd_fill_2
XFILLER_41_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.scs8hd_buf_4_0__A mux_top_track_0.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A1 mux_left_track_3.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A1 mux_top_track_16.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_3.mux_l2_in_2_ left_top_grid_pin_47_ left_top_grid_pin_45_ mux_left_track_3.mux_l2_in_2_/S
+ mux_left_track_3.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XFILLER_27_70 vpwr vgnd scs8hd_fill_2
XFILLER_17_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l1_in_3__A0 _051_/HI vgnd vpwr scs8hd_diode_2
Xmem_top_track_38.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_38.mux_l1_in_1_/S mux_top_track_38.mux_l2_in_0_/S
+ mem_top_track_38.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_23_236 vpwr vgnd scs8hd_fill_2
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 chanx_right_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_14_225 vgnd vpwr scs8hd_fill_1
XFILLER_13_94 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_34.mux_l1_in_0__S mux_top_track_34.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_206 vpwr vgnd scs8hd_fill_2
XFILLER_20_239 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_2__S mux_left_track_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_28 vgnd vpwr scs8hd_fill_1
XFILLER_34_27 vpwr vgnd scs8hd_fill_2
XFILLER_11_239 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.scs8hd_dfxbp_1_3_ prog_clk mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l4_in_0_/S
+ mem_right_track_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_left_track_17.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_17.mux_l1_in_1_/S mux_left_track_17.mux_l2_in_0_/S
+ mem_left_track_17.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_4.mux_l2_in_3_ _065_/HI mux_right_track_4.mux_l1_in_6_/X mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_71 vgnd vpwr scs8hd_decap_4
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_097_ _097_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_10_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_32.mux_l1_in_1__A1 chany_top_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_6 vpwr vgnd scs8hd_fill_2
XFILLER_37_158 vgnd vpwr scs8hd_decap_4
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XFILLER_20_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D mux_left_track_3.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D mux_top_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_128 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_32.mux_l2_in_0__A0 _046_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_33_150 vgnd vpwr scs8hd_decap_3
Xmem_right_track_16.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_8.mux_l4_in_0_/S mux_right_track_16.mux_l1_in_3_/S
+ mem_right_track_16.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l1_in_4_ right_top_grid_pin_48_ right_top_grid_pin_47_ mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A1 mux_right_track_32.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vpwr vgnd scs8hd_fill_2
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_30_131 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l2_in_0__A1 mux_top_track_24.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__D mux_left_track_33.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S mux_right_track_4.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_153 vpwr vgnd scs8hd_fill_2
XFILLER_12_131 vpwr vgnd scs8hd_fill_2
Xmem_top_track_12.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_10.mux_l3_in_0_/S mux_top_track_12.mux_l1_in_0_/S
+ mem_top_track_12.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_32_71 vpwr vgnd scs8hd_fill_2
XFILLER_12_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A0 mux_left_track_17.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_256 vgnd vpwr scs8hd_decap_4
XFILLER_35_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_5__S mux_left_track_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_16 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.mux_l2_in_1_ left_top_grid_pin_43_ chanx_right_in[13] mux_left_track_3.mux_l2_in_2_/S
+ mux_left_track_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D mux_top_track_0.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_201 vgnd vpwr scs8hd_fill_1
XFILLER_17_223 vpwr vgnd scs8hd_fill_2
XFILLER_32_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_3__S mux_left_track_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_3__A0 left_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l1_in_3__A1 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmem_top_track_38.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_36.mux_l2_in_0_/S mux_top_track_38.mux_l1_in_1_/S
+ mem_top_track_38.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__D mux_left_track_5.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0__A1 mux_top_track_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.scs8hd_buf_4_0_ mux_top_track_8.mux_l3_in_0_/X _121_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_9_263 vgnd vpwr scs8hd_decap_12
XFILLER_9_252 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_18 vpwr vgnd scs8hd_fill_2
XFILLER_11_207 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l3_in_0_/S
+ mem_right_track_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_left_track_17.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_9.mux_l4_in_0_/S mux_left_track_17.mux_l1_in_1_/S
+ mem_left_track_17.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_4.mux_l2_in_2_ mux_right_track_4.mux_l1_in_5_/X mux_right_track_4.mux_l1_in_4_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_2__A0 mux_left_track_5.mux_l1_in_5_/X vgnd vpwr
+ scs8hd_diode_2
X_096_ chanx_left_in[8] chanx_right_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_37_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_19 vpwr vgnd scs8hd_fill_2
XFILLER_29_17 vpwr vgnd scs8hd_fill_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_19_148 vpwr vgnd scs8hd_fill_2
XFILLER_35_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l1_in_3__S mux_right_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l2_in_0__A1 mux_top_track_32.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_079_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_3_ _061_/HI chanx_left_in[17] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 chany_top_in[17] vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_3_ right_top_grid_pin_46_ right_top_grid_pin_45_ mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l3_in_1__A0 mux_left_track_5.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_107 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A0 mux_left_track_25.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_40 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_1_ _038_/HI chanx_left_in[13] mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D mux_top_track_0.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_187 vpwr vgnd scs8hd_fill_2
XFILLER_30_154 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vpwr vgnd scs8hd_fill_2
XFILLER_15_195 vpwr vgnd scs8hd_fill_2
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_38_210 vpwr vgnd scs8hd_fill_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_38_265 vgnd vpwr scs8hd_decap_8
XFILLER_29_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.scs8hd_buf_4_0__A mux_top_track_10.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_110 vgnd vpwr scs8hd_decap_8
XFILLER_12_154 vgnd vpwr scs8hd_decap_3
XFILLER_16_51 vpwr vgnd scs8hd_fill_2
XFILLER_16_73 vpwr vgnd scs8hd_fill_2
XFILLER_16_84 vgnd vpwr scs8hd_decap_4
XFILLER_32_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A1 mux_left_track_17.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_268 vpwr vgnd scs8hd_fill_2
XFILLER_35_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l4_in_0__A0 mux_left_track_5.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_8.scs8hd_buf_4_0__A mux_top_track_8.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_180 vgnd vpwr scs8hd_decap_3
XFILLER_26_224 vpwr vgnd scs8hd_fill_2
XFILLER_26_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_28.mux_l1_in_0__A0 chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_41_216 vgnd vpwr scs8hd_decap_4
XFILLER_26_257 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.mux_l2_in_0_ chanx_right_in[4] mux_left_track_3.mux_l1_in_0_/X mux_left_track_3.mux_l2_in_2_/S
+ mux_left_track_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_94 vpwr vgnd scs8hd_fill_2
XFILLER_27_50 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_track_24.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_24.mux_l2_in_1_/S mux_right_track_24.mux_l3_in_0_/S
+ mem_right_track_24.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_3__A1 left_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
Xmem_top_track_4.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l3_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_36.scs8hd_buf_4_0__A mux_top_track_36.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_19 vpwr vgnd scs8hd_fill_2
XFILLER_14_205 vpwr vgnd scs8hd_fill_2
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
XFILLER_14_249 vpwr vgnd scs8hd_fill_2
XFILLER_22_260 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_33.mux_l1_in_1__A0 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_38_71 vpwr vgnd scs8hd_fill_2
XFILLER_38_60 vpwr vgnd scs8hd_fill_2
XFILLER_20_219 vgnd vpwr scs8hd_fill_1
Xmux_top_track_14.scs8hd_buf_4_0_ mux_top_track_14.mux_l2_in_0_/X _118_/A vgnd vpwr
+ scs8hd_buf_1
Xmem_right_track_8.scs8hd_dfxbp_1_3_ prog_clk mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l4_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_275 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l2_in_1_/S
+ mem_right_track_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_16.mux_l2_in_1_ mux_right_track_16.mux_l1_in_3_/X mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_3__S mux_left_track_17.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_72 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_2__A1 mux_left_track_5.mux_l1_in_4_/X vgnd vpwr
+ scs8hd_diode_2
X_095_ chanx_left_in[9] chanx_right_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
XFILLER_27_7 vgnd vpwr scs8hd_fill_1
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_37_127 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_30.mux_l1_in_0__S mux_top_track_30.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l2_in_0__A0 mux_left_track_33.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D mux_left_track_9.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_160 vgnd vpwr scs8hd_decap_4
XFILLER_19_40 vpwr vgnd scs8hd_fill_2
XFILLER_19_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_83 vgnd vpwr scs8hd_decap_3
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
X_078_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_ chanx_left_in[8] right_top_grid_pin_47_ mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_174 vpwr vgnd scs8hd_fill_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 mux_right_track_2.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_2_ right_top_grid_pin_44_ right_top_grid_pin_43_ mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l3_in_1__A1 mux_left_track_5.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A1 mux_left_track_25.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_ chanx_right_in[13] top_left_grid_pin_38_ mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__D mux_left_track_17.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
Xmem_left_track_25.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l3_in_0_/S
+ mem_left_track_25.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_15_163 vpwr vgnd scs8hd_fill_2
XFILLER_15_174 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__D mux_right_track_32.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_36.mux_l1_in_0__A0 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_38_244 vgnd vpwr scs8hd_fill_1
Xmux_top_track_28.mux_l2_in_0_ _044_/HI mux_top_track_28.mux_l1_in_0_/X mux_top_track_28.mux_l2_in_0_/S
+ mux_top_track_28.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l3_in_0__S mux_top_track_8.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_22.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_2__A0 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_266 vpwr vgnd scs8hd_fill_2
XFILLER_12_144 vpwr vgnd scs8hd_fill_2
XFILLER_12_166 vpwr vgnd scs8hd_fill_2
XFILLER_16_63 vgnd vpwr scs8hd_decap_3
XFILLER_16_96 vpwr vgnd scs8hd_fill_2
Xmux_top_track_30.mux_l2_in_0_ _045_/HI mux_top_track_30.mux_l1_in_0_/X mux_top_track_30.mux_l2_in_0_/S
+ mux_top_track_30.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_35_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l4_in_0__A1 mux_left_track_5.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_6.mux_l1_in_3_ _051_/HI chanx_left_in[6] mux_top_track_6.mux_l1_in_0_/S
+ mux_top_track_6.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_269 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_28.mux_l1_in_0__A1 top_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_22.scs8hd_buf_4_0_ mux_top_track_22.mux_l2_in_0_/X _114_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_32_228 vgnd vpwr scs8hd_decap_3
XFILLER_32_206 vgnd vpwr scs8hd_decap_6
XFILLER_17_236 vpwr vgnd scs8hd_fill_2
XFILLER_40_250 vpwr vgnd scs8hd_fill_2
Xmem_right_track_24.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_24.mux_l1_in_1_/S mux_right_track_24.mux_l2_in_1_/S
+ mem_right_track_24.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D mux_top_track_4.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_4.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_4.mux_l1_in_1_/S mux_top_track_4.mux_l2_in_1_/S
+ mem_top_track_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_32.mux_l1_in_1__S mux_right_track_32.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_272 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l3_in_1__A0 mux_right_track_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_228 vpwr vgnd scs8hd_fill_2
XFILLER_13_86 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_33.mux_l1_in_1__A1 chany_top_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_5__S mux_right_track_4.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_8.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l3_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_22.mux_l2_in_0__S mux_top_track_22.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_221 vgnd vpwr scs8hd_decap_8
XFILLER_9_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_3__S mux_left_track_5.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_20.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_20.mux_l1_in_1_/S mux_top_track_20.mux_l2_in_0_/S
+ mem_top_track_20.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_3.mux_l4_in_0__S mux_left_track_3.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[6] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_track_0.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_38.mux_l2_in_0_/S mux_right_track_0.mux_l1_in_1_/S
+ mem_right_track_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_8.mux_l2_in_3__S mux_right_track_8.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_40_84 vpwr vgnd scs8hd_fill_2
X_094_ chanx_left_in[10] chanx_right_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0__S mux_top_track_16.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l3_in_0_ mux_top_track_6.mux_l2_in_1_/X mux_top_track_6.mux_l2_in_0_/X
+ mux_top_track_6.mux_l3_in_0_/S mux_top_track_6.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_0.mux_l4_in_0__A0 mux_right_track_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l3_in_1__S mux_left_track_9.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_139 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_33.mux_l2_in_0__A1 mux_left_track_33.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_183 vpwr vgnd scs8hd_fill_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_19_30 vgnd vpwr scs8hd_decap_4
XFILLER_42_120 vpwr vgnd scs8hd_fill_2
XFILLER_19_85 vpwr vgnd scs8hd_fill_2
XFILLER_19_106 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_38.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_42_153 vpwr vgnd scs8hd_fill_2
XFILLER_42_142 vgnd vpwr scs8hd_fill_1
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
X_077_ _077_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_32_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_142 vpwr vgnd scs8hd_fill_2
XFILLER_18_183 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l1_in_1_ right_top_grid_pin_43_ chany_top_in[17] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_1_ right_top_grid_pin_42_ chany_top_in[15] mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_6.mux_l2_in_1_ mux_top_track_6.mux_l1_in_3_/X mux_top_track_6.mux_l1_in_2_/X
+ mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_131 vpwr vgnd scs8hd_fill_2
XFILLER_24_142 vpwr vgnd scs8hd_fill_2
XFILLER_24_186 vpwr vgnd scs8hd_fill_2
XFILLER_21_53 vgnd vpwr scs8hd_decap_4
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_142 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_25.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_25.mux_l1_in_3_/S mux_left_track_25.mux_l2_in_0_/S
+ mem_left_track_25.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_6.scs8hd_dfxbp_1_1__D mux_top_track_6.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_36.mux_l1_in_0__A1 top_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_18.scs8hd_buf_4_0__A mux_top_track_18.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_223 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_2__A1 right_bottom_grid_pin_1_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_30.scs8hd_buf_4_0_ mux_top_track_30.mux_l2_in_0_/X _110_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_left_track_25.mux_l1_in_1__S mux_left_track_25.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_41 vpwr vgnd scs8hd_fill_2
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.mux_l2_in_1__S mux_right_track_24.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_6__A0 left_bottom_grid_pin_1_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.mux_l1_in_2_ chanx_right_in[11] chanx_right_in[6] mux_top_track_6.mux_l1_in_0_/S
+ mux_top_track_6.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_6.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D mux_right_track_8.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_74 vgnd vpwr scs8hd_fill_1
Xmem_right_track_24.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_16.mux_l3_in_0_/S mux_right_track_24.mux_l1_in_1_/S
+ mem_right_track_24.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
Xmux_top_track_28.mux_l1_in_0_ chanx_left_in[19] top_left_grid_pin_36_ mux_top_track_28.mux_l1_in_0_/S
+ mux_top_track_28.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
Xmem_top_track_4.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_2.mux_l3_in_0_/S mux_top_track_4.mux_l1_in_1_/S
+ mem_top_track_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_9.mux_l3_in_0__A0 mux_left_track_9.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l3_in_1__A1 mux_right_track_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_30.mux_l1_in_0_ chanx_left_in[15] top_left_grid_pin_37_ mux_top_track_30.mux_l1_in_0_/S
+ mux_top_track_30.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_218 vgnd vpwr scs8hd_decap_4
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_84 vpwr vgnd scs8hd_fill_2
XFILLER_38_40 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_251 vpwr vgnd scs8hd_fill_2
XANTENNA__125__A _125_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_20.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_18.mux_l2_in_0_/S mux_top_track_20.mux_l1_in_1_/S
+ mem_top_track_20.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l1_in_0__S mux_top_track_6.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_40_96 vpwr vgnd scs8hd_fill_2
XFILLER_40_41 vpwr vgnd scs8hd_fill_2
X_093_ _093_/A chanx_right_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l4_in_0__A1 mux_right_track_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_5.scs8hd_buf_4_0_ mux_left_track_5.mux_l4_in_0_/X _083_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D mux_top_track_6.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_162 vpwr vgnd scs8hd_fill_2
XFILLER_28_107 vgnd vpwr scs8hd_decap_3
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_184 vgnd vpwr scs8hd_decap_4
XFILLER_42_165 vgnd vpwr scs8hd_decap_3
X_076_ chanx_right_in[8] chanx_left_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_33_187 vgnd vpwr scs8hd_decap_3
XFILLER_33_121 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l1_in_0_ chany_top_in[10] chany_top_in[3] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_173 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[8] chany_top_in[1] mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_6.mux_l2_in_0_ mux_top_track_6.mux_l1_in_1_/X mux_top_track_6.mux_l1_in_0_/X
+ mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_10.mux_l1_in_0__A0 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_17.mux_l2_in_1__S mux_left_track_17.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_65 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_135 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
Xmem_left_track_25.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_17.mux_l3_in_0_/S mux_left_track_25.mux_l1_in_3_/S
+ mem_left_track_25.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_top_track_18.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_059_ _059_/HI _059_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_3 vgnd vpwr scs8hd_decap_4
XFILLER_38_257 vpwr vgnd scs8hd_fill_2
XFILLER_21_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_32_75 vpwr vgnd scs8hd_fill_2
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.scs8hd_dfxbp_1_2__D mux_top_track_10.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_2__S mux_top_track_0.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_7_172 vpwr vgnd scs8hd_fill_2
XFILLER_11_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_6__A1 left_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.mux_l1_in_1_ top_left_grid_pin_41_ top_left_grid_pin_39_ mux_top_track_6.mux_l1_in_0_/S
+ mux_top_track_6.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l1_in_3__S mux_top_track_6.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l3_in_0__S mux_top_track_4.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_17_227 vgnd vpwr scs8hd_decap_3
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l3_in_0__A1 mux_left_track_9.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
Xmem_top_track_28.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_28.mux_l1_in_0_/S mux_top_track_28.mux_l2_in_0_/S
+ mem_top_track_28.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_right_track_8.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_4.mux_l4_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_234 vpwr vgnd scs8hd_fill_2
XFILLER_13_263 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 mux_right_track_4.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_222 vgnd vpwr scs8hd_decap_12
XFILLER_24_21 vpwr vgnd scs8hd_fill_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_3
X_092_ chanx_left_in[12] chanx_right_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_37_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_38.mux_l1_in_1__A0 _049_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_3__A0 _062_/HI vgnd vpwr scs8hd_diode_2
Xmem_right_track_32.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_32.mux_l2_in_0_/S mux_right_track_32.mux_l3_in_0_/S
+ mem_right_track_32.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_1.mux_l2_in_3__S mux_left_track_1.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XFILLER_19_98 vpwr vgnd scs8hd_fill_2
XFILLER_35_97 vpwr vgnd scs8hd_fill_2
XFILLER_35_75 vpwr vgnd scs8hd_fill_2
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_27_130 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
X_075_ chanx_right_in[9] chanx_left_out[10] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_24.mux_l1_in_1__S mux_top_track_24.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_20.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_12.scs8hd_dfxbp_1_1__D mux_top_track_12.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l4_in_0__S mux_right_track_2.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_141 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_12.mux_l1_in_0__S mux_top_track_12.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_1__S mux_left_track_5.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_10.mux_l1_in_0__A1 top_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D mux_top_track_32.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_11 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l3_in_1__S mux_right_track_8.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_38.mux_l2_in_0__A0 mux_top_track_38.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_88 vpwr vgnd scs8hd_fill_2
XFILLER_30_158 vgnd vpwr scs8hd_decap_3
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.scs8hd_buf_4_0__A mux_left_track_5.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_058_ _058_/HI _058_/LO vgnd vpwr scs8hd_conb_1
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
XFILLER_38_247 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 top_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XFILLER_29_258 vpwr vgnd scs8hd_fill_2
XFILLER_29_236 vpwr vgnd scs8hd_fill_2
XFILLER_32_10 vpwr vgnd scs8hd_fill_2
XFILLER_16_55 vgnd vpwr scs8hd_decap_8
XFILLER_32_87 vgnd vpwr scs8hd_decap_3
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XFILLER_35_217 vpwr vgnd scs8hd_fill_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l1_in_0_ top_left_grid_pin_37_ top_left_grid_pin_35_ mux_top_track_6.mux_l1_in_0_/S
+ mux_top_track_6.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_228 vpwr vgnd scs8hd_fill_2
XFILLER_26_206 vpwr vgnd scs8hd_fill_2
XFILLER_34_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XFILLER_27_98 vgnd vpwr scs8hd_decap_4
XFILLER_27_54 vgnd vpwr scs8hd_decap_4
XFILLER_40_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l1_in_2__S mux_left_track_33.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_31_264 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D mux_top_track_38.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_14_209 vgnd vpwr scs8hd_decap_4
Xmem_left_track_33.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_33.mux_l2_in_0_/S ccff_tail
+ mem_left_track_33.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_64 vgnd vpwr scs8hd_decap_4
Xmem_top_track_28.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_24.mux_l2_in_0_/S mux_top_track_28.mux_l1_in_0_/S
+ mem_top_track_28.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_14.scs8hd_dfxbp_1_0__D mux_top_track_12.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 mux_right_track_4.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l3_in_0__S mux_top_track_10.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_39_194 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_34.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_34.scs8hd_dfxbp_1_0__D mux_top_track_32.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_10 vpwr vgnd scs8hd_fill_2
X_091_ chanx_left_in[13] chanx_right_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XFILLER_10_234 vgnd vpwr scs8hd_fill_1
XFILLER_24_44 vgnd vpwr scs8hd_decap_3
XFILLER_24_77 vpwr vgnd scs8hd_fill_2
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_38.mux_l1_in_1__A1 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_36_131 vpwr vgnd scs8hd_fill_2
Xmem_right_track_32.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_32.mux_l1_in_1_/S mux_right_track_32.mux_l2_in_0_/S
+ mem_right_track_32.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_2.mux_l2_in_3__A1 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_19_11 vpwr vgnd scs8hd_fill_2
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_42_178 vgnd vpwr scs8hd_decap_6
XFILLER_42_134 vgnd vpwr scs8hd_decap_8
XFILLER_35_43 vpwr vgnd scs8hd_fill_2
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_074_ chanx_right_in[10] chanx_left_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_2.mux_l1_in_0__S mux_top_track_2.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l3_in_0__A0 mux_top_track_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_112 vpwr vgnd scs8hd_fill_2
XFILLER_18_7 vpwr vgnd scs8hd_fill_2
XFILLER_18_186 vgnd vpwr scs8hd_fill_1
XFILLER_33_178 vgnd vpwr scs8hd_decap_3
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_4.scs8hd_buf_4_0__A mux_right_track_4.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_38.mux_l2_in_0__A1 mux_top_track_38.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_101 vpwr vgnd scs8hd_fill_2
XFILLER_30_104 vpwr vgnd scs8hd_fill_2
XFILLER_15_167 vpwr vgnd scs8hd_fill_2
X_057_ _057_/HI _057_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_38_215 vpwr vgnd scs8hd_fill_2
XFILLER_30_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__D mux_right_track_0.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_115 vgnd vpwr scs8hd_decap_4
XFILLER_21_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 top_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_37_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_12_148 vgnd vpwr scs8hd_decap_3
XFILLER_7_163 vpwr vgnd scs8hd_fill_2
X_109_ _109_/A chany_top_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XFILLER_19_270 vpwr vgnd scs8hd_fill_2
XFILLER_34_273 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l2_in_3_ _059_/HI left_bottom_grid_pin_1_ mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__070__A chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_40_210 vpwr vgnd scs8hd_fill_2
XFILLER_27_66 vpwr vgnd scs8hd_fill_2
XFILLER_27_33 vpwr vgnd scs8hd_fill_2
XFILLER_25_240 vpwr vgnd scs8hd_fill_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_40_254 vgnd vpwr scs8hd_decap_4
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l2_in_3_ _060_/HI chanx_left_in[12] mux_right_track_0.mux_l2_in_1_/S
+ mux_right_track_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_276 vgnd vpwr scs8hd_fill_1
XFILLER_16_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_33.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_33.mux_l1_in_0_/S mux_left_track_33.mux_l2_in_0_/S
+ mem_left_track_33.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_243 vpwr vgnd scs8hd_fill_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vpwr vgnd scs8hd_fill_2
XFILLER_38_10 vpwr vgnd scs8hd_fill_2
XFILLER_9_214 vpwr vgnd scs8hd_fill_2
XFILLER_13_210 vgnd vpwr scs8hd_decap_6
XFILLER_13_232 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_3__S mux_top_track_2.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l3_in_0__S mux_top_track_0.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.mux_l2_in_1__A1 top_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_1__A0 _036_/HI vgnd vpwr scs8hd_diode_2
XFILLER_39_184 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_6.mux_l2_in_1__S mux_top_track_6.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
X_090_ chanx_left_in[14] chanx_right_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_40_88 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
Xmem_top_track_10.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_10.mux_l2_in_0_/S mux_top_track_10.mux_l3_in_0_/S
+ mem_top_track_10.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S mux_left_track_9.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_154 vpwr vgnd scs8hd_fill_2
Xmem_right_track_32.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_24.mux_l3_in_0_/S mux_right_track_32.mux_l1_in_1_/S
+ mem_right_track_32.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D mux_right_track_2.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S mux_right_track_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_073_ _073_/A chanx_left_out[12] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A1 mux_top_track_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_14.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_146 vpwr vgnd scs8hd_fill_2
XFILLER_18_132 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_12.mux_l2_in_0__A0 mux_top_track_12.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.scs8hd_buf_4_0_ mux_right_track_0.mux_l4_in_0_/X _105_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_24_135 vpwr vgnd scs8hd_fill_2
XFILLER_24_146 vgnd vpwr scs8hd_decap_6
XFILLER_24_157 vgnd vpwr scs8hd_decap_8
XANTENNA__073__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_57 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_1_/S mux_left_track_9.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_146 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 chany_top_in[16] vgnd vpwr scs8hd_diode_2
X_125_ _125_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_30_149 vpwr vgnd scs8hd_fill_2
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_056_ _056_/HI _056_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_20.mux_l1_in_1__S mux_top_track_20.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_3__S mux_right_track_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__068__A chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_16_46 vgnd vpwr scs8hd_decap_3
XFILLER_16_68 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l3_in_1__S mux_left_track_1.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_45 vpwr vgnd scs8hd_fill_2
XFILLER_32_23 vgnd vpwr scs8hd_decap_4
XFILLER_12_105 vpwr vgnd scs8hd_fill_2
XFILLER_12_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_36.mux_l2_in_0__S mux_top_track_36.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__D mux_left_track_25.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_5__A0 right_bottom_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l3_in_1__S mux_right_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_108_ _108_/A chany_top_out[17] vgnd vpwr scs8hd_buf_2
X_039_ _039_/HI _039_/LO vgnd vpwr scs8hd_conb_1
Xmux_left_track_17.mux_l1_in_3_ _054_/HI left_top_grid_pin_47_ mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_241 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l2_in_2_ left_top_grid_pin_46_ left_top_grid_pin_42_ mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.mux_l2_in_2_ chanx_left_in[2] right_bottom_grid_pin_1_ mux_right_track_0.mux_l2_in_1_/S
+ mux_right_track_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_20.mux_l1_in_1__A0 _041_/HI vgnd vpwr scs8hd_diode_2
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
Xmux_top_track_12.mux_l2_in_0_ mux_top_track_12.mux_l1_in_1_/X mux_top_track_12.mux_l1_in_0_/X
+ mux_top_track_12.mux_l2_in_0_/S mux_top_track_12.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_28.scs8hd_buf_4_0_ mux_top_track_28.mux_l2_in_0_/X _111_/A vgnd vpwr
+ scs8hd_buf_1
Xmem_left_track_33.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_25.mux_l3_in_0_/S mux_left_track_33.mux_l1_in_0_/S
+ mem_left_track_33.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D mux_right_track_4.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_200 vpwr vgnd scs8hd_fill_2
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XANTENNA__081__A _081_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_88 vpwr vgnd scs8hd_fill_2
XFILLER_9_259 vpwr vgnd scs8hd_fill_2
XFILLER_9_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_18.scs8hd_dfxbp_1_1__D mux_top_track_18.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_1__A1 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_39_152 vpwr vgnd scs8hd_fill_2
XANTENNA__076__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_10_203 vgnd vpwr scs8hd_decap_8
XFILLER_40_45 vpwr vgnd scs8hd_fill_2
XFILLER_40_23 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S mux_left_track_17.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_20.mux_l2_in_0__A0 mux_top_track_20.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l2_in_0__S mux_left_track_33.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_10.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_10.mux_l1_in_0_/S mux_top_track_10.mux_l2_in_0_/S
+ mem_top_track_10.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_top_track_38.scs8hd_dfxbp_1_1__D mux_top_track_38.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.mux_l1_in_1_ _036_/HI chanx_left_in[10] mux_top_track_12.mux_l1_in_0_/S
+ mux_top_track_12.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_32.mux_l3_in_0__S mux_right_track_32.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_166 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_1__A0 top_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_103 vgnd vpwr scs8hd_decap_4
XFILLER_27_188 vgnd vpwr scs8hd_fill_1
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XFILLER_42_147 vgnd vpwr scs8hd_decap_4
X_072_ chanx_right_in[12] chanx_left_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_111 vpwr vgnd scs8hd_fill_2
XFILLER_18_177 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_12.mux_l2_in_0__A1 mux_top_track_12.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_191 vpwr vgnd scs8hd_fill_2
XFILLER_41_180 vgnd vpwr scs8hd_decap_3
Xmem_top_track_36.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_36.mux_l1_in_0_/S mux_top_track_36.mux_l2_in_0_/S
+ mem_top_track_36.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l2_in_1_ mux_left_track_17.mux_l1_in_3_/X mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_2.mux_l1_in_3__A0 _040_/HI vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_1_/S mux_left_track_9.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_36 vpwr vgnd scs8hd_fill_2
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_055_ _055_/HI _055_/LO vgnd vpwr scs8hd_conb_1
X_124_ _124_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_30_139 vgnd vpwr scs8hd_decap_3
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0__A0 mux_top_track_4.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_7 vgnd vpwr scs8hd_fill_1
XFILLER_38_206 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA__084__A _084_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_5__A1 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_107_ _107_/A chany_top_out[18] vgnd vpwr scs8hd_buf_2
X_038_ _038_/HI _038_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_176 vpwr vgnd scs8hd_fill_2
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_ left_top_grid_pin_43_ chanx_right_in[17] mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_36.scs8hd_buf_4_0_ mux_top_track_36.mux_l2_in_0_/X _107_/A vgnd vpwr
+ scs8hd_buf_1
Xmux_left_track_9.mux_l2_in_1_ chanx_right_in[16] chanx_right_in[6] mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__079__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_40_267 vgnd vpwr scs8hd_decap_8
XFILLER_25_264 vgnd vpwr scs8hd_decap_12
XFILLER_25_231 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.mux_l2_in_1_ right_top_grid_pin_48_ right_top_grid_pin_46_ mux_right_track_0.mux_l2_in_1_/S
+ mux_right_track_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_16_220 vpwr vgnd scs8hd_fill_2
XFILLER_16_264 vpwr vgnd scs8hd_fill_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_20.mux_l1_in_1__A1 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_31_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_234 vgnd vpwr scs8hd_decap_3
XFILLER_22_256 vpwr vgnd scs8hd_fill_2
XFILLER_22_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D mux_right_track_16.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XFILLER_38_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l3_in_0__S mux_left_track_25.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_238 vgnd vpwr scs8hd_decap_6
XFILLER_13_245 vgnd vpwr scs8hd_decap_4
XFILLER_13_267 vgnd vpwr scs8hd_decap_8
XFILLER_8_260 vgnd vpwr scs8hd_decap_12
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XFILLER_24_25 vpwr vgnd scs8hd_fill_2
XFILLER_40_68 vpwr vgnd scs8hd_fill_2
XANTENNA__092__A chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_20.mux_l2_in_0__A1 mux_top_track_20.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_10.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_8.mux_l3_in_0_/S mux_top_track_10.mux_l1_in_0_/S
+ mem_top_track_10.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_top_track_12.mux_l1_in_0_ chanx_right_in[10] top_left_grid_pin_36_ mux_top_track_12.mux_l1_in_0_/S
+ mux_top_track_12.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_80 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1__S mux_right_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_145 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S mux_top_track_24.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A1 top_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_36 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_35_79 vpwr vgnd scs8hd_fill_2
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_156 vpwr vgnd scs8hd_fill_2
XFILLER_27_134 vgnd vpwr scs8hd_fill_1
X_071_ chanx_right_in[13] chanx_left_out[14] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_2.mux_l2_in_1__S mux_top_track_2.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_145 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l1_in_0__S mux_left_track_9.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_104 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_36.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_34.mux_l2_in_0_/S mux_top_track_36.mux_l1_in_0_/S
+ mem_top_track_36.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 chany_top_in[11] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l1_in_3_ _040_/HI chanx_left_in[4] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_104 vpwr vgnd scs8hd_fill_2
Xmux_right_track_24.mux_l1_in_3_ _063_/HI chanx_left_in[18] mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_3__A1 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_15_159 vpwr vgnd scs8hd_fill_2
XFILLER_23_170 vpwr vgnd scs8hd_fill_2
X_123_ _123_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_054_ _054_/HI _054_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
Xmux_top_track_24.mux_l1_in_1_ _043_/HI chanx_left_in[18] mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A1 mux_top_track_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.scs8hd_buf_4_0_ mux_top_track_4.mux_l3_in_0_/X _123_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_16_7 vgnd vpwr scs8hd_decap_12
XFILLER_14_181 vpwr vgnd scs8hd_fill_2
XFILLER_37_240 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_162 vpwr vgnd scs8hd_fill_2
XFILLER_28_251 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_ chanx_right_in[8] chany_top_in[17] mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_106_ _106_/A chany_top_out[19] vgnd vpwr scs8hd_buf_2
X_037_ _037_/HI _037_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_155 vpwr vgnd scs8hd_fill_2
XFILLER_11_184 vgnd vpwr scs8hd_decap_4
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l2_in_0_ chany_top_in[18] mux_left_track_9.mux_l1_in_0_/X mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_34_232 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_2__A0 left_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XFILLER_27_58 vgnd vpwr scs8hd_fill_1
XFILLER_40_235 vgnd vpwr scs8hd_decap_4
XFILLER_25_276 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A chanx_left_in[9] vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l2_in_0__S mux_top_track_32.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_210 vgnd vpwr scs8hd_decap_4
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_17_80 vpwr vgnd scs8hd_fill_2
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_268 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l3_in_1__S mux_right_track_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_2__S mux_left_track_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_38_68 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D mux_right_track_8.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_38.mux_l1_in_1__S mux_top_track_38.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l3_in_1__A0 mux_left_track_1.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_5.scs8hd_dfxbp_1_3_ prog_clk mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l4_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_272 vgnd vpwr scs8hd_decap_3
Xmem_top_track_18.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_18.mux_l1_in_1_/S mux_top_track_18.mux_l2_in_0_/S
+ mem_top_track_18.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_top_track_12.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_1_ right_top_grid_pin_44_ right_top_grid_pin_42_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_238 vgnd vpwr scs8hd_decap_8
XFILLER_10_249 vgnd vpwr scs8hd_decap_8
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l1_in_3_/X mux_top_track_2.mux_l1_in_2_/X
+ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_24.mux_l2_in_1_ mux_right_track_24.mux_l1_in_3_/X mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_1_/S mux_right_track_24.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.scs8hd_buf_4_0__A mux_top_track_6.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_36_179 vpwr vgnd scs8hd_fill_2
XFILLER_36_135 vgnd vpwr scs8hd_decap_4
XFILLER_27_102 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l4_in_0__A0 mux_left_track_1.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_116 vpwr vgnd scs8hd_fill_2
XFILLER_35_47 vgnd vpwr scs8hd_decap_4
XFILLER_35_14 vpwr vgnd scs8hd_fill_2
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
X_070_ chanx_right_in[14] chanx_left_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_33_116 vgnd vpwr scs8hd_decap_3
XFILLER_18_102 vgnd vpwr scs8hd_decap_3
XFILLER_41_160 vpwr vgnd scs8hd_fill_2
XPHY_80 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_3__A0 _033_/HI vgnd vpwr scs8hd_diode_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_34.scs8hd_buf_4_0__A mux_top_track_34.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_91 vpwr vgnd scs8hd_fill_2
Xmem_top_track_2.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l3_in_0_/S
+ mem_top_track_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_2_ chanx_right_in[4] chanx_right_in[3] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_24.mux_l1_in_2_ chanx_left_in[9] right_top_grid_pin_48_ mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_32_182 vpwr vgnd scs8hd_fill_2
XFILLER_32_171 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D mux_right_track_32.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_20.scs8hd_dfxbp_1_1__D mux_top_track_20.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__098__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_30_108 vpwr vgnd scs8hd_fill_2
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
X_122_ _122_/A chany_top_out[3] vgnd vpwr scs8hd_buf_2
X_053_ _053_/HI _053_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 top_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_0__A1 mux_left_track_3.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[18] top_left_grid_pin_34_ mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_119 vgnd vpwr scs8hd_fill_1
XFILLER_29_219 vpwr vgnd scs8hd_fill_2
Xmux_top_track_36.mux_l2_in_0_ _048_/HI mux_top_track_36.mux_l1_in_0_/X mux_top_track_36.mux_l2_in_0_/S
+ mux_top_track_36.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_10.scs8hd_buf_4_0_ mux_top_track_10.mux_l3_in_0_/X _120_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
XFILLER_28_263 vpwr vgnd scs8hd_fill_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_11_141 vpwr vgnd scs8hd_fill_2
XFILLER_11_163 vgnd vpwr scs8hd_fill_1
X_105_ _105_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
Xmux_left_track_17.mux_l1_in_0_ chany_top_in[10] chany_top_in[3] mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_167 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
X_036_ _036_/HI _036_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_81 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l2_in_2__A1 left_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XFILLER_27_37 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_18.mux_l2_in_0__S mux_top_track_18.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_203 vgnd vpwr scs8hd_decap_6
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_6.mux_l1_in_2__A0 chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_38_36 vpwr vgnd scs8hd_fill_2
XFILLER_13_236 vgnd vpwr scs8hd_decap_8
XFILLER_9_229 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l3_in_1__A1 mux_left_track_1.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_ chany_top_in[11] chany_top_in[4] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_left_track_5.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l3_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_28_80 vpwr vgnd scs8hd_fill_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
Xmem_top_track_18.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_16.mux_l2_in_0_/S mux_top_track_18.mux_l1_in_1_/S
+ mem_top_track_18.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_199 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.mux_l1_in_0_ chany_top_in[13] chany_top_in[6] mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__D mux_left_track_1.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_49 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_32.mux_l1_in_0__A0 chanx_left_in[11] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_1_/S mux_right_track_24.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_22.scs8hd_dfxbp_1_0__D mux_top_track_20.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l2_in_1__A0 mux_top_track_6.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_81 vgnd vpwr scs8hd_decap_3
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_decap_4
XFILLER_39_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l4_in_0__A1 mux_left_track_1.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 top_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XFILLER_41_172 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_3__A1 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_3__S mux_right_track_16.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_2.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_2.mux_l1_in_1_/S mux_top_track_2.mux_l2_in_0_/S
+ mem_top_track_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_top_track_2.mux_l1_in_1_ top_left_grid_pin_41_ top_left_grid_pin_39_ mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_24.mux_l1_in_1_ right_top_grid_pin_44_ chany_top_in[18] mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__A0 mux_top_track_6.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_3__A0 _061_/HI vgnd vpwr scs8hd_diode_2
X_121_ _121_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
X_052_ _052_/HI _052_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_49 vgnd vpwr scs8hd_decap_3
XFILLER_20_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_2__S mux_top_track_4.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_120 vpwr vgnd scs8hd_fill_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
X_035_ _035_/HI _035_/LO vgnd vpwr scs8hd_conb_1
X_104_ _104_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XFILLER_21_7 vpwr vgnd scs8hd_fill_2
XFILLER_34_245 vgnd vpwr scs8hd_decap_3
Xmux_left_track_5.mux_l1_in_6_ left_bottom_grid_pin_1_ left_top_grid_pin_49_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_6_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D mux_left_track_3.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_36.mux_l1_in_0_ chanx_left_in[3] top_left_grid_pin_40_ mux_top_track_36.mux_l1_in_0_/S
+ mux_top_track_36.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_2__A1 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 left_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XFILLER_22_204 vgnd vpwr scs8hd_decap_8
XFILLER_13_259 vpwr vgnd scs8hd_fill_2
XFILLER_21_270 vpwr vgnd scs8hd_fill_2
Xmem_left_track_5.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_5.mux_l1_in_0_/S mux_left_track_5.mux_l2_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_16.scs8hd_buf_4_0__A mux_top_track_16.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_39_123 vpwr vgnd scs8hd_fill_2
XFILLER_24_17 vpwr vgnd scs8hd_fill_2
XFILLER_40_27 vpwr vgnd scs8hd_fill_2
XFILLER_10_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l1_in_0__A1 top_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l2_in_1__A1 mux_top_track_6.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_18.mux_l1_in_1__A0 _039_/HI vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vpwr vgnd scs8hd_fill_2
XFILLER_30_60 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A0 mux_left_track_5.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_22.mux_l1_in_0__S mux_top_track_22.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_2__S mux_right_track_2.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_3__S mux_left_track_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l1_in_3__A0 _063_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__S mux_left_track_3.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_126 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_18_137 vpwr vgnd scs8hd_fill_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_2.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_0.mux_l4_in_0_/S mux_top_track_2.mux_l1_in_1_/S
+ mem_top_track_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_9.mux_l2_in_1__S mux_left_track_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_3__A0 _056_/HI vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_37_ top_left_grid_pin_35_ mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_24.mux_l1_in_0_ chany_top_in[11] chany_top_in[4] mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_18.mux_l2_in_0__A0 mux_top_track_18.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A0 mux_left_track_5.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D mux_left_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__A1 mux_top_track_6.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_3__A1 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _120_/A chany_top_out[5] vgnd vpwr scs8hd_buf_2
X_051_ _051_/HI _051_/LO vgnd vpwr scs8hd_conb_1
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.scs8hd_buf_4_0__A mux_right_track_16.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_254 vpwr vgnd scs8hd_fill_2
XFILLER_37_243 vgnd vpwr scs8hd_fill_1
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_147 vgnd vpwr scs8hd_decap_8
XFILLER_11_154 vgnd vpwr scs8hd_decap_3
X_034_ _034_/HI _034_/LO vgnd vpwr scs8hd_conb_1
X_103_ _103_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_22_50 vpwr vgnd scs8hd_fill_2
XFILLER_34_257 vpwr vgnd scs8hd_fill_2
XFILLER_34_224 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_5_ left_top_grid_pin_48_ left_top_grid_pin_47_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_5_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_254 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.scs8hd_buf_4_0_ mux_left_track_1.mux_l4_in_0_/X _085_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__D mux_left_track_33.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_16_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_10.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_71 vpwr vgnd scs8hd_fill_2
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_268 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_24.mux_l1_in_1__S mux_right_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_6__S mux_left_track_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_38_27 vpwr vgnd scs8hd_fill_2
XFILLER_13_216 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D mux_top_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_5.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_3.mux_l4_in_0_/S mux_left_track_5.mux_l1_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_14.mux_l2_in_0__S mux_top_track_14.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_271 vgnd vpwr scs8hd_decap_4
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_39_179 vpwr vgnd scs8hd_fill_2
XFILLER_39_113 vpwr vgnd scs8hd_fill_2
XFILLER_24_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A1 mux_left_track_5.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_18.mux_l1_in_1__A1 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_39_70 vgnd vpwr scs8hd_decap_4
XFILLER_36_149 vgnd vpwr scs8hd_decap_4
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l1_in_3__A1 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.mux_l2_in_3__A1 left_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_108 vpwr vgnd scs8hd_fill_2
XFILLER_32_163 vpwr vgnd scs8hd_fill_2
XFILLER_17_193 vpwr vgnd scs8hd_fill_2
XFILLER_21_19 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l2_in_3_ _058_/HI mux_left_track_5.mux_l1_in_6_/X mux_left_track_5.mux_l2_in_0_/S
+ mux_left_track_5.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_18.mux_l2_in_0__A1 mux_top_track_18.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A1 mux_left_track_5.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_141 vgnd vpwr scs8hd_decap_4
XFILLER_23_174 vgnd vpwr scs8hd_decap_3
X_050_ _050_/HI _050_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vpwr vgnd scs8hd_fill_2
XFILLER_14_152 vgnd vpwr scs8hd_fill_1
XFILLER_14_185 vpwr vgnd scs8hd_fill_2
XFILLER_35_3 vpwr vgnd scs8hd_fill_2
XFILLER_37_266 vpwr vgnd scs8hd_fill_2
XFILLER_16_19 vgnd vpwr scs8hd_decap_12
XFILLER_32_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_20_122 vgnd vpwr scs8hd_fill_1
XFILLER_20_166 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_28_255 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1__S mux_left_track_17.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
X_033_ _033_/HI _033_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_159 vpwr vgnd scs8hd_fill_2
X_102_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D mux_top_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_222 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_1__S mux_right_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l1_in_4_ left_top_grid_pin_46_ left_top_grid_pin_45_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_266 vpwr vgnd scs8hd_fill_2
XFILLER_27_29 vpwr vgnd scs8hd_fill_2
XFILLER_25_214 vpwr vgnd scs8hd_fill_2
XFILLER_40_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_236 vpwr vgnd scs8hd_fill_2
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_16_247 vpwr vgnd scs8hd_fill_2
XFILLER_17_51 vpwr vgnd scs8hd_fill_2
XFILLER_17_62 vgnd vpwr scs8hd_decap_3
XFILLER_17_84 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S mux_left_track_5.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_239 vgnd vpwr scs8hd_decap_3
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_28.scs8hd_dfxbp_1_0__D mux_top_track_24.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_239 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A1 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.scs8hd_buf_4_0__A mux_left_track_3.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_34.mux_l2_in_0__A0 _047_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D mux_left_track_9.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__D mux_right_track_24.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_29_180 vgnd vpwr scs8hd_decap_3
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
XFILLER_35_18 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_3__A0 _054_/HI vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XPHY_84 vgnd vpwr scs8hd_decap_3
XFILLER_41_164 vpwr vgnd scs8hd_fill_2
XFILLER_41_142 vpwr vgnd scs8hd_fill_2
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_150 vgnd vpwr scs8hd_fill_1
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_40 vpwr vgnd scs8hd_fill_2
XFILLER_41_72 vgnd vpwr scs8hd_decap_4
XANTENNA__112__A top_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D mux_top_track_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_172 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_38.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_186 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.mux_l2_in_2_ mux_left_track_5.mux_l1_in_5_/X mux_left_track_5.mux_l1_in_4_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D mux_left_track_9.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
XFILLER_36_83 vgnd vpwr scs8hd_decap_3
XFILLER_36_50 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_3__S mux_right_track_4.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_223 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_1__S mux_left_track_5.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_3 vgnd vpwr scs8hd_fill_1
XFILLER_20_189 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XFILLER_28_267 vgnd vpwr scs8hd_decap_8
XFILLER_28_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_123 vpwr vgnd scs8hd_fill_2
X_101_ _101_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_22_85 vgnd vpwr scs8hd_fill_1
XFILLER_34_237 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_3_ left_top_grid_pin_44_ left_top_grid_pin_43_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_5__A0 left_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_33_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_215 vgnd vpwr scs8hd_fill_1
XFILLER_17_30 vgnd vpwr scs8hd_decap_6
XFILLER_24_270 vgnd vpwr scs8hd_decap_4
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_6.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.scs8hd_buf_4_0__A mux_right_track_2.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
XFILLER_28_84 vpwr vgnd scs8hd_fill_2
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_8_200 vgnd vpwr scs8hd_fill_1
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_34.mux_l2_in_0__A1 mux_top_track_34.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_148 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_32.mux_l1_in_2__S mux_right_track_32.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_3__A0 _055_/HI vgnd vpwr scs8hd_diode_2
XFILLER_38_181 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_41 vpwr vgnd scs8hd_fill_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_14_86 vpwr vgnd scs8hd_fill_2
XFILLER_39_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_6__S mux_right_track_4.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_192 vgnd vpwr scs8hd_decap_3
XFILLER_29_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l2_in_0__S mux_top_track_10.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_3
XFILLER_35_162 vpwr vgnd scs8hd_fill_2
XFILLER_35_151 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_3__A1 left_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XFILLER_26_162 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_107 vpwr vgnd scs8hd_fill_2
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_187 vpwr vgnd scs8hd_fill_2
XFILLER_41_176 vpwr vgnd scs8hd_fill_2
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l1_in_1__S mux_top_track_16.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_85 vgnd vpwr scs8hd_decap_4
XFILLER_41_62 vgnd vpwr scs8hd_fill_1
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_132 vpwr vgnd scs8hd_fill_2
XFILLER_17_151 vgnd vpwr scs8hd_decap_3
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_24.scs8hd_buf_4_0__A mux_top_track_24.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_98 vgnd vpwr scs8hd_decap_8
XFILLER_14_154 vpwr vgnd scs8hd_fill_2
XFILLER_42_6 vpwr vgnd scs8hd_fill_2
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_20_146 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l2_in_0__A1 mux_left_track_9.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_18.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
X_100_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
Xmux_top_track_16.scs8hd_buf_4_0_ mux_top_track_16.mux_l2_in_0_/X _117_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_34_205 vpwr vgnd scs8hd_fill_2
XFILLER_19_235 vgnd vpwr scs8hd_decap_3
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l1_in_2_ left_top_grid_pin_42_ chanx_right_in[14] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_25.mux_l1_in_3_ _055_/HI left_top_grid_pin_48_ mux_left_track_25.mux_l1_in_3_/S
+ mux_left_track_25.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_6.scs8hd_dfxbp_1_2__D mux_top_track_6.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_5__A1 left_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XFILLER_40_219 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l1_in_2__S mux_left_track_25.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_18.mux_l2_in_0_ mux_top_track_18.mux_l1_in_1_/X mux_top_track_18.mux_l1_in_0_/X
+ mux_top_track_18.mux_l2_in_0_/S mux_top_track_18.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_97 vpwr vgnd scs8hd_fill_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_263 vpwr vgnd scs8hd_fill_2
Xmux_top_track_20.mux_l2_in_0_ mux_top_track_20.mux_l1_in_1_/X mux_top_track_20.mux_l1_in_0_/X
+ mux_top_track_20.mux_l2_in_0_/S mux_top_track_20.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_24.scs8hd_buf_4_0__A mux_right_track_24.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_219 vpwr vgnd scs8hd_fill_2
XFILLER_21_230 vpwr vgnd scs8hd_fill_2
XFILLER_21_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D mux_right_track_16.mux_l1_in_3_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_28_63 vpwr vgnd scs8hd_fill_2
XFILLER_12_241 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_25.mux_l1_in_3__A1 left_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_39_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 mux_right_track_4.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_18.mux_l1_in_1_ _039_/HI chanx_left_in[14] mux_top_track_18.mux_l1_in_1_/S
+ mux_top_track_18.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_193 vpwr vgnd scs8hd_fill_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_86 vgnd vpwr scs8hd_decap_4
XFILLER_30_64 vpwr vgnd scs8hd_fill_2
XFILLER_36_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_10.scs8hd_dfxbp_1_0__D mux_top_track_8.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_20.mux_l1_in_1_ _041_/HI chanx_left_in[16] mux_top_track_20.mux_l1_in_1_/S
+ mux_top_track_20.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_38.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_30.scs8hd_dfxbp_1_0__D mux_top_track_28.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_2__A0 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l1_in_1__S mux_top_track_6.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_41_100 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_185 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XFILLER_41_199 vpwr vgnd scs8hd_fill_2
XFILLER_41_41 vpwr vgnd scs8hd_fill_2
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D mux_top_track_8.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_20.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_left_track_25.mux_l2_in_1_ mux_left_track_25.mux_l1_in_3_/X mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_166 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.scs8hd_buf_4_0_ mux_top_track_24.mux_l2_in_0_/X _113_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_36_30 vgnd vpwr scs8hd_fill_1
XFILLER_36_41 vgnd vpwr scs8hd_decap_3
XFILLER_14_144 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.mux_l3_in_1__A0 mux_right_track_2.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_258 vpwr vgnd scs8hd_fill_2
XFILLER_37_236 vgnd vpwr scs8hd_decap_4
XFILLER_20_158 vgnd vpwr scs8hd_fill_1
XFILLER_11_114 vgnd vpwr scs8hd_decap_4
XFILLER_22_32 vgnd vpwr scs8hd_decap_3
XFILLER_22_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_228 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_1_ chanx_right_in[5] chany_top_in[19] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_203 vpwr vgnd scs8hd_fill_2
XFILLER_19_258 vpwr vgnd scs8hd_fill_2
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
Xmux_left_track_25.mux_l1_in_2_ left_top_grid_pin_44_ chanx_right_in[18] mux_left_track_25.mux_l1_in_3_/S
+ mux_left_track_25.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 chany_top_in[15] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_1__S mux_left_track_1.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_36.mux_l1_in_0__S mux_top_track_36.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_206 vpwr vgnd scs8hd_fill_2
XFILLER_17_10 vpwr vgnd scs8hd_fill_2
XFILLER_17_43 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_75 vgnd vpwr scs8hd_decap_4
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_209 vgnd vpwr scs8hd_fill_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l4_in_0__A0 mux_right_track_2.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_3__S mux_top_track_0.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
Xmem_top_track_34.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_34.mux_l1_in_0_/S mux_top_track_34.mux_l2_in_0_/S
+ mem_top_track_34.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XFILLER_12_253 vpwr vgnd scs8hd_fill_2
XFILLER_39_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 top_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_18.mux_l1_in_0_ chanx_right_in[14] top_left_grid_pin_39_ mux_top_track_18.mux_l1_in_1_/S
+ mux_top_track_18.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_36.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_99 vpwr vgnd scs8hd_fill_2
XFILLER_30_10 vpwr vgnd scs8hd_fill_2
XFILLER_39_74 vgnd vpwr scs8hd_fill_1
Xmux_top_track_20.mux_l1_in_0_ chanx_right_in[16] top_left_grid_pin_40_ mux_top_track_20.mux_l1_in_1_/S
+ mux_top_track_20.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_38.mux_l1_in_0__A1 top_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XFILLER_35_175 vpwr vgnd scs8hd_fill_2
Xmux_top_track_32.mux_l2_in_0_ _046_/HI mux_top_track_32.mux_l1_in_0_/X mux_top_track_32.mux_l2_in_0_/S
+ mux_top_track_32.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_2__A1 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_32.scs8hd_buf_4_0_ mux_top_track_32.mux_l2_in_0_/X _109_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_41_123 vgnd vpwr scs8hd_decap_4
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_142 vpwr vgnd scs8hd_fill_2
XFILLER_26_131 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_41_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l1_in_0__S mux_left_track_33.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_178 vpwr vgnd scs8hd_fill_2
XFILLER_32_167 vpwr vgnd scs8hd_fill_2
XFILLER_32_145 vpwr vgnd scs8hd_fill_2
XFILLER_32_112 vpwr vgnd scs8hd_fill_2
XFILLER_17_197 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_101 vpwr vgnd scs8hd_fill_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l2_in_3__A0 _059_/HI vgnd vpwr scs8hd_diode_2
XFILLER_36_75 vpwr vgnd scs8hd_fill_2
XFILLER_14_112 vpwr vgnd scs8hd_fill_2
XFILLER_14_189 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_2.mux_l3_in_1__A1 mux_right_track_2.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_1__S mux_top_track_12.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XFILLER_20_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_28.mux_l2_in_0__S mux_top_track_28.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_159 vgnd vpwr scs8hd_decap_4
XFILLER_22_77 vpwr vgnd scs8hd_fill_2
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_ chany_top_in[12] chany_top_in[5] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_240 vgnd vpwr scs8hd_decap_4
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l4_in_0__S mux_left_track_9.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_25.mux_l1_in_1_ chanx_right_in[9] chany_top_in[16] mux_left_track_25.mux_l1_in_3_/S
+ mux_left_track_25.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_089_ _089_/A chanx_right_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
XFILLER_25_218 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S mux_top_track_8.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_55 vgnd vpwr scs8hd_decap_4
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l4_in_0__A1 mux_right_track_2.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_221 vpwr vgnd scs8hd_fill_2
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S mux_right_track_32.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_top_track_0.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l4_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
Xmem_top_track_34.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_32.mux_l2_in_0_/S mux_top_track_34.mux_l1_in_0_/S
+ mem_top_track_34.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_254 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_3
XFILLER_0_147 vgnd vpwr scs8hd_decap_8
XFILLER_28_76 vpwr vgnd scs8hd_fill_2
XFILLER_12_210 vgnd vpwr scs8hd_fill_1
XFILLER_8_203 vpwr vgnd scs8hd_fill_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_1_ _052_/HI chanx_left_in[8] mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_0.mux_l2_in_0__A1 mux_top_track_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_0.scs8hd_buf_4_0_ mux_top_track_0.mux_l4_in_0_/X _125_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D mux_right_track_0.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0__A0 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_38_140 vgnd vpwr scs8hd_fill_1
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_25.mux_l2_in_0__S mux_left_track_25.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_77 vpwr vgnd scs8hd_fill_2
Xmux_right_track_32.mux_l2_in_1_ _064_/HI mux_right_track_32.mux_l1_in_2_/X mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_86 vpwr vgnd scs8hd_fill_2
XFILLER_29_184 vgnd vpwr scs8hd_decap_3
XFILLER_29_162 vpwr vgnd scs8hd_fill_2
XFILLER_29_140 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_14.scs8hd_dfxbp_1_1__D mux_top_track_14.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l3_in_0__S mux_right_track_24.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_41_146 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_34.scs8hd_dfxbp_1_1__D mux_top_track_34.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_25_11 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_176 vgnd vpwr scs8hd_fill_1
XFILLER_32_124 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_track_32.mux_l1_in_2_ chanx_left_in[10] right_top_grid_pin_49_ mux_right_track_32.mux_l1_in_1_/S
+ mux_right_track_32.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_135 vgnd vpwr scs8hd_decap_4
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_3__A1 left_bottom_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_36_54 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_1__S mux_top_track_2.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
Xmem_left_track_3.scs8hd_dfxbp_1_3_ prog_clk mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l4_in_0_/S
+ mem_left_track_3.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_top_track_32.mux_l1_in_0_ chanx_left_in[11] top_left_grid_pin_38_ mux_top_track_32.mux_l1_in_0_/S
+ mux_top_track_32.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_top_track_16.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_16.mux_l1_in_1_/S mux_top_track_16.mux_l2_in_0_/S
+ mem_top_track_16.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_10.mux_l2_in_1__A0 _035_/HI vgnd vpwr scs8hd_diode_2
XFILLER_28_238 vpwr vgnd scs8hd_fill_2
XFILLER_11_127 vgnd vpwr scs8hd_fill_1
XFILLER_22_12 vpwr vgnd scs8hd_fill_2
XFILLER_22_23 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_4__A0 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_19_216 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.scs8hd_buf_4_0__A mux_top_track_4.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_25.mux_l1_in_0_ chany_top_in[9] chany_top_in[2] mux_left_track_25.mux_l1_in_3_/S
+ mux_left_track_25.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_40_6 vpwr vgnd scs8hd_fill_2
X_088_ chanx_left_in[16] chanx_right_out[17] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D mux_right_track_0.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_67 vpwr vgnd scs8hd_fill_2
XFILLER_24_241 vpwr vgnd scs8hd_fill_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_11 vpwr vgnd scs8hd_fill_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_274 vgnd vpwr scs8hd_fill_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_32.scs8hd_buf_4_0__A mux_top_track_32.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l3_in_0__A0 mux_top_track_10.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_255 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l3_in_1_/S
+ mem_top_track_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_20.mux_l1_in_0__A0 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D mux_top_track_14.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__A0 _065_/HI vgnd vpwr scs8hd_diode_2
XFILLER_21_266 vpwr vgnd scs8hd_fill_2
XANTENNA__071__A chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_28_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l3_in_0__S mux_left_track_17.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_36.scs8hd_dfxbp_1_0__D mux_top_track_34.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_4.scs8hd_dfxbp_1_3_ prog_clk mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l4_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_248 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l1_in_0__S mux_top_track_32.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_ chanx_right_in[15] mux_top_track_8.mux_l1_in_0_/X mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0__A1 top_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XANTENNA__066__A chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_38_185 vpwr vgnd scs8hd_fill_2
XFILLER_30_45 vgnd vpwr scs8hd_decap_4
XFILLER_30_23 vgnd vpwr scs8hd_decap_4
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_39_54 vpwr vgnd scs8hd_fill_2
XFILLER_39_10 vpwr vgnd scs8hd_fill_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_0_/S mux_right_track_32.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D mux_left_track_17.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l3_in_1__S mux_top_track_0.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_35_155 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 top_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_114 vpwr vgnd scs8hd_fill_2
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_32.scs8hd_buf_4_0__A mux_right_track_32.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.scs8hd_buf_4_0_ mux_left_track_17.mux_l3_in_0_/X _077_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__D mux_right_track_2.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_32.mux_l1_in_1_ right_top_grid_pin_45_ chany_top_in[19] mux_right_track_32.mux_l1_in_1_/S
+ mux_right_track_32.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_2__A0 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_36_88 vpwr vgnd scs8hd_fill_2
XFILLER_36_22 vpwr vgnd scs8hd_fill_2
XFILLER_14_158 vgnd vpwr scs8hd_decap_4
Xmem_left_track_3.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_3.mux_l2_in_2_/S mux_left_track_3.mux_l3_in_1_/S
+ mem_left_track_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_top_track_16.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_14.mux_l2_in_0_/S mux_top_track_16.mux_l1_in_1_/S
+ mem_top_track_16.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XFILLER_9_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l2_in_1__A1 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_28_206 vgnd vpwr scs8hd_decap_8
XANTENNA__074__A chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_106 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l1_in_4__A1 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XFILLER_42_253 vgnd vpwr scs8hd_decap_8
XFILLER_34_209 vgnd vpwr scs8hd_decap_3
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_087_ chanx_left_in[17] chanx_right_out[18] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_1__A0 mux_top_track_2.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_250 vpwr vgnd scs8hd_fill_2
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_34 vpwr vgnd scs8hd_fill_2
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_45 vpwr vgnd scs8hd_fill_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l3_in_0__A1 mux_top_track_10.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_0.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_0.mux_l1_in_0_/S mux_top_track_0.mux_l2_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_267 vgnd vpwr scs8hd_decap_8
XFILLER_30_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_20.mux_l1_in_0__A1 top_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l4_in_0__S mux_left_track_5.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__A1 mux_right_track_4.mux_l1_in_6_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_3__A0 _034_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_234 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l4_in_0__S mux_right_track_8.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_18.mux_l1_in_0__S mux_top_track_18.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
Xmem_right_track_4.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l3_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l3_in_0__A0 mux_top_track_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D mux_right_track_4.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_3_ _053_/HI left_bottom_grid_pin_1_ mux_left_track_1.mux_l2_in_2_/S
+ mux_left_track_1.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_39_66 vpwr vgnd scs8hd_fill_2
Xmux_left_track_25.scs8hd_buf_4_0_ mux_left_track_25.mux_l3_in_0_/X _073_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_29_197 vgnd vpwr scs8hd_decap_3
XFILLER_29_175 vgnd vpwr scs8hd_decap_3
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_35_101 vpwr vgnd scs8hd_fill_2
XFILLER_35_189 vgnd vpwr scs8hd_decap_3
XFILLER_35_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_26_189 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _077_/A vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_25_35 vgnd vpwr scs8hd_decap_3
XFILLER_41_45 vpwr vgnd scs8hd_fill_2
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_41_78 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[8] top_left_grid_pin_34_ mux_top_track_8.mux_l1_in_0_/S
+ mux_top_track_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_33.mux_l2_in_1__S mux_left_track_33.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_17_101 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_3
XFILLER_17_156 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_track_32.mux_l1_in_0_ chany_top_in[12] chany_top_in[5] mux_right_track_32.mux_l1_in_1_/S
+ mux_right_track_32.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_2__A1 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_39_270 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A0 left_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S mux_left_track_1.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_left_track_3.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_3.mux_l1_in_0_/S mux_left_track_3.mux_l2_in_2_/S
+ mem_left_track_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_14.scs8hd_buf_4_0__A mux_top_track_14.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA__090__A chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
XFILLER_42_265 vgnd vpwr scs8hd_decap_12
XFILLER_42_232 vpwr vgnd scs8hd_fill_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_086_ chanx_left_in[18] chanx_right_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XFILLER_26_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 mux_top_track_2.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_1__A0 left_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XFILLER_33_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_14.mux_l1_in_1__A0 _037_/HI vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_8.mux_l2_in_1_/S mux_top_track_8.mux_l3_in_0_/S
+ mem_top_track_8.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_17_14 vpwr vgnd scs8hd_fill_2
XFILLER_17_36 vgnd vpwr scs8hd_fill_1
XFILLER_17_47 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_top_track_0.mux_l1_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_15_210 vgnd vpwr scs8hd_fill_1
XFILLER_15_254 vpwr vgnd scs8hd_fill_2
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
X_069_ _069_/A chanx_left_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_24_3 vgnd vpwr scs8hd_decap_3
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_21_213 vpwr vgnd scs8hd_fill_2
Xmux_left_track_33.scs8hd_buf_4_0_ mux_left_track_33.mux_l3_in_0_/X _069_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_top_track_0.mux_l2_in_3__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0__S mux_top_track_8.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_4.mux_l1_in_3_/S mux_right_track_4.mux_l2_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_239 vgnd vpwr scs8hd_decap_6
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XFILLER_12_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0__A0 mux_top_track_14.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A0 mux_left_track_1.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l3_in_0__A1 mux_top_track_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_261 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.scs8hd_buf_4_0_ mux_right_track_2.mux_l4_in_0_/X _104_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_38_154 vpwr vgnd scs8hd_fill_2
XFILLER_38_132 vpwr vgnd scs8hd_fill_2
XFILLER_38_110 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l2_in_2_ left_top_grid_pin_48_ left_top_grid_pin_46_ mux_left_track_1.mux_l2_in_2_/S
+ mux_left_track_1.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D mux_right_track_24.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_12.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_41_138 vpwr vgnd scs8hd_fill_2
XFILLER_41_105 vpwr vgnd scs8hd_fill_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_157 vgnd vpwr scs8hd_decap_3
XFILLER_26_146 vgnd vpwr scs8hd_decap_4
XFILLER_26_135 vpwr vgnd scs8hd_fill_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_41_57 vpwr vgnd scs8hd_fill_2
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_149 vpwr vgnd scs8hd_fill_2
XFILLER_32_116 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A0 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_17_168 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0__S mux_left_track_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_3_ _062_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_1_/S
+ mux_right_track_2.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_17.scs8hd_buf_4_0__A mux_left_track_17.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XFILLER_39_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D mux_right_track_4.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_46 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_36_79 vpwr vgnd scs8hd_fill_2
XFILLER_14_116 vpwr vgnd scs8hd_fill_2
XFILLER_22_160 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_left_track_3.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_1.mux_l4_in_0_/S mux_left_track_3.mux_l1_in_0_/S
+ mem_left_track_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_22.mux_l1_in_1__A0 _042_/HI vgnd vpwr scs8hd_diode_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_160 vpwr vgnd scs8hd_fill_2
XFILLER_20_119 vgnd vpwr scs8hd_fill_1
XFILLER_9_197 vpwr vgnd scs8hd_fill_2
XFILLER_36_274 vgnd vpwr scs8hd_fill_1
XFILLER_36_252 vpwr vgnd scs8hd_fill_2
XFILLER_22_37 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l3_in_1__A0 mux_right_track_8.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__S mux_top_track_6.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_42_244 vgnd vpwr scs8hd_fill_1
XFILLER_10_130 vgnd vpwr scs8hd_decap_4
XFILLER_10_141 vgnd vpwr scs8hd_fill_1
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
X_085_ _085_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_33_266 vpwr vgnd scs8hd_fill_2
XFILLER_33_211 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_1__A1 mux_left_track_1.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_1__A1 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_8.mux_l1_in_0_/S mux_top_track_8.mux_l2_in_1_/S
+ mem_top_track_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_24_211 vgnd vpwr scs8hd_fill_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_22.mux_l2_in_0__A0 mux_top_track_22.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
XFILLER_15_266 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S mux_right_track_2.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_91 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_28.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_068_ chanx_right_in[16] chanx_left_out[17] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_6.mux_l1_in_1__A0 top_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l4_in_0__A0 mux_right_track_8.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_258 vpwr vgnd scs8hd_fill_2
XFILLER_28_36 vpwr vgnd scs8hd_fill_2
Xmem_top_track_24.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_24.mux_l1_in_1_/S mux_top_track_24.mux_l2_in_0_/S
+ mem_top_track_24.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__096__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_2.mux_l4_in_0_/S mux_right_track_4.mux_l1_in_3_/S
+ mem_right_track_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_207 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_14.mux_l2_in_0__A1 mux_top_track_14.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A1 mux_left_track_1.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_16.scs8hd_buf_4_0_ mux_right_track_16.mux_l3_in_0_/X _097_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_20.mux_l2_in_0__S mux_top_track_20.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_273 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l2_in_1_ left_top_grid_pin_44_ mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_2_/S mux_left_track_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_3.mux_l2_in_3__S mux_left_track_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_3__A0 _050_/HI vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l4_in_0__S mux_left_track_1.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__D mux_right_track_8.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_166 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_6.mux_l2_in_0__A0 mux_top_track_6.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l4_in_0__S mux_right_track_4.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0__S mux_top_track_14.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_20_70 vgnd vpwr scs8hd_decap_3
XFILLER_35_158 vpwr vgnd scs8hd_fill_2
XFILLER_35_114 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_41_14 vpwr vgnd scs8hd_fill_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_40_194 vgnd vpwr scs8hd_fill_1
XFILLER_32_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A1 right_bottom_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_15_70 vgnd vpwr scs8hd_fill_1
XFILLER_15_81 vgnd vpwr scs8hd_decap_4
Xmux_top_track_38.scs8hd_buf_4_0_ mux_top_track_38.mux_l2_in_0_/X _106_/A vgnd vpwr
+ scs8hd_buf_1
Xmux_left_track_1.mux_l1_in_2_ left_top_grid_pin_42_ chanx_right_in[12] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l2_in_2_ chanx_left_in[4] right_top_grid_pin_49_ mux_right_track_2.mux_l2_in_1_/S
+ mux_right_track_2.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2__A0 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_14_139 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.scs8hd_buf_4_0__A mux_left_track_1.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_183 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.mux_l2_in_0_ mux_top_track_14.mux_l1_in_1_/X mux_top_track_14.mux_l1_in_0_/X
+ mux_top_track_14.mux_l2_in_0_/S mux_top_track_14.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_22.mux_l1_in_1__A1 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_9_110 vgnd vpwr scs8hd_decap_3
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XFILLER_36_264 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D mux_left_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_30.mux_l2_in_0__A0 _045_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l3_in_1__A1 mux_right_track_8.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_264 vpwr vgnd scs8hd_fill_2
XFILLER_10_186 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_30.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_4
X_084_ _084_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_19_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A0 mux_right_track_16.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_14.mux_l1_in_1_ _037_/HI chanx_left_in[12] mux_top_track_14.mux_l1_in_0_/S
+ mux_top_track_14.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_top_track_8.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_6.mux_l3_in_0_/S mux_top_track_8.mux_l1_in_0_/S
+ mem_top_track_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_24_245 vpwr vgnd scs8hd_fill_2
XFILLER_33_15 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_22.mux_l2_in_0__A1 mux_top_track_22.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_24.scs8hd_buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _093_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_30_215 vgnd vpwr scs8hd_decap_4
XFILLER_30_204 vpwr vgnd scs8hd_fill_2
X_067_ chanx_right_in[17] chanx_left_out[18] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l4_in_0__A1 mux_right_track_8.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_1__A1 top_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
Xmem_top_track_24.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_22.mux_l2_in_0_/S mux_top_track_24.mux_l1_in_1_/S
+ mem_top_track_24.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_28_59 vpwr vgnd scs8hd_fill_2
XFILLER_12_204 vgnd vpwr scs8hd_decap_6
XFILLER_12_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l3_in_0__A0 mux_right_track_16.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
X_119_ _119_/A chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_38_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_2_/S mux_left_track_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_189 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_3__A1 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_58 vgnd vpwr scs8hd_decap_3
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.scs8hd_buf_4_0_ mux_top_track_6.mux_l3_in_0_/X _122_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_top_track_6.mux_l2_in_0__A1 mux_top_track_6.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 mux_left_track_5.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_18.mux_l1_in_0__A0 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_20_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_24.mux_l1_in_2__A0 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_26_104 vpwr vgnd scs8hd_fill_2
XFILLER_41_118 vpwr vgnd scs8hd_fill_2
XFILLER_34_192 vpwr vgnd scs8hd_fill_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D mux_left_track_1.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_22.scs8hd_dfxbp_1_1__D mux_top_track_22.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_184 vpwr vgnd scs8hd_fill_2
XFILLER_40_140 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_1_ chanx_right_in[2] chany_top_in[14] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_81 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.mux_l2_in_2__A0 left_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.scs8hd_buf_4_0__A mux_right_track_0.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l2_in_1_ right_top_grid_pin_47_ right_top_grid_pin_45_ mux_right_track_2.mux_l2_in_1_/S
+ mux_right_track_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_173 vgnd vpwr scs8hd_decap_4
XFILLER_39_240 vpwr vgnd scs8hd_fill_2
XFILLER_36_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2__A1 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A0 mux_right_track_24.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_173 vpwr vgnd scs8hd_fill_2
XFILLER_13_184 vgnd vpwr scs8hd_decap_3
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_36_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_30.mux_l2_in_0__A1 mux_top_track_30.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_32.scs8hd_buf_4_0_ mux_right_track_32.mux_l3_in_0_/X _089_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_27_210 vgnd vpwr scs8hd_decap_4
XFILLER_42_213 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_3.mux_l3_in_1__A0 mux_left_track_3.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_221 vgnd vpwr scs8hd_decap_3
XFILLER_10_154 vpwr vgnd scs8hd_fill_2
X_083_ _083_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_18_210 vpwr vgnd scs8hd_fill_2
XFILLER_18_254 vpwr vgnd scs8hd_fill_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A1 mux_right_track_16.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__S mux_left_track_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_14.mux_l1_in_0_ chanx_right_in[12] top_left_grid_pin_37_ mux_top_track_14.mux_l1_in_0_/S
+ mux_top_track_14.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_39 vpwr vgnd scs8hd_fill_2
XFILLER_33_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l3_in_0__A0 mux_right_track_24.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_3__S mux_top_track_4.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_30_238 vpwr vgnd scs8hd_fill_2
XFILLER_15_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l3_in_0__S mux_top_track_2.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
X_066_ chanx_right_in[18] chanx_left_out[19] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 chany_top_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_22.scs8hd_buf_4_0__A mux_top_track_22.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l4_in_0__A0 mux_left_track_3.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__D mux_left_track_3.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_1__S mux_top_track_8.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D mux_top_track_22.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__A1 mux_right_track_16.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_3_ _050_/HI chanx_left_in[5] mux_top_track_4.mux_l1_in_1_/S
+ mux_top_track_4.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
X_118_ _118_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
X_049_ _049_/HI _049_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_32.mux_l1_in_2__A0 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_38_102 vpwr vgnd scs8hd_fill_2
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail mux_left_track_33.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_0__A1 mux_left_track_5.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_18.mux_l1_in_0__A1 top_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XFILLER_29_70 vgnd vpwr scs8hd_decap_3
XFILLER_35_127 vgnd vpwr scs8hd_decap_3
Xmux_top_track_12.scs8hd_buf_4_0_ mux_top_track_12.mux_l2_in_0_/X _119_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_right_track_24.mux_l1_in_2__A1 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__D mux_left_track_25.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_160 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_32.mux_l2_in_1__A0 _064_/HI vgnd vpwr scs8hd_diode_2
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XFILLER_40_130 vpwr vgnd scs8hd_fill_2
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_ chany_top_in[7] chany_top_in[0] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_2__A1 left_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_22.mux_l1_in_1__S mux_top_track_22.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_3__S mux_right_track_2.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_4__S mux_left_track_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.scs8hd_buf_4_0__A mux_left_track_9.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l1_in_0__S mux_top_track_10.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l4_in_0__S mux_right_track_0.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_3.mux_l3_in_1__S mux_left_track_3.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_274 vgnd vpwr scs8hd_decap_3
Xmux_left_track_33.mux_l2_in_1_ _057_/HI mux_left_track_33.mux_l1_in_2_/X mux_left_track_33.mux_l2_in_0_/S
+ mux_left_track_33.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_38.mux_l2_in_0__S mux_top_track_38.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_163 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_24.mux_l2_in_1__A1 mux_right_track_24.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_2__S mux_left_track_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_32.mux_l3_in_0__A0 mux_right_track_32.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D mux_left_track_5.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_247 vgnd vpwr scs8hd_fill_1
XFILLER_42_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l3_in_1__A1 mux_left_track_3.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_082_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
Xmux_right_track_2.mux_l1_in_1_ right_top_grid_pin_43_ chany_top_in[14] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_258 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l1_in_3_/X mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_33.mux_l1_in_2_ left_top_grid_pin_49_ left_top_grid_pin_45_ mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_34.mux_l1_in_0__A0 chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_17_18 vgnd vpwr scs8hd_decap_12
XFILLER_33_28 vgnd vpwr scs8hd_decap_4
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_203 vpwr vgnd scs8hd_fill_2
XFILLER_24_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.mux_l3_in_0__A1 mux_right_track_24.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_1__A0 _052_/HI vgnd vpwr scs8hd_diode_2
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
XFILLER_15_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.scs8hd_buf_4_0__A mux_left_track_25.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
X_065_ _065_/HI _065_/LO vgnd vpwr scs8hd_conb_1
XFILLER_17_6 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_21_217 vpwr vgnd scs8hd_fill_2
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l4_in_0__A1 mux_left_track_3.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_228 vgnd vpwr scs8hd_decap_4
Xmux_top_track_4.mux_l1_in_2_ chanx_right_in[7] chanx_right_in[5] mux_top_track_4.mux_l1_in_1_/S
+ mux_top_track_4.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_83 vpwr vgnd scs8hd_fill_2
X_117_ _117_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
Xmux_top_track_20.scs8hd_buf_4_0_ mux_top_track_20.mux_l2_in_0_/X _115_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_34_93 vpwr vgnd scs8hd_fill_2
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.mux_l1_in_2__S mux_right_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l1_in_2__A1 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
X_048_ _048_/HI _048_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_158 vpwr vgnd scs8hd_fill_2
XFILLER_38_136 vpwr vgnd scs8hd_fill_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l3_in_0__A0 mux_top_track_8.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_29 vpwr vgnd scs8hd_fill_2
XFILLER_39_27 vpwr vgnd scs8hd_fill_2
XFILLER_29_136 vgnd vpwr scs8hd_decap_4
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_37_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
Xmux_top_track_38.mux_l2_in_0_ mux_top_track_38.mux_l1_in_1_/X mux_top_track_38.mux_l1_in_0_/X
+ mux_top_track_38.mux_l2_in_0_/S mux_top_track_38.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_62 vpwr vgnd scs8hd_fill_2
XFILLER_20_84 vgnd vpwr scs8hd_decap_4
XFILLER_29_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__D mux_top_track_0.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_191 vgnd vpwr scs8hd_decap_4
XFILLER_41_109 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2__A0 left_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l2_in_1__A1 mux_right_track_32.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.scs8hd_buf_4_0__A mux_right_track_8.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_15_62 vgnd vpwr scs8hd_decap_8
XFILLER_15_73 vpwr vgnd scs8hd_fill_2
XFILLER_17_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 chany_top_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__S mux_top_track_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA__102__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
Xmem_top_track_32.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_32.mux_l1_in_0_/S mux_top_track_32.mux_l2_in_0_/S
+ mem_top_track_32.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_142 vpwr vgnd scs8hd_fill_2
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_0_/S mux_left_track_33.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_38.mux_l1_in_1_ _049_/HI chanx_left_in[1] mux_top_track_38.mux_l1_in_1_/S
+ mux_top_track_38.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_71 vpwr vgnd scs8hd_fill_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A0 mux_left_track_17.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_36_256 vpwr vgnd scs8hd_fill_2
XFILLER_36_223 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_32.mux_l3_in_0__A1 mux_right_track_32.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_134 vgnd vpwr scs8hd_fill_1
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
X_081_ _081_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_37_71 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[7] chany_top_in[0] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_223 vpwr vgnd scs8hd_fill_2
XFILLER_18_267 vgnd vpwr scs8hd_decap_8
XFILLER_41_270 vgnd vpwr scs8hd_decap_6
Xmux_left_track_33.mux_l1_in_1_ chanx_right_in[10] chany_top_in[15] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_4__A0 left_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_34.mux_l1_in_0__A1 top_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2__S mux_left_track_17.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l3_in_0__A0 mux_left_track_17.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_40 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vpwr vgnd scs8hd_fill_2
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
X_064_ _064_/HI _064_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D mux_top_track_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_1__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D mux_left_track_5.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_1_ top_left_grid_pin_40_ top_left_grid_pin_38_ mux_top_track_4.mux_l1_in_1_/S
+ mux_top_track_4.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_116_ _116_/A chany_top_out[9] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_3__A0 _058_/HI vgnd vpwr scs8hd_diode_2
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_28.scs8hd_dfxbp_1_1__D mux_top_track_28.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
X_047_ _047_/HI _047_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_25.mux_l1_in_2__A0 left_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l3_in_0__A1 mux_top_track_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_1__S mux_top_track_4.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.scs8hd_buf_4_0_ mux_right_track_8.mux_l4_in_0_/X _101_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D mux_left_track_17.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__D mux_right_track_32.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_41_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2__A1 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vpwr vgnd scs8hd_fill_2
XFILLER_25_162 vpwr vgnd scs8hd_fill_2
XFILLER_15_85 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l2_in_1__A0 mux_left_track_25.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_40 vpwr vgnd scs8hd_fill_2
Xmem_top_track_32.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_30.mux_l2_in_0_/S mux_top_track_32.mux_l1_in_0_/S
+ mem_top_track_32.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
XFILLER_31_110 vpwr vgnd scs8hd_fill_2
XFILLER_16_173 vpwr vgnd scs8hd_fill_2
XFILLER_31_165 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_3.scs8hd_buf_4_0_ mux_left_track_3.mux_l4_in_0_/X _084_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_39_254 vgnd vpwr scs8hd_decap_4
XFILLER_39_210 vgnd vpwr scs8hd_decap_3
XFILLER_36_18 vpwr vgnd scs8hd_fill_2
Xmux_top_track_38.mux_l1_in_0_ chanx_right_in[0] top_left_grid_pin_41_ mux_top_track_38.mux_l1_in_1_/S
+ mux_top_track_38.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_22_132 vpwr vgnd scs8hd_fill_2
XFILLER_22_154 vgnd vpwr scs8hd_decap_6
XFILLER_22_187 vpwr vgnd scs8hd_fill_2
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XFILLER_26_40 vgnd vpwr scs8hd_fill_1
XFILLER_42_94 vpwr vgnd scs8hd_fill_2
XFILLER_9_158 vpwr vgnd scs8hd_fill_2
XFILLER_9_147 vpwr vgnd scs8hd_fill_2
XFILLER_13_110 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D mux_top_track_4.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A1 mux_left_track_17.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_235 vpwr vgnd scs8hd_fill_2
XFILLER_36_268 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_32.mux_l1_in_0__S mux_right_track_32.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A0 mux_left_track_25.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_268 vgnd vpwr scs8hd_decap_8
XFILLER_27_235 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__D mux_left_track_9.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
X_080_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_34.mux_l2_in_0__S mux_top_track_34.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_4__S mux_right_track_4.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_94 vpwr vgnd scs8hd_fill_2
XFILLER_33_238 vgnd vpwr scs8hd_decap_4
XFILLER_33_205 vgnd vpwr scs8hd_decap_4
Xmux_left_track_33.mux_l1_in_0_ chany_top_in[8] chany_top_in[1] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l3_in_1__S mux_right_track_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_2__S mux_left_track_5.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_4__A1 left_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_2__S mux_right_track_8.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_208 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_17.mux_l3_in_0__A1 mux_left_track_17.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_28.mux_l1_in_0__S mux_top_track_28.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_063_ _063_/HI _063_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l1_in_2__A0 left_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l3_in_0__S mux_left_track_9.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_28.mux_l2_in_0__A0 _044_/HI vgnd vpwr scs8hd_diode_2
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_36_ top_left_grid_pin_34_ mux_top_track_4.mux_l1_in_1_/S
+ mux_top_track_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_84 vpwr vgnd scs8hd_fill_2
XFILLER_34_73 vpwr vgnd scs8hd_fill_2
XFILLER_34_51 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.scs8hd_dfxbp_1_3_ prog_clk mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l4_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
X_115_ _115_/A chany_top_out[10] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_5.mux_l2_in_3__A1 mux_left_track_5.mux_l1_in_6_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_245 vpwr vgnd scs8hd_fill_2
XFILLER_11_252 vgnd vpwr scs8hd_decap_4
XFILLER_11_263 vpwr vgnd scs8hd_fill_2
X_046_ _046_/HI _046_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__121__A _121_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_14.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_14.mux_l1_in_0_/S mux_top_track_14.mux_l2_in_0_/S
+ mem_top_track_14.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_6 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_25.mux_l1_in_2__A1 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_38_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_33.mux_l2_in_1__A0 _057_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.scs8hd_buf_4_0__A mux_top_track_2.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_6.scs8hd_dfxbp_1_0__D mux_top_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_108 vpwr vgnd scs8hd_fill_2
XFILLER_19_193 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XFILLER_40_188 vgnd vpwr scs8hd_decap_6
XFILLER_40_100 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_25.mux_l2_in_1__A1 mux_left_track_25.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__S mux_left_track_25.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_30.scs8hd_buf_4_0__A mux_top_track_30.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_273 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l3_in_0__A0 mux_left_track_33.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_22.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l2_in_1__S mux_top_track_10.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
.ends

