version https://git-lfs.github.com/spec/v1
oid sha256:5ea86ad5b43ac7b2709cf0c8cf84478705705f49ef25dba6b5ca1a9f654fbc3a
size 36467042
