//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog netlist for pre-configured FPGA fabric by design: top
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Nov 24 18:04:19 2020
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

module top_top_formal_verification (
input [0:0] a_fm,
input [0:0] b_fm,
output [0:0] out_c_fm);

// ----- Local wires for FPGA fabric -----
wire [0:0] prog_clk;
wire [0:0] Test_en;
wire [0:0] IO_ISOL_N;
wire [0:0] clk;
wire [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_IN;
wire [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT;
wire [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR;
wire [0:0] ccff_head;
wire [0:0] ccff_tail;

// ----- FPGA top-level module to be capsulated -----
	fpga_core U0_formal_verification (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.IO_ISOL_N(IO_ISOL_N[0]),
		.clk(clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0:95]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0:95]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0:95]),
		.ccff_head(ccff_head[0]),
		.ccff_tail(ccff_tail[0]),
		.sc_head(sc_head[0]),
		.sc_tail(sc_tail[0])
		);

// ----- Begin Connect Global ports of FPGA top module -----
	assign Test_en[0] = 1'b0;
	assign prog_clk[0] = 1'b0;
	assign IO_ISOL_N[0] = 1'b1;
// ----- End Connect Global ports of FPGA top module -----

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input a is mapped to FPGA IOPAD gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4] -----
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4] = a_fm[0];

// ----- Blif Benchmark input b is mapped to FPGA IOPAD gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3] -----
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3] = b_fm[0];

// ----- Blif Benchmark output out:c is mapped to FPGA IOPAD gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] -----
	assign out_c_fm[0] = gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95] = 1'b0;

	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95] = 1'b0;

// ----- Begin load bitstream to configuration memories -----
`ifdef ICARUS_SIMULATOR
// ----- Begin assign bitstream to configuration memories -----
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = 17'b00000000110000001;
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = 2'b01;
	assign U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	// assign U0_formal_verification.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_top_top_2__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_top_top_3__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_top_top_4__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_top_top_5__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_top_top_6__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b0;
	// assign U0_formal_verification.grid_io_top_top_7__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_top_top_8__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_right_right_9__7_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_right_right_9__6_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_right_right_9__5_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_right_right_9__4_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_right_right_9__3_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_right_right_9__2_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_right_right_9__1_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_left_left_0__2_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_left_left_0__3_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_left_left_0__4_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_left_left_0__5_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_left_left_0__6_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_left_left_0__7_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	// assign U0_formal_verification.grid_io_left_left_0__8_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__4_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__5_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__6_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__7_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__8_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__4_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__5_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__7_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__8_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__4_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__5_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__7_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__8_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__4_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__5_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__7_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_right_track_4.mem_out[0:3] = {4{1'b1}};
	assign U0_formal_verification.sb_3__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_3__8_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__1_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__2_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__3_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__4_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__5_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__7_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_right_track_4.mem_out[0:3] = {4{1'b1}};
	assign U0_formal_verification.sb_4__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_4__8_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__1_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__2_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__3_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__4_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__5_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_top_track_4.mem_out[0:4] = 5'b00101;
	assign U0_formal_verification.sb_5__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__7_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_right_track_8.mem_out[0:3] = 4'b0101;
	assign U0_formal_verification.sb_5__8_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_1.mem_out[0:2] = 3'b100;
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_3.mem_out[0:2] = 3'b010;
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_5__8_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__1_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__2_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__3_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__4_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__5_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__7_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_6__8_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__1_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__2_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__3_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__4_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__5_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__7_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_7__8_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__0_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__1_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__2_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__3_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__4_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__5_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__6_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__7_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_8__8_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_3__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__0_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__0_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__0_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__0_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__0_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_4__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__0_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__0_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__0_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__0_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__0_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_5__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__0_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__0_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__0_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__0_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__0_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_bottom_ipin_0.mem_out[0:3] = 4'b1101;
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_6__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__0_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__0_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__0_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__0_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__0_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_7__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__0_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__0_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__0_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__0_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__0_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_8__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_3__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_4__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_12.mem_out[0:3] = 4'b0111;
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_13.mem_out[0:3] = 4'b0111;
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_5__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_6__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_7__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_8__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
// ----- End assign bitstream to configuration memories -----
`else
// ----- Begin deposit bitstream to configuration memories -----
initial begin
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_4__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], 17'b00000000110000001);
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.grid_clb_5__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_6__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_7__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__1_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__2_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__3_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__4_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__5_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__6_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__7_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_0.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_1.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_2.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_3.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_4.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_5.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_6.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.ltile_fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_8__8_.ltile_clb_mode__0.ltile_fle_7.ltile_fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_top_2__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_top_3__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_top_4__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_top_5__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_top_6__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_top_7__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_top_8__9_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_right_9__7_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_right_9__6_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_right_9__5_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_right_9__4_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_right_9__3_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_right_9__2_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_right_9__1_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_left_0__2_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_left_0__3_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_left_0__4_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_left_0__5_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_left_0__6_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_left_0__7_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_left_0__8_.logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_top_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_12.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_14.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_top_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_12.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_14.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_right_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__4_.mem_bottom_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_top_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_12.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_14.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_right_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__5_.mem_bottom_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_top_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_12.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_14.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_right_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__6_.mem_bottom_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_top_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_12.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_14.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_right_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__7_.mem_bottom_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_right_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_bottom_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_bottom_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_bottom_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__8_.mem_bottom_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__4_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__5_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__6_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__7_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_bottom_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__8_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__4_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__5_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__6_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__7_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_bottom_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__8_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__4_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__5_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__6_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__7_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_right_track_4.mem_out[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_3__8_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_bottom_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_3__8_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_top_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__0_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__1_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__2_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__3_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__4_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__5_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__6_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__7_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_right_track_4.mem_out[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_4__8_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_bottom_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_4__8_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_top_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__0_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__1_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__2_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__3_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__4_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__5_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__6_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_top_track_4.mem_out[0:4], 5'b00101);
	$deposit(U0_formal_verification.sb_5__7_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__7_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_right_track_8.mem_out[0:3], 4'b0101);
	$deposit(U0_formal_verification.sb_5__8_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_1.mem_out[0:2], 3'b100);
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_3.mem_out[0:2], 3'b010);
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_bottom_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_5__8_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_top_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__0_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__1_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__2_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__3_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__4_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__5_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__6_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__7_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_bottom_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_6__8_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_top_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__0_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__1_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__2_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__3_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__4_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__5_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__6_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__7_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_bottom_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_7__8_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_top_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__0_.mem_left_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_top_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_bottom_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_13.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_15.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__1_.mem_left_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_top_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_bottom_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_13.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_15.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__2_.mem_left_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_top_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_bottom_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_13.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_15.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__3_.mem_left_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_top_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_bottom_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_13.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_15.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__4_.mem_left_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_top_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_bottom_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_13.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_15.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__5_.mem_left_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_top_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_bottom_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_13.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_15.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__6_.mem_left_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_top_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_bottom_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_13.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_15.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__7_.mem_left_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_bottom_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_8__8_.mem_left_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__4_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__5_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__6_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__7_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__8_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__4_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__5_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__6_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__7_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__8_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__4_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__5_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__6_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__7_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_3__8_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__0_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__0_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__0_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__0_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__0_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__1_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__2_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__3_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__4_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__5_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__6_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__7_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_4__8_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__0_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__0_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__0_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__0_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__0_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__0_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__0_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__0_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__0_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__1_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__2_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__3_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__4_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__5_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__6_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__7_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_5__8_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__0_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__0_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__0_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__0_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__0_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__0_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__0_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__0_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__0_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__1_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__2_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__3_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__4_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__5_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__6_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__7_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_bottom_ipin_0.mem_out[0:3], 4'b1101);
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_6__8_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__0_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__0_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__0_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__0_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__0_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__0_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__0_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__0_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__0_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__1_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__2_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__3_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__4_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__5_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__6_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__7_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_7__8_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__0_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__0_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__0_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__0_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__0_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__0_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__0_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__0_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__0_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__1_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__2_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__3_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__4_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__5_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__6_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__7_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_8__8_.mem_top_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__7_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__8_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__4_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__5_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__6_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__7_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__8_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__4_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__5_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__6_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__7_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__8_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__4_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__5_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__6_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__7_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_3__8_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__1_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__2_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__3_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__4_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__5_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__6_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__7_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_4__8_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__1_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__2_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__3_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__4_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__5_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__6_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__7_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_12.mem_out[0:3], 4'b0111);
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_13.mem_out[0:3], 4'b0111);
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_5__8_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__1_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__2_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__3_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__4_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__5_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__6_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__7_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_6__8_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__1_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__2_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__3_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__4_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__5_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__6_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__7_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_7__8_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__1_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__2_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__3_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__4_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__5_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__6_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__7_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_8__8_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
end
// ----- End deposit bitstream to configuration memories -----
`endif
// ----- End load bitstream to configuration memories -----
endmodule
// ----- END Verilog module for top_top_formal_verification -----

