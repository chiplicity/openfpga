VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 137.630 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.940 0.000 24.220 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.420 0.000 41.700 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.900 0.000 59.180 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.380 0.000 76.660 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.860 0.000 94.140 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.340 0.000 111.620 2.400 ;
    END
  END address[5]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 6.840 137.630 7.440 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 12.280 137.630 12.880 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 17.040 137.630 17.640 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 22.480 137.630 23.080 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 27.920 137.630 28.520 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 32.680 137.630 33.280 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 38.120 137.630 38.720 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 43.560 137.630 44.160 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 48.320 137.630 48.920 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.230 53.760 137.630 54.360 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.230 58.520 137.630 59.120 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.230 63.960 137.630 64.560 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.230 69.400 137.630 70.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.230 74.160 137.630 74.760 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.230 79.600 137.630 80.200 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.230 85.040 137.630 85.640 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.230 89.800 137.630 90.400 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.230 95.240 137.630 95.840 ;
    END
  END chanx_right_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.420 137.600 41.700 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.480 137.600 46.760 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.540 137.600 51.820 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.600 137.600 56.880 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.120 137.600 62.400 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.180 137.600 67.460 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.240 137.600 72.520 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.300 137.600 77.580 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.820 137.600 83.100 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.880 137.600 88.160 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.940 137.600 93.220 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.000 137.600 98.280 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.520 137.600 103.800 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.580 137.600 108.860 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.640 137.600 113.920 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.700 137.600 118.980 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.220 137.600 124.500 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.280 137.600 129.560 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.820 0.000 129.100 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.460 0.000 6.740 2.400 ;
    END
  END enable
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 126.520 137.630 127.120 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 131.280 137.630 131.880 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 136.720 137.630 137.320 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 100.000 137.630 100.600 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 105.440 137.630 106.040 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 110.880 137.630 111.480 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 115.640 137.630 116.240 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 121.080 137.630 121.680 ;
    END
  END right_bottom_grid_pin_9_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.230 2.080 137.630 2.680 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.780 137.600 26.060 140.000 ;
    END
  END top_left_grid_pin_11_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.840 137.600 31.120 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.900 137.600 36.180 140.000 ;
    END
  END top_left_grid_pin_15_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.020 137.600 0.300 140.000 ;
    END
  END top_left_grid_pin_1_
  PIN top_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.080 137.600 5.360 140.000 ;
    END
  END top_left_grid_pin_3_
  PIN top_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.140 137.600 10.420 140.000 ;
    END
  END top_left_grid_pin_5_
  PIN top_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.200 137.600 15.480 140.000 ;
    END
  END top_left_grid_pin_7_
  PIN top_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.720 137.600 21.000 140.000 ;
    END
  END top_left_grid_pin_9_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.340 137.600 134.620 140.000 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 25.685 10.640 27.285 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 49.015 10.640 50.615 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 3.150 10.795 131.950 127.925 ;
      LAYER met1 ;
        RECT 0.000 0.380 136.020 128.080 ;
      LAYER met2 ;
        RECT 0.580 137.320 4.800 137.770 ;
        RECT 5.640 137.320 9.860 137.770 ;
        RECT 10.700 137.320 14.920 137.770 ;
        RECT 15.760 137.320 20.440 137.770 ;
        RECT 21.280 137.320 25.500 137.770 ;
        RECT 26.340 137.320 30.560 137.770 ;
        RECT 31.400 137.320 35.620 137.770 ;
        RECT 36.460 137.320 41.140 137.770 ;
        RECT 41.980 137.320 46.200 137.770 ;
        RECT 47.040 137.320 51.260 137.770 ;
        RECT 52.100 137.320 56.320 137.770 ;
        RECT 57.160 137.320 61.840 137.770 ;
        RECT 62.680 137.320 66.900 137.770 ;
        RECT 67.740 137.320 71.960 137.770 ;
        RECT 72.800 137.320 77.020 137.770 ;
        RECT 77.860 137.320 82.540 137.770 ;
        RECT 83.380 137.320 87.600 137.770 ;
        RECT 88.440 137.320 92.660 137.770 ;
        RECT 93.500 137.320 97.720 137.770 ;
        RECT 98.560 137.320 103.240 137.770 ;
        RECT 104.080 137.320 108.300 137.770 ;
        RECT 109.140 137.320 113.360 137.770 ;
        RECT 114.200 137.320 118.420 137.770 ;
        RECT 119.260 137.320 123.940 137.770 ;
        RECT 124.780 137.320 129.000 137.770 ;
        RECT 129.840 137.320 134.060 137.770 ;
        RECT 134.900 137.320 136.000 137.770 ;
        RECT 0.030 2.680 136.000 137.320 ;
        RECT 0.030 0.270 6.180 2.680 ;
        RECT 7.020 0.270 23.660 2.680 ;
        RECT 24.500 0.270 41.140 2.680 ;
        RECT 41.980 0.270 58.620 2.680 ;
        RECT 59.460 0.270 76.100 2.680 ;
        RECT 76.940 0.270 93.580 2.680 ;
        RECT 94.420 0.270 111.060 2.680 ;
        RECT 111.900 0.270 128.540 2.680 ;
        RECT 129.380 0.270 136.000 2.680 ;
      LAYER met3 ;
        RECT 25.680 136.320 134.830 136.720 ;
        RECT 25.680 132.280 136.280 136.320 ;
        RECT 25.680 130.880 134.830 132.280 ;
        RECT 25.680 127.520 136.280 130.880 ;
        RECT 25.680 126.120 134.830 127.520 ;
        RECT 25.680 122.080 136.280 126.120 ;
        RECT 25.680 120.680 134.830 122.080 ;
        RECT 25.680 116.640 136.280 120.680 ;
        RECT 25.680 115.240 134.830 116.640 ;
        RECT 25.680 111.880 136.280 115.240 ;
        RECT 25.680 110.480 134.830 111.880 ;
        RECT 25.680 106.440 136.280 110.480 ;
        RECT 25.680 105.040 134.830 106.440 ;
        RECT 25.680 101.000 136.280 105.040 ;
        RECT 25.680 99.600 134.830 101.000 ;
        RECT 25.680 96.240 136.280 99.600 ;
        RECT 25.680 94.840 134.830 96.240 ;
        RECT 25.680 90.800 136.280 94.840 ;
        RECT 25.680 89.400 134.830 90.800 ;
        RECT 25.680 86.040 136.280 89.400 ;
        RECT 25.680 84.640 134.830 86.040 ;
        RECT 25.680 80.600 136.280 84.640 ;
        RECT 25.680 79.200 134.830 80.600 ;
        RECT 25.680 75.160 136.280 79.200 ;
        RECT 25.680 73.760 134.830 75.160 ;
        RECT 25.680 70.400 136.280 73.760 ;
        RECT 25.680 69.000 134.830 70.400 ;
        RECT 25.680 64.960 136.280 69.000 ;
        RECT 25.680 63.560 134.830 64.960 ;
        RECT 25.680 59.520 136.280 63.560 ;
        RECT 25.680 58.120 134.830 59.520 ;
        RECT 25.680 54.760 136.280 58.120 ;
        RECT 25.680 53.360 134.830 54.760 ;
        RECT 25.680 49.320 136.280 53.360 ;
        RECT 25.680 47.920 134.830 49.320 ;
        RECT 25.680 44.560 136.280 47.920 ;
        RECT 25.680 43.160 134.830 44.560 ;
        RECT 25.680 39.120 136.280 43.160 ;
        RECT 25.680 37.720 134.830 39.120 ;
        RECT 25.680 33.680 136.280 37.720 ;
        RECT 25.680 32.280 134.830 33.680 ;
        RECT 25.680 28.920 136.280 32.280 ;
        RECT 25.680 27.520 134.830 28.920 ;
        RECT 25.680 23.480 136.280 27.520 ;
        RECT 25.680 22.080 134.830 23.480 ;
        RECT 25.680 18.040 136.280 22.080 ;
        RECT 25.680 16.640 134.830 18.040 ;
        RECT 25.680 13.280 136.280 16.640 ;
        RECT 25.680 11.880 134.830 13.280 ;
        RECT 25.680 7.840 136.280 11.880 ;
        RECT 25.680 7.440 134.830 7.840 ;
      LAYER met4 ;
        RECT 27.685 10.640 48.615 128.080 ;
        RECT 51.015 10.640 136.255 128.080 ;
  END
END sb_0__0_
END LIBRARY

