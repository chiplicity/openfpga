VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__1_
  CLASS BLOCK ;
  FOREIGN sb_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN bottom_left_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 2.400 ;
    END
  END bottom_left_grid_pin_34_
  PIN bottom_left_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 2.400 ;
    END
  END bottom_left_grid_pin_35_
  PIN bottom_left_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.400 ;
    END
  END bottom_left_grid_pin_36_
  PIN bottom_left_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END bottom_left_grid_pin_37_
  PIN bottom_left_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END bottom_left_grid_pin_38_
  PIN bottom_left_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 2.400 ;
    END
  END bottom_left_grid_pin_39_
  PIN bottom_left_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 2.400 ;
    END
  END bottom_left_grid_pin_40_
  PIN bottom_left_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 2.400 ;
    END
  END bottom_left_grid_pin_41_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 2.400 2.000 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 2.400 30.560 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 2.400 36.680 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.400 39.400 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 2.400 42.800 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 2.400 45.520 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 2.400 48.240 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 2.400 50.960 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 2.400 10.160 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.400 13.560 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 2.400 16.280 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.400 19.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 2.400 25.120 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 2.400 27.840 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 2.400 89.040 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 2.400 92.440 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 2.400 95.160 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 2.400 97.880 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 2.400 104.000 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.400 106.720 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.400 112.840 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 2.400 115.560 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 2.400 72.040 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.400 83.600 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.400 86.320 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 1.400 140.000 2.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 29.960 140.000 30.560 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 33.360 140.000 33.960 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 36.080 140.000 36.680 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.800 140.000 39.400 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 42.200 140.000 42.800 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.920 140.000 45.520 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 47.640 140.000 48.240 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 50.360 140.000 50.960 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 53.760 140.000 54.360 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 56.480 140.000 57.080 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 4.120 140.000 4.720 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 6.840 140.000 7.440 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 9.560 140.000 10.160 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 12.960 140.000 13.560 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 15.680 140.000 16.280 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 18.400 140.000 19.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 21.800 140.000 22.400 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 24.520 140.000 25.120 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 27.240 140.000 27.840 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 59.200 140.000 59.800 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 88.440 140.000 89.040 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 91.840 140.000 92.440 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 94.560 140.000 95.160 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 97.280 140.000 97.880 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 100.000 140.000 100.600 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 103.400 140.000 104.000 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 106.120 140.000 106.720 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 108.840 140.000 109.440 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 112.240 140.000 112.840 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 114.960 140.000 115.560 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 62.600 140.000 63.200 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 65.320 140.000 65.920 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 68.040 140.000 68.640 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 71.440 140.000 72.040 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 74.160 140.000 74.760 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 76.880 140.000 77.480 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 79.600 140.000 80.200 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 83.000 140.000 83.600 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 85.720 140.000 86.320 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.400 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 137.600 24.750 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 137.600 54.190 140.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 137.600 56.950 140.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 137.600 59.710 140.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 137.600 62.930 140.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 137.600 65.690 140.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 137.600 68.450 140.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.390 137.600 71.670 140.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.150 137.600 74.430 140.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 137.600 77.190 140.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 137.600 80.410 140.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 137.600 27.970 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 137.600 30.730 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 137.600 33.490 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 137.600 36.710 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.190 137.600 39.470 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 137.600 42.230 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 137.600 45.450 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 137.600 48.210 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 137.600 50.970 140.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 137.600 83.170 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.870 137.600 112.150 140.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 137.600 115.370 140.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.850 137.600 118.130 140.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 137.600 120.890 140.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 137.600 124.110 140.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 137.600 126.870 140.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.350 137.600 129.630 140.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 137.600 132.850 140.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 137.600 135.610 140.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.090 137.600 138.370 140.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 137.600 85.930 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 137.600 89.150 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.630 137.600 91.910 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.390 137.600 94.670 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 137.600 97.890 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 137.600 100.650 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.130 137.600 103.410 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.350 137.600 106.630 140.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.110 137.600 109.390 140.000 ;
    END
  END chany_top_out[9]
  PIN left_top_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 2.400 118.280 ;
    END
  END left_top_grid_pin_42_
  PIN left_top_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 2.400 121.000 ;
    END
  END left_top_grid_pin_43_
  PIN left_top_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 2.400 124.400 ;
    END
  END left_top_grid_pin_44_
  PIN left_top_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END left_top_grid_pin_45_
  PIN left_top_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 2.400 129.840 ;
    END
  END left_top_grid_pin_46_
  PIN left_top_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 2.400 133.240 ;
    END
  END left_top_grid_pin_47_
  PIN left_top_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 2.400 135.960 ;
    END
  END left_top_grid_pin_48_
  PIN left_top_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 2.400 138.680 ;
    END
  END left_top_grid_pin_49_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END prog_clk
  PIN right_top_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 117.680 140.000 118.280 ;
    END
  END right_top_grid_pin_42_
  PIN right_top_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 120.400 140.000 121.000 ;
    END
  END right_top_grid_pin_43_
  PIN right_top_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 123.800 140.000 124.400 ;
    END
  END right_top_grid_pin_44_
  PIN right_top_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 126.520 140.000 127.120 ;
    END
  END right_top_grid_pin_45_
  PIN right_top_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.240 140.000 129.840 ;
    END
  END right_top_grid_pin_46_
  PIN right_top_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 132.640 140.000 133.240 ;
    END
  END right_top_grid_pin_47_
  PIN right_top_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 135.360 140.000 135.960 ;
    END
  END right_top_grid_pin_48_
  PIN right_top_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 138.080 140.000 138.680 ;
    END
  END right_top_grid_pin_49_
  PIN top_left_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 137.600 1.750 140.000 ;
    END
  END top_left_grid_pin_34_
  PIN top_left_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 137.600 4.510 140.000 ;
    END
  END top_left_grid_pin_35_
  PIN top_left_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 137.600 7.270 140.000 ;
    END
  END top_left_grid_pin_36_
  PIN top_left_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 137.600 10.490 140.000 ;
    END
  END top_left_grid_pin_37_
  PIN top_left_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 137.600 13.250 140.000 ;
    END
  END top_left_grid_pin_38_
  PIN top_left_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 137.600 16.010 140.000 ;
    END
  END top_left_grid_pin_39_
  PIN top_left_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 137.600 19.230 140.000 ;
    END
  END top_left_grid_pin_40_
  PIN top_left_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 137.600 21.990 140.000 ;
    END
  END top_left_grid_pin_41_
  PIN vpwr
    USE POWER ; 
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ; 
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 132.855 ;
      LAYER met1 ;
        RECT 2.830 1.060 134.320 134.260 ;
      LAYER met2 ;
        RECT 0.090 137.320 1.190 138.565 ;
        RECT 2.030 137.320 3.950 138.565 ;
        RECT 4.790 137.320 6.710 138.565 ;
        RECT 7.550 137.320 9.930 138.565 ;
        RECT 10.770 137.320 12.690 138.565 ;
        RECT 13.530 137.320 15.450 138.565 ;
        RECT 16.290 137.320 18.670 138.565 ;
        RECT 19.510 137.320 21.430 138.565 ;
        RECT 22.270 137.320 24.190 138.565 ;
        RECT 25.030 137.320 27.410 138.565 ;
        RECT 28.250 137.320 30.170 138.565 ;
        RECT 31.010 137.320 32.930 138.565 ;
        RECT 33.770 137.320 36.150 138.565 ;
        RECT 36.990 137.320 38.910 138.565 ;
        RECT 39.750 137.320 41.670 138.565 ;
        RECT 42.510 137.320 44.890 138.565 ;
        RECT 45.730 137.320 47.650 138.565 ;
        RECT 48.490 137.320 50.410 138.565 ;
        RECT 51.250 137.320 53.630 138.565 ;
        RECT 54.470 137.320 56.390 138.565 ;
        RECT 57.230 137.320 59.150 138.565 ;
        RECT 59.990 137.320 62.370 138.565 ;
        RECT 63.210 137.320 65.130 138.565 ;
        RECT 65.970 137.320 67.890 138.565 ;
        RECT 68.730 137.320 71.110 138.565 ;
        RECT 71.950 137.320 73.870 138.565 ;
        RECT 74.710 137.320 76.630 138.565 ;
        RECT 77.470 137.320 79.850 138.565 ;
        RECT 80.690 137.320 82.610 138.565 ;
        RECT 83.450 137.320 85.370 138.565 ;
        RECT 86.210 137.320 88.590 138.565 ;
        RECT 89.430 137.320 91.350 138.565 ;
        RECT 92.190 137.320 94.110 138.565 ;
        RECT 94.950 137.320 97.330 138.565 ;
        RECT 98.170 137.320 100.090 138.565 ;
        RECT 100.930 137.320 102.850 138.565 ;
        RECT 103.690 137.320 106.070 138.565 ;
        RECT 106.910 137.320 108.830 138.565 ;
        RECT 109.670 137.320 111.590 138.565 ;
        RECT 112.430 137.320 114.810 138.565 ;
        RECT 115.650 137.320 117.570 138.565 ;
        RECT 118.410 137.320 120.330 138.565 ;
        RECT 121.170 137.320 123.550 138.565 ;
        RECT 124.390 137.320 126.310 138.565 ;
        RECT 127.150 137.320 129.070 138.565 ;
        RECT 129.910 137.320 132.290 138.565 ;
        RECT 133.130 137.320 135.050 138.565 ;
        RECT 135.890 137.320 137.810 138.565 ;
        RECT 0.090 2.680 138.370 137.320 ;
        RECT 0.090 0.155 0.730 2.680 ;
        RECT 1.570 0.155 3.030 2.680 ;
        RECT 3.870 0.155 5.790 2.680 ;
        RECT 6.630 0.155 8.550 2.680 ;
        RECT 9.390 0.155 11.310 2.680 ;
        RECT 12.150 0.155 14.070 2.680 ;
        RECT 14.910 0.155 16.830 2.680 ;
        RECT 17.670 0.155 19.590 2.680 ;
        RECT 20.430 0.155 22.350 2.680 ;
        RECT 23.190 0.155 25.110 2.680 ;
        RECT 25.950 0.155 27.870 2.680 ;
        RECT 28.710 0.155 30.630 2.680 ;
        RECT 31.470 0.155 33.390 2.680 ;
        RECT 34.230 0.155 36.150 2.680 ;
        RECT 36.990 0.155 38.910 2.680 ;
        RECT 39.750 0.155 41.670 2.680 ;
        RECT 42.510 0.155 44.430 2.680 ;
        RECT 45.270 0.155 47.190 2.680 ;
        RECT 48.030 0.155 49.950 2.680 ;
        RECT 50.790 0.155 52.710 2.680 ;
        RECT 53.550 0.155 55.470 2.680 ;
        RECT 56.310 0.155 58.230 2.680 ;
        RECT 59.070 0.155 60.990 2.680 ;
        RECT 61.830 0.155 63.750 2.680 ;
        RECT 64.590 0.155 66.510 2.680 ;
        RECT 67.350 0.155 69.270 2.680 ;
        RECT 70.110 0.155 71.570 2.680 ;
        RECT 72.410 0.155 74.330 2.680 ;
        RECT 75.170 0.155 77.090 2.680 ;
        RECT 77.930 0.155 79.850 2.680 ;
        RECT 80.690 0.155 82.610 2.680 ;
        RECT 83.450 0.155 85.370 2.680 ;
        RECT 86.210 0.155 88.130 2.680 ;
        RECT 88.970 0.155 90.890 2.680 ;
        RECT 91.730 0.155 93.650 2.680 ;
        RECT 94.490 0.155 96.410 2.680 ;
        RECT 97.250 0.155 99.170 2.680 ;
        RECT 100.010 0.155 101.930 2.680 ;
        RECT 102.770 0.155 104.690 2.680 ;
        RECT 105.530 0.155 107.450 2.680 ;
        RECT 108.290 0.155 110.210 2.680 ;
        RECT 111.050 0.155 112.970 2.680 ;
        RECT 113.810 0.155 115.730 2.680 ;
        RECT 116.570 0.155 118.490 2.680 ;
        RECT 119.330 0.155 121.250 2.680 ;
        RECT 122.090 0.155 124.010 2.680 ;
        RECT 124.850 0.155 126.770 2.680 ;
        RECT 127.610 0.155 129.530 2.680 ;
        RECT 130.370 0.155 132.290 2.680 ;
        RECT 133.130 0.155 135.050 2.680 ;
        RECT 135.890 0.155 137.810 2.680 ;
      LAYER met3 ;
        RECT 2.800 137.680 137.200 138.545 ;
        RECT 0.065 136.360 138.395 137.680 ;
        RECT 2.800 134.960 137.200 136.360 ;
        RECT 0.065 133.640 138.395 134.960 ;
        RECT 2.800 132.240 137.200 133.640 ;
        RECT 0.065 130.240 138.395 132.240 ;
        RECT 2.800 128.840 137.200 130.240 ;
        RECT 0.065 127.520 138.395 128.840 ;
        RECT 2.800 126.120 137.200 127.520 ;
        RECT 0.065 124.800 138.395 126.120 ;
        RECT 2.800 123.400 137.200 124.800 ;
        RECT 0.065 121.400 138.395 123.400 ;
        RECT 2.800 120.000 137.200 121.400 ;
        RECT 0.065 118.680 138.395 120.000 ;
        RECT 2.800 117.280 137.200 118.680 ;
        RECT 0.065 115.960 138.395 117.280 ;
        RECT 2.800 114.560 137.200 115.960 ;
        RECT 0.065 113.240 138.395 114.560 ;
        RECT 2.800 111.840 137.200 113.240 ;
        RECT 0.065 109.840 138.395 111.840 ;
        RECT 2.800 108.440 137.200 109.840 ;
        RECT 0.065 107.120 138.395 108.440 ;
        RECT 2.800 105.720 137.200 107.120 ;
        RECT 0.065 104.400 138.395 105.720 ;
        RECT 2.800 103.000 137.200 104.400 ;
        RECT 0.065 101.000 138.395 103.000 ;
        RECT 2.800 99.600 137.200 101.000 ;
        RECT 0.065 98.280 138.395 99.600 ;
        RECT 2.800 96.880 137.200 98.280 ;
        RECT 0.065 95.560 138.395 96.880 ;
        RECT 2.800 94.160 137.200 95.560 ;
        RECT 0.065 92.840 138.395 94.160 ;
        RECT 2.800 91.440 137.200 92.840 ;
        RECT 0.065 89.440 138.395 91.440 ;
        RECT 2.800 88.040 137.200 89.440 ;
        RECT 0.065 86.720 138.395 88.040 ;
        RECT 2.800 85.320 137.200 86.720 ;
        RECT 0.065 84.000 138.395 85.320 ;
        RECT 2.800 82.600 137.200 84.000 ;
        RECT 0.065 80.600 138.395 82.600 ;
        RECT 2.800 79.200 137.200 80.600 ;
        RECT 0.065 77.880 138.395 79.200 ;
        RECT 2.800 76.480 137.200 77.880 ;
        RECT 0.065 75.160 138.395 76.480 ;
        RECT 2.800 73.760 137.200 75.160 ;
        RECT 0.065 72.440 138.395 73.760 ;
        RECT 2.800 71.040 137.200 72.440 ;
        RECT 0.065 69.040 138.395 71.040 ;
        RECT 2.800 67.640 137.200 69.040 ;
        RECT 0.065 66.320 138.395 67.640 ;
        RECT 2.800 64.920 137.200 66.320 ;
        RECT 0.065 63.600 138.395 64.920 ;
        RECT 2.800 62.200 137.200 63.600 ;
        RECT 0.065 60.200 138.395 62.200 ;
        RECT 2.800 58.800 137.200 60.200 ;
        RECT 0.065 57.480 138.395 58.800 ;
        RECT 2.800 56.080 137.200 57.480 ;
        RECT 0.065 54.760 138.395 56.080 ;
        RECT 2.800 53.360 137.200 54.760 ;
        RECT 0.065 51.360 138.395 53.360 ;
        RECT 2.800 49.960 137.200 51.360 ;
        RECT 0.065 48.640 138.395 49.960 ;
        RECT 2.800 47.240 137.200 48.640 ;
        RECT 0.065 45.920 138.395 47.240 ;
        RECT 2.800 44.520 137.200 45.920 ;
        RECT 0.065 43.200 138.395 44.520 ;
        RECT 2.800 41.800 137.200 43.200 ;
        RECT 0.065 39.800 138.395 41.800 ;
        RECT 2.800 38.400 137.200 39.800 ;
        RECT 0.065 37.080 138.395 38.400 ;
        RECT 2.800 35.680 137.200 37.080 ;
        RECT 0.065 34.360 138.395 35.680 ;
        RECT 2.800 32.960 137.200 34.360 ;
        RECT 0.065 30.960 138.395 32.960 ;
        RECT 2.800 29.560 137.200 30.960 ;
        RECT 0.065 28.240 138.395 29.560 ;
        RECT 2.800 26.840 137.200 28.240 ;
        RECT 0.065 25.520 138.395 26.840 ;
        RECT 2.800 24.120 137.200 25.520 ;
        RECT 0.065 22.800 138.395 24.120 ;
        RECT 2.800 21.400 137.200 22.800 ;
        RECT 0.065 19.400 138.395 21.400 ;
        RECT 2.800 18.000 137.200 19.400 ;
        RECT 0.065 16.680 138.395 18.000 ;
        RECT 2.800 15.280 137.200 16.680 ;
        RECT 0.065 13.960 138.395 15.280 ;
        RECT 2.800 12.560 137.200 13.960 ;
        RECT 0.065 10.560 138.395 12.560 ;
        RECT 2.800 9.160 137.200 10.560 ;
        RECT 0.065 7.840 138.395 9.160 ;
        RECT 2.800 6.440 137.200 7.840 ;
        RECT 0.065 5.120 138.395 6.440 ;
        RECT 2.800 3.720 137.200 5.120 ;
        RECT 0.065 2.400 138.395 3.720 ;
        RECT 2.800 1.000 137.200 2.400 ;
        RECT 0.065 0.175 138.395 1.000 ;
      LAYER met4 ;
        RECT 7.230 128.480 134.450 133.105 ;
        RECT 7.230 10.240 27.655 128.480 ;
        RECT 30.055 10.240 50.985 128.480 ;
        RECT 53.385 10.240 134.450 128.480 ;
        RECT 7.230 0.855 134.450 10.240 ;
      LAYER met5 ;
        RECT 7.020 4.300 134.660 128.300 ;
  END
END sb_1__1_
END LIBRARY

