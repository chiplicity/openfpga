VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__3_
  CLASS BLOCK ;
  FOREIGN cbx_1__3_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 80.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.070 77.600 6.350 80.000 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 77.600 18.770 80.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 77.600 31.190 80.000 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 2.400 14.240 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 77.600 43.610 80.000 ;
    END
  END address[6]
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.750 77.600 56.030 80.000 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 77.600 68.450 80.000 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 2.760 200.000 3.360 ;
    END
  END bottom_grid_pin_8_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 8.880 200.000 9.480 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.050 77.600 81.330 80.000 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 2.400 20.360 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.470 77.600 93.750 80.000 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 15.680 200.000 16.280 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 77.600 106.170 80.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.400 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 22.480 200.000 23.080 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 29.280 200.000 29.880 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.310 77.600 118.590 80.000 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 2.400 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 2.400 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 36.080 200.000 36.680 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 42.880 200.000 43.480 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 77.600 131.010 80.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 49.000 200.000 49.600 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.610 77.600 143.890 80.000 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.030 77.600 156.310 80.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 55.800 200.000 56.400 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 62.600 200.000 63.200 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 2.400 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 2.400 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.450 77.600 168.730 80.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.400 37.360 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 69.400 200.000 70.000 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.870 77.600 181.150 80.000 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 2.400 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 2.400 60.480 ;
    END
  END chanx_right_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END enable
  PIN top_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 76.200 200.000 76.800 ;
    END
  END top_grid_pin_0_
  PIN top_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END top_grid_pin_10_
  PIN top_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.290 77.600 193.570 80.000 ;
    END
  END top_grid_pin_12_
  PIN top_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 2.400 ;
    END
  END top_grid_pin_14_
  PIN top_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END top_grid_pin_2_
  PIN top_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 2.400 ;
    END
  END top_grid_pin_4_
  PIN top_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 2.400 72.040 ;
    END
  END top_grid_pin_6_
  PIN top_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 2.400 ;
    END
  END top_grid_pin_8_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 38.055 10.640 39.655 68.240 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 71.385 10.640 72.985 68.240 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 68.085 ;
      LAYER met1 ;
        RECT 0.070 0.380 198.190 78.160 ;
      LAYER met2 ;
        RECT 0.090 77.320 5.790 78.190 ;
        RECT 6.630 77.320 18.210 78.190 ;
        RECT 19.050 77.320 30.630 78.190 ;
        RECT 31.470 77.320 43.050 78.190 ;
        RECT 43.890 77.320 55.470 78.190 ;
        RECT 56.310 77.320 67.890 78.190 ;
        RECT 68.730 77.320 80.770 78.190 ;
        RECT 81.610 77.320 93.190 78.190 ;
        RECT 94.030 77.320 105.610 78.190 ;
        RECT 106.450 77.320 118.030 78.190 ;
        RECT 118.870 77.320 130.450 78.190 ;
        RECT 131.290 77.320 143.330 78.190 ;
        RECT 144.170 77.320 155.750 78.190 ;
        RECT 156.590 77.320 168.170 78.190 ;
        RECT 169.010 77.320 180.590 78.190 ;
        RECT 181.430 77.320 193.010 78.190 ;
        RECT 193.850 77.320 198.170 78.190 ;
        RECT 0.090 2.680 198.170 77.320 ;
        RECT 0.090 0.155 6.710 2.680 ;
        RECT 7.550 0.155 20.970 2.680 ;
        RECT 21.810 0.155 35.230 2.680 ;
        RECT 36.070 0.155 49.490 2.680 ;
        RECT 50.330 0.155 63.750 2.680 ;
        RECT 64.590 0.155 78.010 2.680 ;
        RECT 78.850 0.155 92.270 2.680 ;
        RECT 93.110 0.155 106.530 2.680 ;
        RECT 107.370 0.155 120.790 2.680 ;
        RECT 121.630 0.155 135.050 2.680 ;
        RECT 135.890 0.155 149.310 2.680 ;
        RECT 150.150 0.155 163.570 2.680 ;
        RECT 164.410 0.155 177.830 2.680 ;
        RECT 178.670 0.155 192.090 2.680 ;
        RECT 192.930 0.155 198.170 2.680 ;
      LAYER met3 ;
        RECT 2.800 76.480 197.200 76.880 ;
        RECT 0.310 75.800 197.200 76.480 ;
        RECT 0.310 72.440 198.450 75.800 ;
        RECT 2.800 71.040 198.450 72.440 ;
        RECT 0.310 70.400 198.450 71.040 ;
        RECT 0.310 69.000 197.200 70.400 ;
        RECT 0.310 66.320 198.450 69.000 ;
        RECT 2.800 64.920 198.450 66.320 ;
        RECT 0.310 63.600 198.450 64.920 ;
        RECT 0.310 62.200 197.200 63.600 ;
        RECT 0.310 60.880 198.450 62.200 ;
        RECT 2.800 59.480 198.450 60.880 ;
        RECT 0.310 56.800 198.450 59.480 ;
        RECT 0.310 55.400 197.200 56.800 ;
        RECT 0.310 54.760 198.450 55.400 ;
        RECT 2.800 53.360 198.450 54.760 ;
        RECT 0.310 50.000 198.450 53.360 ;
        RECT 0.310 49.320 197.200 50.000 ;
        RECT 2.800 48.600 197.200 49.320 ;
        RECT 2.800 47.920 198.450 48.600 ;
        RECT 0.310 43.880 198.450 47.920 ;
        RECT 2.800 42.480 197.200 43.880 ;
        RECT 0.310 37.760 198.450 42.480 ;
        RECT 2.800 37.080 198.450 37.760 ;
        RECT 2.800 36.360 197.200 37.080 ;
        RECT 0.310 35.680 197.200 36.360 ;
        RECT 0.310 32.320 198.450 35.680 ;
        RECT 2.800 30.920 198.450 32.320 ;
        RECT 0.310 30.280 198.450 30.920 ;
        RECT 0.310 28.880 197.200 30.280 ;
        RECT 0.310 26.200 198.450 28.880 ;
        RECT 2.800 24.800 198.450 26.200 ;
        RECT 0.310 23.480 198.450 24.800 ;
        RECT 0.310 22.080 197.200 23.480 ;
        RECT 0.310 20.760 198.450 22.080 ;
        RECT 2.800 19.360 198.450 20.760 ;
        RECT 0.310 16.680 198.450 19.360 ;
        RECT 0.310 15.280 197.200 16.680 ;
        RECT 0.310 14.640 198.450 15.280 ;
        RECT 2.800 13.240 198.450 14.640 ;
        RECT 0.310 9.880 198.450 13.240 ;
        RECT 0.310 9.200 197.200 9.880 ;
        RECT 2.800 8.480 197.200 9.200 ;
        RECT 2.800 7.800 198.450 8.480 ;
        RECT 0.310 3.760 198.450 7.800 ;
        RECT 2.800 2.360 197.200 3.760 ;
        RECT 0.310 0.175 198.450 2.360 ;
      LAYER met4 ;
        RECT 40.055 10.640 70.985 68.240 ;
        RECT 73.385 10.640 198.425 68.240 ;
      LAYER met5 ;
        RECT 47.500 51.900 118.100 53.500 ;
  END
END cbx_1__3_
END LIBRARY

